magic
tech EFS8A
magscale 1 2
timestamp 1602524379
<< locali >>
rect 9919 35785 10057 35819
rect 7475 33065 7481 33099
rect 7475 32997 7509 33065
rect 8211 30889 8217 30923
rect 8211 30821 8245 30889
rect 8217 27523 8251 27557
rect 8217 27489 8378 27523
rect 9321 26911 9355 27013
rect 1995 26401 2030 26435
rect 3007 26401 3042 26435
rect 4295 25925 4387 25959
rect 4353 25687 4387 25925
rect 11287 25313 11322 25347
rect 1869 24225 2030 24259
rect 1869 24191 1903 24225
rect 7199 23511 7233 23579
rect 7199 23477 7205 23511
rect 11287 22049 11322 22083
rect 8119 21097 8125 21131
rect 8119 21029 8153 21097
rect 4629 19873 4755 19907
rect 4629 19703 4663 19873
rect 8159 18785 8194 18819
rect 2605 18275 2639 18377
rect 12851 16609 12886 16643
rect 11287 15521 11322 15555
rect 5267 14807 5301 14875
rect 5267 14773 5273 14807
rect 6469 13719 6503 14025
rect 4353 12767 4387 12937
rect 1777 8415 1811 8517
rect 8211 8041 8217 8075
rect 5376 7973 5444 8007
rect 8211 7973 8245 8041
rect 8211 6953 8217 6987
rect 8211 6885 8245 6953
rect 10977 6239 11011 6409
rect 5583 5729 5710 5763
rect 6469 5151 6503 5321
rect 8125 5151 8159 5321
rect 3065 4063 3099 4097
rect 3065 4029 3226 4063
rect 6279 3689 6285 3723
rect 6279 3621 6313 3689
rect 8159 3621 8204 3655
rect 7239 2533 7284 2567
<< viali >>
rect 10057 35785 10091 35819
rect 6904 35581 6938 35615
rect 7297 35581 7331 35615
rect 8953 35581 8987 35615
rect 9816 35581 9850 35615
rect 10241 35581 10275 35615
rect 8125 35513 8159 35547
rect 8309 35513 8343 35547
rect 8401 35513 8435 35547
rect 6975 35445 7009 35479
rect 6837 35241 6871 35275
rect 8493 35241 8527 35275
rect 9873 35241 9907 35275
rect 7113 35173 7147 35207
rect 5968 35105 6002 35139
rect 9689 35105 9723 35139
rect 6055 35037 6089 35071
rect 6469 35037 6503 35071
rect 7021 35037 7055 35071
rect 7665 35037 7699 35071
rect 8309 34901 8343 34935
rect 5549 34697 5583 34731
rect 6193 34697 6227 34731
rect 9689 34697 9723 34731
rect 10241 34697 10275 34731
rect 12633 34697 12667 34731
rect 5825 34629 5859 34663
rect 7573 34629 7607 34663
rect 7021 34561 7055 34595
rect 8585 34561 8619 34595
rect 9229 34561 9263 34595
rect 5641 34493 5675 34527
rect 10057 34493 10091 34527
rect 10609 34493 10643 34527
rect 12449 34493 12483 34527
rect 13001 34493 13035 34527
rect 6653 34425 6687 34459
rect 7113 34425 7147 34459
rect 8677 34425 8711 34459
rect 7941 34357 7975 34391
rect 8401 34357 8435 34391
rect 8309 34153 8343 34187
rect 8585 34153 8619 34187
rect 7710 34085 7744 34119
rect 9873 34085 9907 34119
rect 6101 34017 6135 34051
rect 6285 34017 6319 34051
rect 6561 34017 6595 34051
rect 7389 34017 7423 34051
rect 4813 33949 4847 33983
rect 9781 33949 9815 33983
rect 10057 33949 10091 33983
rect 7021 33813 7055 33847
rect 7757 33609 7791 33643
rect 9505 33609 9539 33643
rect 10149 33609 10183 33643
rect 4537 33541 4571 33575
rect 4813 33405 4847 33439
rect 5089 33405 5123 33439
rect 6561 33405 6595 33439
rect 6837 33405 6871 33439
rect 8585 33405 8619 33439
rect 5917 33337 5951 33371
rect 7159 33337 7193 33371
rect 8033 33337 8067 33371
rect 8401 33337 8435 33371
rect 8906 33337 8940 33371
rect 4721 33269 4755 33303
rect 6193 33269 6227 33303
rect 9781 33269 9815 33303
rect 4629 33065 4663 33099
rect 7481 33065 7515 33099
rect 8033 33065 8067 33099
rect 5134 32997 5168 33031
rect 4813 32861 4847 32895
rect 7113 32861 7147 32895
rect 8585 32793 8619 32827
rect 5733 32725 5767 32759
rect 6009 32725 6043 32759
rect 6561 32725 6595 32759
rect 6929 32725 6963 32759
rect 10057 32725 10091 32759
rect 7849 32521 7883 32555
rect 6561 32453 6595 32487
rect 4353 32385 4387 32419
rect 5273 32385 5307 32419
rect 6193 32385 6227 32419
rect 3525 32317 3559 32351
rect 3617 32317 3651 32351
rect 4077 32317 4111 32351
rect 6837 32317 6871 32351
rect 7389 32317 7423 32351
rect 8677 32317 8711 32351
rect 8861 32317 8895 32351
rect 9965 32317 9999 32351
rect 10425 32317 10459 32351
rect 5365 32249 5399 32283
rect 5917 32249 5951 32283
rect 8309 32249 8343 32283
rect 4905 32181 4939 32215
rect 6929 32181 6963 32215
rect 8493 32181 8527 32215
rect 9781 32181 9815 32215
rect 10057 32181 10091 32215
rect 3709 31977 3743 32011
rect 4813 31977 4847 32011
rect 9781 31977 9815 32011
rect 11391 31977 11425 32011
rect 5318 31909 5352 31943
rect 6929 31909 6963 31943
rect 7849 31909 7883 31943
rect 9689 31841 9723 31875
rect 10241 31841 10275 31875
rect 11320 31841 11354 31875
rect 4997 31773 5031 31807
rect 6837 31773 6871 31807
rect 7113 31773 7147 31807
rect 5917 31637 5951 31671
rect 8493 31637 8527 31671
rect 10701 31637 10735 31671
rect 7389 31433 7423 31467
rect 11437 31433 11471 31467
rect 5825 31365 5859 31399
rect 7021 31365 7055 31399
rect 10701 31365 10735 31399
rect 4813 31297 4847 31331
rect 7849 31297 7883 31331
rect 8309 31297 8343 31331
rect 10149 31297 10183 31331
rect 3617 31229 3651 31263
rect 3893 31229 3927 31263
rect 4077 31229 4111 31263
rect 4905 31229 4939 31263
rect 6101 31229 6135 31263
rect 9689 31229 9723 31263
rect 3249 31161 3283 31195
rect 5226 31161 5260 31195
rect 8630 31161 8664 31195
rect 10241 31161 10275 31195
rect 4445 31093 4479 31127
rect 8125 31093 8159 31127
rect 9229 31093 9263 31127
rect 11069 31093 11103 31127
rect 3433 30889 3467 30923
rect 8217 30889 8251 30923
rect 8769 30889 8803 30923
rect 10701 30889 10735 30923
rect 4491 30821 4525 30855
rect 5641 30821 5675 30855
rect 6193 30821 6227 30855
rect 9873 30821 9907 30855
rect 10425 30821 10459 30855
rect 4404 30753 4438 30787
rect 5549 30685 5583 30719
rect 7849 30685 7883 30719
rect 9781 30685 9815 30719
rect 11253 30685 11287 30719
rect 4997 30549 5031 30583
rect 3893 30345 3927 30379
rect 5825 30345 5859 30379
rect 9781 30345 9815 30379
rect 11437 30345 11471 30379
rect 7757 30277 7791 30311
rect 8125 30277 8159 30311
rect 9229 30277 9263 30311
rect 8309 30209 8343 30243
rect 10425 30209 10459 30243
rect 4629 30141 4663 30175
rect 4721 30141 4755 30175
rect 5181 30141 5215 30175
rect 6872 30141 6906 30175
rect 7297 30141 7331 30175
rect 4261 30073 4295 30107
rect 8630 30073 8664 30107
rect 10149 30073 10183 30107
rect 10241 30073 10275 30107
rect 11069 30073 11103 30107
rect 4813 30005 4847 30039
rect 6101 30005 6135 30039
rect 6975 30005 7009 30039
rect 4169 29801 4203 29835
rect 8401 29801 8435 29835
rect 9781 29801 9815 29835
rect 10701 29801 10735 29835
rect 6837 29733 6871 29767
rect 7021 29733 7055 29767
rect 7113 29733 7147 29767
rect 8033 29733 8067 29767
rect 4077 29665 4111 29699
rect 4537 29665 4571 29699
rect 5952 29665 5986 29699
rect 8560 29665 8594 29699
rect 9689 29665 9723 29699
rect 10149 29665 10183 29699
rect 7665 29597 7699 29631
rect 6055 29461 6089 29495
rect 8631 29461 8665 29495
rect 8953 29461 8987 29495
rect 5917 29257 5951 29291
rect 9689 29189 9723 29223
rect 3341 29121 3375 29155
rect 4169 29121 4203 29155
rect 6929 29121 6963 29155
rect 7573 29121 7607 29155
rect 8493 29121 8527 29155
rect 9137 29121 9171 29155
rect 4077 28985 4111 29019
rect 4490 28985 4524 29019
rect 7021 28985 7055 29019
rect 8585 28985 8619 29019
rect 3709 28917 3743 28951
rect 5089 28917 5123 28951
rect 6653 28917 6687 28951
rect 7849 28917 7883 28951
rect 8309 28917 8343 28951
rect 10057 28917 10091 28951
rect 1593 28713 1627 28747
rect 4353 28713 4387 28747
rect 7389 28713 7423 28747
rect 4813 28645 4847 28679
rect 6514 28645 6548 28679
rect 8125 28645 8159 28679
rect 8953 28645 8987 28679
rect 1409 28577 1443 28611
rect 3008 28577 3042 28611
rect 7113 28577 7147 28611
rect 9756 28577 9790 28611
rect 3111 28509 3145 28543
rect 4721 28509 4755 28543
rect 5365 28509 5399 28543
rect 6193 28509 6227 28543
rect 8033 28509 8067 28543
rect 8309 28509 8343 28543
rect 5641 28373 5675 28407
rect 7757 28373 7791 28407
rect 9827 28373 9861 28407
rect 10149 28373 10183 28407
rect 4813 28169 4847 28203
rect 6193 28169 6227 28203
rect 6975 28169 7009 28203
rect 9781 28169 9815 28203
rect 3433 28101 3467 28135
rect 7941 28101 7975 28135
rect 3019 28033 3053 28067
rect 4997 28033 5031 28067
rect 5641 28033 5675 28067
rect 9965 28033 9999 28067
rect 10241 28033 10275 28067
rect 1685 27965 1719 27999
rect 2932 27965 2966 27999
rect 3960 27965 3994 27999
rect 6872 27965 6906 27999
rect 8125 27965 8159 27999
rect 4353 27897 4387 27931
rect 5089 27897 5123 27931
rect 6561 27897 6595 27931
rect 8446 27897 8480 27931
rect 9413 27897 9447 27931
rect 10057 27897 10091 27931
rect 3709 27829 3743 27863
rect 4031 27829 4065 27863
rect 7297 27829 7331 27863
rect 9045 27829 9079 27863
rect 3525 27625 3559 27659
rect 4353 27625 4387 27659
rect 4721 27625 4755 27659
rect 7297 27625 7331 27659
rect 7941 27625 7975 27659
rect 11621 27625 11655 27659
rect 5549 27557 5583 27591
rect 6698 27557 6732 27591
rect 8217 27557 8251 27591
rect 9873 27557 9907 27591
rect 4813 27489 4847 27523
rect 5273 27489 5307 27523
rect 11437 27489 11471 27523
rect 6377 27421 6411 27455
rect 8447 27421 8481 27455
rect 9781 27421 9815 27455
rect 10241 27421 10275 27455
rect 8769 27353 8803 27387
rect 5825 27285 5859 27319
rect 9137 27285 9171 27319
rect 4537 27081 4571 27115
rect 6377 27081 6411 27115
rect 7941 27081 7975 27115
rect 8401 27081 8435 27115
rect 11069 27081 11103 27115
rect 4905 27013 4939 27047
rect 9321 27013 9355 27047
rect 5089 26945 5123 26979
rect 8585 26945 8619 26979
rect 9229 26945 9263 26979
rect 3709 26877 3743 26911
rect 3985 26877 4019 26911
rect 6929 26877 6963 26911
rect 7389 26877 7423 26911
rect 9321 26877 9355 26911
rect 9965 26877 9999 26911
rect 10057 26877 10091 26911
rect 10517 26877 10551 26911
rect 3341 26809 3375 26843
rect 4169 26809 4203 26843
rect 5181 26809 5215 26843
rect 5733 26809 5767 26843
rect 7665 26809 7699 26843
rect 8677 26809 8711 26843
rect 6009 26741 6043 26775
rect 9505 26741 9539 26775
rect 10149 26741 10183 26775
rect 11437 26741 11471 26775
rect 3433 26537 3467 26571
rect 7113 26537 7147 26571
rect 8769 26537 8803 26571
rect 9045 26537 9079 26571
rect 9413 26537 9447 26571
rect 4715 26469 4749 26503
rect 6285 26469 6319 26503
rect 8170 26469 8204 26503
rect 9873 26469 9907 26503
rect 10425 26469 10459 26503
rect 1961 26401 1995 26435
rect 2973 26401 3007 26435
rect 11304 26401 11338 26435
rect 4353 26333 4387 26367
rect 6193 26333 6227 26367
rect 6653 26333 6687 26367
rect 7849 26333 7883 26367
rect 9781 26333 9815 26367
rect 11391 26333 11425 26367
rect 2099 26265 2133 26299
rect 3111 26197 3145 26231
rect 5273 26197 5307 26231
rect 5549 26197 5583 26231
rect 2605 25993 2639 26027
rect 4537 25993 4571 26027
rect 6193 25993 6227 26027
rect 6469 25993 6503 26027
rect 9689 25993 9723 26027
rect 10885 25993 10919 26027
rect 2053 25925 2087 25959
rect 4261 25925 4295 25959
rect 5641 25925 5675 25959
rect 2421 25789 2455 25823
rect 3709 25789 3743 25823
rect 3893 25789 3927 25823
rect 4169 25789 4203 25823
rect 8125 25857 8159 25891
rect 10241 25857 10275 25891
rect 6872 25789 6906 25823
rect 7297 25789 7331 25823
rect 5089 25721 5123 25755
rect 5181 25721 5215 25755
rect 8446 25721 8480 25755
rect 9965 25721 9999 25755
rect 10057 25721 10091 25755
rect 3065 25653 3099 25687
rect 4353 25653 4387 25687
rect 4905 25653 4939 25687
rect 6975 25653 7009 25687
rect 7941 25653 7975 25687
rect 9045 25653 9079 25687
rect 9413 25653 9447 25687
rect 11345 25653 11379 25687
rect 3157 25449 3191 25483
rect 4353 25449 4387 25483
rect 5825 25449 5859 25483
rect 8631 25449 8665 25483
rect 8953 25449 8987 25483
rect 10701 25449 10735 25483
rect 11391 25449 11425 25483
rect 4950 25381 4984 25415
rect 7665 25381 7699 25415
rect 8309 25381 8343 25415
rect 9873 25381 9907 25415
rect 2973 25313 3007 25347
rect 5549 25313 5583 25347
rect 6929 25313 6963 25347
rect 7389 25313 7423 25347
rect 8528 25313 8562 25347
rect 11253 25313 11287 25347
rect 3525 25245 3559 25279
rect 4629 25245 4663 25279
rect 9781 25245 9815 25279
rect 10149 25245 10183 25279
rect 2513 25177 2547 25211
rect 6837 25109 6871 25143
rect 7941 25109 7975 25143
rect 4169 24905 4203 24939
rect 4905 24905 4939 24939
rect 9505 24905 9539 24939
rect 9735 24905 9769 24939
rect 10425 24905 10459 24939
rect 11253 24905 11287 24939
rect 3157 24837 3191 24871
rect 4629 24837 4663 24871
rect 6193 24837 6227 24871
rect 9137 24837 9171 24871
rect 5641 24769 5675 24803
rect 7113 24769 7147 24803
rect 2973 24701 3007 24735
rect 3985 24701 4019 24735
rect 8636 24701 8670 24735
rect 9664 24701 9698 24735
rect 10057 24701 10091 24735
rect 5181 24633 5215 24667
rect 5273 24633 5307 24667
rect 7205 24633 7239 24667
rect 7757 24633 7791 24667
rect 8401 24633 8435 24667
rect 8723 24633 8757 24667
rect 3433 24565 3467 24599
rect 3893 24565 3927 24599
rect 6561 24565 6595 24599
rect 8033 24565 8067 24599
rect 3111 24361 3145 24395
rect 3893 24361 3927 24395
rect 4445 24361 4479 24395
rect 5733 24361 5767 24395
rect 6423 24361 6457 24395
rect 2099 24293 2133 24327
rect 6101 24293 6135 24327
rect 7481 24293 7515 24327
rect 3008 24225 3042 24259
rect 4629 24225 4663 24259
rect 4813 24225 4847 24259
rect 6320 24225 6354 24259
rect 1869 24157 1903 24191
rect 7389 24157 7423 24191
rect 8033 24157 8067 24191
rect 6837 24089 6871 24123
rect 1685 24021 1719 24055
rect 3433 24021 3467 24055
rect 5457 24021 5491 24055
rect 8677 24021 8711 24055
rect 1547 23817 1581 23851
rect 2881 23817 2915 23851
rect 4997 23817 5031 23851
rect 6285 23817 6319 23851
rect 13645 23817 13679 23851
rect 3525 23749 3559 23783
rect 10287 23749 10321 23783
rect 8677 23681 8711 23715
rect 8953 23681 8987 23715
rect 1476 23613 1510 23647
rect 3433 23613 3467 23647
rect 3709 23613 3743 23647
rect 5181 23613 5215 23647
rect 5641 23613 5675 23647
rect 6837 23613 6871 23647
rect 7757 23613 7791 23647
rect 10184 23613 10218 23647
rect 10609 23613 10643 23647
rect 13461 23613 13495 23647
rect 14013 23613 14047 23647
rect 5917 23545 5951 23579
rect 8493 23545 8527 23579
rect 8769 23545 8803 23579
rect 2053 23477 2087 23511
rect 3249 23477 3283 23511
rect 3893 23477 3927 23511
rect 4537 23477 4571 23511
rect 7205 23477 7239 23511
rect 8033 23477 8067 23511
rect 1593 23273 1627 23307
rect 4445 23273 4479 23307
rect 7849 23273 7883 23307
rect 6647 23205 6681 23239
rect 8217 23205 8251 23239
rect 8769 23205 8803 23239
rect 9781 23205 9815 23239
rect 9873 23205 9907 23239
rect 1409 23137 1443 23171
rect 3040 23137 3074 23171
rect 4721 23137 4755 23171
rect 5273 23137 5307 23171
rect 5457 23069 5491 23103
rect 6285 23069 6319 23103
rect 8125 23069 8159 23103
rect 10057 23069 10091 23103
rect 3111 23001 3145 23035
rect 7205 23001 7239 23035
rect 3433 22933 3467 22967
rect 3893 22933 3927 22967
rect 7481 22933 7515 22967
rect 9045 22933 9079 22967
rect 1685 22729 1719 22763
rect 2697 22729 2731 22763
rect 4721 22729 4755 22763
rect 6285 22729 6319 22763
rect 6653 22729 6687 22763
rect 7941 22729 7975 22763
rect 10149 22729 10183 22763
rect 10471 22661 10505 22695
rect 3249 22593 3283 22627
rect 3893 22593 3927 22627
rect 7021 22593 7055 22627
rect 9781 22593 9815 22627
rect 2212 22525 2246 22559
rect 3157 22525 3191 22559
rect 3433 22525 3467 22559
rect 4169 22525 4203 22559
rect 5181 22525 5215 22559
rect 5641 22525 5675 22559
rect 5917 22525 5951 22559
rect 10400 22525 10434 22559
rect 10793 22525 10827 22559
rect 7342 22457 7376 22491
rect 8861 22457 8895 22491
rect 8953 22457 8987 22491
rect 9505 22457 9539 22491
rect 2283 22389 2317 22423
rect 2973 22389 3007 22423
rect 8217 22389 8251 22423
rect 8677 22389 8711 22423
rect 6285 22185 6319 22219
rect 7481 22185 7515 22219
rect 9045 22185 9079 22219
rect 11391 22185 11425 22219
rect 3157 22117 3191 22151
rect 3893 22117 3927 22151
rect 6653 22117 6687 22151
rect 7205 22117 7239 22151
rect 8217 22117 8251 22151
rect 9873 22117 9907 22151
rect 1409 22049 1443 22083
rect 3065 22049 3099 22083
rect 4169 22049 4203 22083
rect 4445 22049 4479 22083
rect 11253 22049 11287 22083
rect 2329 21981 2363 22015
rect 4905 21981 4939 22015
rect 6561 21981 6595 22015
rect 8125 21981 8159 22015
rect 9781 21981 9815 22015
rect 10057 21981 10091 22015
rect 3433 21913 3467 21947
rect 4261 21913 4295 21947
rect 8677 21913 8711 21947
rect 1869 21845 1903 21879
rect 5181 21845 5215 21879
rect 5641 21845 5675 21879
rect 7849 21845 7883 21879
rect 2605 21641 2639 21675
rect 4169 21641 4203 21675
rect 4813 21641 4847 21675
rect 6561 21641 6595 21675
rect 7297 21641 7331 21675
rect 8677 21641 8711 21675
rect 8953 21641 8987 21675
rect 9965 21641 9999 21675
rect 5825 21573 5859 21607
rect 10333 21573 10367 21607
rect 10977 21505 11011 21539
rect 1593 21437 1627 21471
rect 3065 21437 3099 21471
rect 3157 21437 3191 21471
rect 3341 21437 3375 21471
rect 4905 21437 4939 21471
rect 6101 21437 6135 21471
rect 7757 21437 7791 21471
rect 10517 21437 10551 21471
rect 2237 21369 2271 21403
rect 3801 21369 3835 21403
rect 5226 21369 5260 21403
rect 7573 21369 7607 21403
rect 8078 21369 8112 21403
rect 11345 21369 11379 21403
rect 2973 21301 3007 21335
rect 9505 21301 9539 21335
rect 10701 21301 10735 21335
rect 1869 21097 1903 21131
rect 2237 21097 2271 21131
rect 3433 21097 3467 21131
rect 4905 21097 4939 21131
rect 7205 21097 7239 21131
rect 8125 21097 8159 21131
rect 8677 21097 8711 21131
rect 3157 21029 3191 21063
rect 6929 21029 6963 21063
rect 9781 21029 9815 21063
rect 9873 21029 9907 21063
rect 1409 20961 1443 20995
rect 2421 20961 2455 20995
rect 2697 20961 2731 20995
rect 3801 20961 3835 20995
rect 4445 20961 4479 20995
rect 4721 20961 4755 20995
rect 6193 20961 6227 20995
rect 6745 20961 6779 20995
rect 7757 20893 7791 20927
rect 1593 20825 1627 20859
rect 2513 20825 2547 20859
rect 4537 20825 4571 20859
rect 10333 20825 10367 20859
rect 4353 20757 4387 20791
rect 5549 20757 5583 20791
rect 7573 20757 7607 20791
rect 9045 20757 9079 20791
rect 4077 20553 4111 20587
rect 5273 20553 5307 20587
rect 5917 20553 5951 20587
rect 8125 20553 8159 20587
rect 9689 20553 9723 20587
rect 10149 20553 10183 20587
rect 1869 20485 1903 20519
rect 9137 20485 9171 20519
rect 10885 20485 10919 20519
rect 4721 20417 4755 20451
rect 8217 20417 8251 20451
rect 1685 20349 1719 20383
rect 2605 20349 2639 20383
rect 3341 20349 3375 20383
rect 4261 20349 4295 20383
rect 4353 20349 4387 20383
rect 4537 20349 4571 20383
rect 6193 20349 6227 20383
rect 7021 20349 7055 20383
rect 7665 20349 7699 20383
rect 9965 20349 9999 20383
rect 10517 20349 10551 20383
rect 3433 20281 3467 20315
rect 3709 20281 3743 20315
rect 6561 20281 6595 20315
rect 6837 20281 6871 20315
rect 8538 20281 8572 20315
rect 2237 20213 2271 20247
rect 7113 20213 7147 20247
rect 1961 20009 1995 20043
rect 3433 20009 3467 20043
rect 4813 20009 4847 20043
rect 7205 20009 7239 20043
rect 9781 20009 9815 20043
rect 2329 19941 2363 19975
rect 6423 19941 6457 19975
rect 7843 19941 7877 19975
rect 8677 19941 8711 19975
rect 1409 19873 1443 19907
rect 3065 19873 3099 19907
rect 5181 19873 5215 19907
rect 6336 19873 6370 19907
rect 9689 19873 9723 19907
rect 10149 19873 10183 19907
rect 3157 19805 3191 19839
rect 7481 19805 7515 19839
rect 6101 19737 6135 19771
rect 1593 19669 1627 19703
rect 3801 19669 3835 19703
rect 4445 19669 4479 19703
rect 4629 19669 4663 19703
rect 5825 19669 5859 19703
rect 6929 19669 6963 19703
rect 8401 19669 8435 19703
rect 4629 19465 4663 19499
rect 2513 19397 2547 19431
rect 3387 19397 3421 19431
rect 3525 19397 3559 19431
rect 4905 19397 4939 19431
rect 7941 19397 7975 19431
rect 9229 19397 9263 19431
rect 2145 19329 2179 19363
rect 3157 19329 3191 19363
rect 3617 19329 3651 19363
rect 7573 19329 7607 19363
rect 8493 19329 8527 19363
rect 8677 19329 8711 19363
rect 10149 19329 10183 19363
rect 1501 19261 1535 19295
rect 4813 19261 4847 19295
rect 5089 19261 5123 19295
rect 7113 19261 7147 19295
rect 7297 19261 7331 19295
rect 3249 19193 3283 19227
rect 8769 19193 8803 19227
rect 10609 19193 10643 19227
rect 3893 19125 3927 19159
rect 4261 19125 4295 19159
rect 5273 19125 5307 19159
rect 5825 19125 5859 19159
rect 6377 19125 6411 19159
rect 9689 19125 9723 19159
rect 2881 18921 2915 18955
rect 3801 18921 3835 18955
rect 6009 18921 6043 18955
rect 8585 18921 8619 18955
rect 9781 18921 9815 18955
rect 2329 18853 2363 18887
rect 5175 18853 5209 18887
rect 7297 18853 7331 18887
rect 7573 18853 7607 18887
rect 1409 18785 1443 18819
rect 2421 18785 2455 18819
rect 2697 18785 2731 18819
rect 6377 18785 6411 18819
rect 6561 18785 6595 18819
rect 7113 18785 7147 18819
rect 8125 18785 8159 18819
rect 9689 18785 9723 18819
rect 10149 18785 10183 18819
rect 3433 18717 3467 18751
rect 4813 18717 4847 18751
rect 1593 18649 1627 18683
rect 2513 18649 2547 18683
rect 4629 18649 4663 18683
rect 1869 18581 1903 18615
rect 5733 18581 5767 18615
rect 8263 18581 8297 18615
rect 10701 18581 10735 18615
rect 2421 18377 2455 18411
rect 2605 18377 2639 18411
rect 2789 18377 2823 18411
rect 4077 18377 4111 18411
rect 4353 18377 4387 18411
rect 8125 18377 8159 18411
rect 10149 18377 10183 18411
rect 1869 18309 1903 18343
rect 3065 18309 3099 18343
rect 5549 18309 5583 18343
rect 2605 18241 2639 18275
rect 3433 18241 3467 18275
rect 6929 18241 6963 18275
rect 7205 18241 7239 18275
rect 9781 18241 9815 18275
rect 10425 18241 10459 18275
rect 10701 18241 10735 18275
rect 2012 18173 2046 18207
rect 2973 18173 3007 18207
rect 3249 18173 3283 18207
rect 4721 18173 4755 18207
rect 4997 18173 5031 18207
rect 6193 18173 6227 18207
rect 2099 18105 2133 18139
rect 5273 18105 5307 18139
rect 7021 18105 7055 18139
rect 8861 18105 8895 18139
rect 8953 18105 8987 18139
rect 9505 18105 9539 18139
rect 10517 18105 10551 18139
rect 6653 18037 6687 18071
rect 8585 18037 8619 18071
rect 1593 17833 1627 17867
rect 1961 17833 1995 17867
rect 3341 17833 3375 17867
rect 5273 17833 5307 17867
rect 7205 17833 7239 17867
rect 4353 17765 4387 17799
rect 5549 17765 5583 17799
rect 5825 17765 5859 17799
rect 5917 17765 5951 17799
rect 9873 17765 9907 17799
rect 2973 17697 3007 17731
rect 7297 17697 7331 17731
rect 7849 17697 7883 17731
rect 11288 17697 11322 17731
rect 2329 17629 2363 17663
rect 4261 17629 4295 17663
rect 6745 17629 6779 17663
rect 8033 17629 8067 17663
rect 9505 17629 9539 17663
rect 9781 17629 9815 17663
rect 10425 17629 10459 17663
rect 4813 17561 4847 17595
rect 6377 17561 6411 17595
rect 10701 17561 10735 17595
rect 8861 17493 8895 17527
rect 11391 17493 11425 17527
rect 2237 17289 2271 17323
rect 4077 17289 4111 17323
rect 4997 17289 5031 17323
rect 12587 17289 12621 17323
rect 13001 17289 13035 17323
rect 13645 17289 13679 17323
rect 4307 17221 4341 17255
rect 11713 17221 11747 17255
rect 2697 17153 2731 17187
rect 5273 17153 5307 17187
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 9229 17153 9263 17187
rect 11069 17153 11103 17187
rect 4236 17085 4270 17119
rect 4629 17085 4663 17119
rect 5917 17085 5951 17119
rect 12516 17085 12550 17119
rect 13461 17085 13495 17119
rect 1869 17017 1903 17051
rect 2421 17017 2455 17051
rect 2513 17017 2547 17051
rect 5365 17017 5399 17051
rect 6561 17017 6595 17051
rect 7710 17017 7744 17051
rect 8585 17017 8619 17051
rect 9321 17017 9355 17051
rect 9873 17017 9907 17051
rect 10793 17017 10827 17051
rect 10885 17017 10919 17051
rect 14013 17017 14047 17051
rect 3341 16949 3375 16983
rect 6193 16949 6227 16983
rect 8309 16949 8343 16983
rect 9045 16949 9079 16983
rect 10149 16949 10183 16983
rect 10517 16949 10551 16983
rect 1409 16745 1443 16779
rect 7481 16745 7515 16779
rect 8585 16745 8619 16779
rect 10701 16745 10735 16779
rect 2329 16677 2363 16711
rect 2605 16677 2639 16711
rect 4261 16677 4295 16711
rect 5917 16677 5951 16711
rect 6009 16677 6043 16711
rect 7986 16677 8020 16711
rect 9873 16677 9907 16711
rect 11437 16677 11471 16711
rect 11989 16677 12023 16711
rect 6929 16609 6963 16643
rect 12817 16609 12851 16643
rect 2513 16541 2547 16575
rect 4169 16541 4203 16575
rect 4813 16541 4847 16575
rect 6193 16541 6227 16575
rect 7665 16541 7699 16575
rect 9781 16541 9815 16575
rect 10425 16541 10459 16575
rect 11345 16541 11379 16575
rect 3065 16473 3099 16507
rect 1869 16405 1903 16439
rect 3433 16405 3467 16439
rect 5273 16405 5307 16439
rect 5641 16405 5675 16439
rect 9229 16405 9263 16439
rect 12955 16405 12989 16439
rect 4261 16201 4295 16235
rect 6193 16201 6227 16235
rect 7297 16201 7331 16235
rect 8309 16201 8343 16235
rect 10057 16201 10091 16235
rect 10793 16201 10827 16235
rect 11345 16201 11379 16235
rect 11713 16201 11747 16235
rect 12173 16201 12207 16235
rect 2053 16133 2087 16167
rect 8953 16133 8987 16167
rect 11023 16133 11057 16167
rect 1501 16065 1535 16099
rect 5089 16065 5123 16099
rect 9137 16065 9171 16099
rect 10333 16065 10367 16099
rect 2513 15997 2547 16031
rect 2973 15997 3007 16031
rect 6653 15997 6687 16031
rect 7389 15997 7423 16031
rect 10952 15997 10986 16031
rect 1593 15929 1627 15963
rect 3294 15929 3328 15963
rect 4813 15929 4847 15963
rect 4905 15929 4939 15963
rect 7710 15929 7744 15963
rect 9499 15929 9533 15963
rect 2789 15861 2823 15895
rect 3893 15861 3927 15895
rect 4537 15861 4571 15895
rect 5917 15861 5951 15895
rect 8585 15861 8619 15895
rect 12817 15861 12851 15895
rect 1685 15657 1719 15691
rect 2145 15657 2179 15691
rect 3157 15657 3191 15691
rect 6423 15657 6457 15691
rect 8861 15657 8895 15691
rect 11391 15657 11425 15691
rect 12403 15657 12437 15691
rect 2558 15589 2592 15623
rect 4858 15589 4892 15623
rect 6837 15589 6871 15623
rect 7802 15589 7836 15623
rect 9137 15589 9171 15623
rect 9873 15589 9907 15623
rect 10425 15589 10459 15623
rect 5457 15521 5491 15555
rect 6320 15521 6354 15555
rect 11253 15521 11287 15555
rect 12332 15521 12366 15555
rect 2237 15453 2271 15487
rect 3433 15453 3467 15487
rect 4537 15453 4571 15487
rect 7481 15453 7515 15487
rect 9781 15453 9815 15487
rect 5825 15385 5859 15419
rect 3801 15317 3835 15351
rect 4445 15317 4479 15351
rect 7205 15317 7239 15351
rect 8401 15317 8435 15351
rect 2329 15113 2363 15147
rect 5825 15113 5859 15147
rect 6285 15113 6319 15147
rect 8677 15113 8711 15147
rect 9873 15113 9907 15147
rect 10241 15113 10275 15147
rect 12633 15113 12667 15147
rect 4445 15045 4479 15079
rect 4813 15045 4847 15079
rect 7849 15045 7883 15079
rect 11437 15045 11471 15079
rect 4905 14977 4939 15011
rect 8953 14977 8987 15011
rect 9597 14977 9631 15011
rect 10793 14977 10827 15011
rect 1593 14909 1627 14943
rect 2789 14909 2823 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 6837 14909 6871 14943
rect 7389 14909 7423 14943
rect 1409 14841 1443 14875
rect 1961 14841 1995 14875
rect 2697 14841 2731 14875
rect 9045 14841 9079 14875
rect 10517 14841 10551 14875
rect 10609 14841 10643 14875
rect 2881 14773 2915 14807
rect 5273 14773 5307 14807
rect 6929 14773 6963 14807
rect 8217 14773 8251 14807
rect 1547 14569 1581 14603
rect 4353 14569 4387 14603
rect 6101 14569 6135 14603
rect 9505 14569 9539 14603
rect 9965 14569 9999 14603
rect 10701 14569 10735 14603
rect 3157 14501 3191 14535
rect 5502 14501 5536 14535
rect 7665 14501 7699 14535
rect 1476 14433 1510 14467
rect 2513 14433 2547 14467
rect 3433 14433 3467 14467
rect 4169 14433 4203 14467
rect 6929 14433 6963 14467
rect 7389 14433 7423 14467
rect 8528 14433 8562 14467
rect 9689 14433 9723 14467
rect 10149 14433 10183 14467
rect 1961 14365 1995 14399
rect 5181 14365 5215 14399
rect 8953 14365 8987 14399
rect 2329 14229 2363 14263
rect 4813 14229 4847 14263
rect 8631 14229 8665 14263
rect 1593 14025 1627 14059
rect 2697 14025 2731 14059
rect 4629 14025 4663 14059
rect 5733 14025 5767 14059
rect 6469 14025 6503 14059
rect 7941 14025 7975 14059
rect 8309 14025 8343 14059
rect 9689 14025 9723 14059
rect 10103 14025 10137 14059
rect 2053 13957 2087 13991
rect 3525 13889 3559 13923
rect 1409 13821 1443 13855
rect 2881 13821 2915 13855
rect 3617 13821 3651 13855
rect 4997 13821 5031 13855
rect 5273 13821 5307 13855
rect 6193 13753 6227 13787
rect 10425 13889 10459 13923
rect 6929 13821 6963 13855
rect 7389 13821 7423 13855
rect 8401 13821 8435 13855
rect 8861 13821 8895 13855
rect 10016 13821 10050 13855
rect 2881 13685 2915 13719
rect 4169 13685 4203 13719
rect 4813 13685 4847 13719
rect 6469 13685 6503 13719
rect 6561 13685 6595 13719
rect 6929 13685 6963 13719
rect 8677 13685 8711 13719
rect 1685 13481 1719 13515
rect 2421 13481 2455 13515
rect 3157 13481 3191 13515
rect 3433 13481 3467 13515
rect 4537 13481 4571 13515
rect 5181 13481 5215 13515
rect 6285 13481 6319 13515
rect 7021 13481 7055 13515
rect 10149 13481 10183 13515
rect 5727 13413 5761 13447
rect 8217 13413 8251 13447
rect 1961 13345 1995 13379
rect 2973 13345 3007 13379
rect 4353 13345 4387 13379
rect 9724 13345 9758 13379
rect 2881 13277 2915 13311
rect 5365 13277 5399 13311
rect 8125 13277 8159 13311
rect 9827 13277 9861 13311
rect 2145 13209 2179 13243
rect 7297 13209 7331 13243
rect 8677 13209 8711 13243
rect 4813 13141 4847 13175
rect 2237 12937 2271 12971
rect 2605 12937 2639 12971
rect 2881 12937 2915 12971
rect 4353 12937 4387 12971
rect 4537 12937 4571 12971
rect 6193 12937 6227 12971
rect 10517 12937 10551 12971
rect 3893 12869 3927 12903
rect 3249 12801 3283 12835
rect 9781 12869 9815 12903
rect 5273 12801 5307 12835
rect 8493 12801 8527 12835
rect 8769 12801 8803 12835
rect 1685 12733 1719 12767
rect 2697 12733 2731 12767
rect 3709 12733 3743 12767
rect 4353 12733 4387 12767
rect 4997 12733 5031 12767
rect 5181 12733 5215 12767
rect 6837 12733 6871 12767
rect 7297 12733 7331 12767
rect 10032 12733 10066 12767
rect 4261 12665 4295 12699
rect 8585 12665 8619 12699
rect 1869 12597 1903 12631
rect 3525 12597 3559 12631
rect 5825 12597 5859 12631
rect 6561 12597 6595 12631
rect 7113 12597 7147 12631
rect 7941 12597 7975 12631
rect 8217 12597 8251 12631
rect 10103 12597 10137 12631
rect 4629 12393 4663 12427
rect 6837 12393 6871 12427
rect 8493 12393 8527 12427
rect 8861 12393 8895 12427
rect 7342 12325 7376 12359
rect 9781 12325 9815 12359
rect 9873 12325 9907 12359
rect 1961 12257 1995 12291
rect 2973 12257 3007 12291
rect 3433 12257 3467 12291
rect 4445 12257 4479 12291
rect 5641 12257 5675 12291
rect 6009 12257 6043 12291
rect 11320 12257 11354 12291
rect 6193 12189 6227 12223
rect 7021 12189 7055 12223
rect 10241 12189 10275 12223
rect 1777 12121 1811 12155
rect 3157 12121 3191 12155
rect 7941 12121 7975 12155
rect 2145 12053 2179 12087
rect 4905 12053 4939 12087
rect 6469 12053 6503 12087
rect 11391 12053 11425 12087
rect 1593 11849 1627 11883
rect 2421 11849 2455 11883
rect 3433 11849 3467 11883
rect 4537 11849 4571 11883
rect 4997 11849 5031 11883
rect 6193 11849 6227 11883
rect 9873 11849 9907 11883
rect 2053 11781 2087 11815
rect 5917 11713 5951 11747
rect 8677 11713 8711 11747
rect 1409 11645 1443 11679
rect 3433 11645 3467 11679
rect 5273 11645 5307 11679
rect 5641 11645 5675 11679
rect 7021 11645 7055 11679
rect 8217 11645 8251 11679
rect 7342 11577 7376 11611
rect 8861 11577 8895 11611
rect 8953 11577 8987 11611
rect 9505 11577 9539 11611
rect 10425 11577 10459 11611
rect 10517 11577 10551 11611
rect 11069 11577 11103 11611
rect 3065 11509 3099 11543
rect 4169 11509 4203 11543
rect 6653 11509 6687 11543
rect 7941 11509 7975 11543
rect 10149 11509 10183 11543
rect 11437 11509 11471 11543
rect 1593 11305 1627 11339
rect 5181 11305 5215 11339
rect 5641 11305 5675 11339
rect 8217 11305 8251 11339
rect 9505 11305 9539 11339
rect 3157 11237 3191 11271
rect 7618 11237 7652 11271
rect 9873 11237 9907 11271
rect 11437 11237 11471 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 4077 11169 4111 11203
rect 4169 11169 4203 11203
rect 4353 11169 4387 11203
rect 5733 11169 5767 11203
rect 6193 11169 6227 11203
rect 2329 11101 2363 11135
rect 4537 11101 4571 11135
rect 6469 11101 6503 11135
rect 7297 11101 7331 11135
rect 9781 11101 9815 11135
rect 10241 11101 10275 11135
rect 10701 11101 10735 11135
rect 11345 11101 11379 11135
rect 11621 11101 11655 11135
rect 2513 11033 2547 11067
rect 3709 10965 3743 10999
rect 7021 10965 7055 10999
rect 8769 10965 8803 10999
rect 4997 10761 5031 10795
rect 6193 10761 6227 10795
rect 8585 10761 8619 10795
rect 8953 10761 8987 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 11621 10761 11655 10795
rect 8309 10693 8343 10727
rect 3157 10625 3191 10659
rect 3709 10625 3743 10659
rect 11253 10625 11287 10659
rect 1961 10557 1995 10591
rect 2697 10557 2731 10591
rect 3617 10557 3651 10591
rect 3893 10557 3927 10591
rect 4629 10557 4663 10591
rect 5457 10557 5491 10591
rect 5733 10557 5767 10591
rect 7389 10557 7423 10591
rect 2789 10489 2823 10523
rect 5917 10489 5951 10523
rect 6653 10489 6687 10523
rect 7297 10489 7331 10523
rect 7751 10489 7785 10523
rect 9229 10489 9263 10523
rect 9321 10489 9355 10523
rect 9873 10489 9907 10523
rect 3525 10421 3559 10455
rect 4077 10421 4111 10455
rect 2329 10217 2363 10251
rect 2881 10217 2915 10251
rect 5273 10217 5307 10251
rect 5641 10217 5675 10251
rect 8217 10217 8251 10251
rect 9229 10217 9263 10251
rect 9827 10217 9861 10251
rect 1685 10149 1719 10183
rect 6469 10149 6503 10183
rect 7113 10149 7147 10183
rect 7659 10149 7693 10183
rect 2421 10081 2455 10115
rect 2513 10081 2547 10115
rect 2697 10081 2731 10115
rect 4261 10081 4295 10115
rect 5733 10081 5767 10115
rect 6193 10081 6227 10115
rect 7297 10081 7331 10115
rect 9756 10081 9790 10115
rect 3709 10013 3743 10047
rect 4813 10013 4847 10047
rect 2145 9673 2179 9707
rect 2789 9673 2823 9707
rect 3157 9673 3191 9707
rect 3525 9673 3559 9707
rect 4997 9673 5031 9707
rect 5365 9673 5399 9707
rect 6009 9673 6043 9707
rect 8401 9673 8435 9707
rect 8907 9673 8941 9707
rect 9597 9673 9631 9707
rect 10333 9673 10367 9707
rect 11253 9673 11287 9707
rect 4077 9605 4111 9639
rect 5733 9605 5767 9639
rect 2513 9537 2547 9571
rect 4721 9537 4755 9571
rect 6561 9537 6595 9571
rect 2973 9469 3007 9503
rect 3985 9469 4019 9503
rect 4261 9469 4295 9503
rect 5549 9469 5583 9503
rect 7021 9469 7055 9503
rect 7573 9469 7607 9503
rect 8836 9469 8870 9503
rect 9848 9469 9882 9503
rect 10860 9469 10894 9503
rect 7757 9401 7791 9435
rect 9321 9401 9355 9435
rect 3801 9333 3835 9367
rect 8125 9333 8159 9367
rect 9919 9333 9953 9367
rect 10931 9333 10965 9367
rect 2973 9129 3007 9163
rect 5181 9129 5215 9163
rect 5549 9129 5583 9163
rect 4813 9061 4847 9095
rect 6101 9061 6135 9095
rect 9873 9061 9907 9095
rect 4077 8993 4111 9027
rect 4169 8993 4203 9027
rect 4353 8993 4387 9027
rect 7481 8993 7515 9027
rect 7941 8993 7975 9027
rect 11288 8993 11322 9027
rect 6009 8925 6043 8959
rect 6653 8925 6687 8959
rect 8217 8925 8251 8959
rect 9781 8925 9815 8959
rect 10333 8857 10367 8891
rect 7113 8789 7147 8823
rect 11391 8789 11425 8823
rect 1593 8585 1627 8619
rect 4629 8585 4663 8619
rect 4997 8585 5031 8619
rect 7849 8585 7883 8619
rect 10609 8585 10643 8619
rect 11529 8585 11563 8619
rect 1777 8517 1811 8551
rect 2053 8517 2087 8551
rect 4353 8517 4387 8551
rect 5825 8517 5859 8551
rect 7481 8517 7515 8551
rect 6929 8449 6963 8483
rect 9229 8449 9263 8483
rect 1409 8381 1443 8415
rect 1777 8381 1811 8415
rect 3192 8381 3226 8415
rect 3617 8381 3651 8415
rect 4169 8381 4203 8415
rect 10768 8381 10802 8415
rect 11161 8381 11195 8415
rect 3295 8313 3329 8347
rect 5273 8313 5307 8347
rect 5365 8313 5399 8347
rect 7021 8313 7055 8347
rect 9045 8313 9079 8347
rect 9298 8313 9332 8347
rect 9873 8313 9907 8347
rect 3985 8245 4019 8279
rect 6193 8245 6227 8279
rect 6653 8245 6687 8279
rect 8217 8245 8251 8279
rect 10241 8245 10275 8279
rect 10839 8245 10873 8279
rect 3111 8041 3145 8075
rect 3801 8041 3835 8075
rect 4215 8041 4249 8075
rect 6653 8041 6687 8075
rect 7297 8041 7331 8075
rect 8217 8041 8251 8075
rect 9229 8041 9263 8075
rect 4629 7973 4663 8007
rect 5342 7973 5376 8007
rect 9873 7973 9907 8007
rect 10425 7973 10459 8007
rect 3008 7905 3042 7939
rect 4144 7905 4178 7939
rect 6837 7905 6871 7939
rect 7849 7905 7883 7939
rect 11320 7905 11354 7939
rect 5089 7837 5123 7871
rect 9781 7837 9815 7871
rect 8769 7769 8803 7803
rect 3525 7701 3559 7735
rect 4997 7701 5031 7735
rect 6009 7701 6043 7735
rect 6285 7701 6319 7735
rect 7021 7701 7055 7735
rect 11391 7701 11425 7735
rect 2973 7497 3007 7531
rect 4445 7497 4479 7531
rect 5917 7497 5951 7531
rect 9689 7497 9723 7531
rect 9965 7497 9999 7531
rect 11529 7497 11563 7531
rect 6193 7429 6227 7463
rect 4169 7361 4203 7395
rect 4997 7361 5031 7395
rect 7021 7361 7055 7395
rect 8769 7361 8803 7395
rect 10609 7361 10643 7395
rect 10885 7361 10919 7395
rect 3433 7293 3467 7327
rect 3985 7293 4019 7327
rect 5318 7225 5352 7259
rect 7383 7225 7417 7259
rect 9090 7225 9124 7259
rect 10425 7225 10459 7259
rect 10701 7225 10735 7259
rect 4905 7157 4939 7191
rect 6561 7157 6595 7191
rect 7941 7157 7975 7191
rect 8217 7157 8251 7191
rect 8585 7157 8619 7191
rect 3433 6953 3467 6987
rect 7021 6953 7055 6987
rect 7757 6953 7791 6987
rect 8217 6953 8251 6987
rect 9045 6953 9079 6987
rect 9505 6953 9539 6987
rect 10701 6953 10735 6987
rect 5181 6885 5215 6919
rect 5825 6885 5859 6919
rect 6193 6885 6227 6919
rect 6745 6885 6779 6919
rect 9873 6885 9907 6919
rect 10425 6885 10459 6919
rect 4721 6817 4755 6851
rect 4905 6817 4939 6851
rect 12332 6817 12366 6851
rect 6101 6749 6135 6783
rect 7849 6749 7883 6783
rect 9781 6749 9815 6783
rect 11253 6749 11287 6783
rect 5457 6613 5491 6647
rect 8769 6613 8803 6647
rect 12403 6613 12437 6647
rect 5733 6409 5767 6443
rect 8953 6409 8987 6443
rect 10149 6409 10183 6443
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 11253 6409 11287 6443
rect 4077 6341 4111 6375
rect 6009 6341 6043 6375
rect 10839 6341 10873 6375
rect 7665 6273 7699 6307
rect 8309 6273 8343 6307
rect 9229 6273 9263 6307
rect 4445 6205 4479 6239
rect 4813 6205 4847 6239
rect 4997 6205 5031 6239
rect 6653 6205 6687 6239
rect 6929 6205 6963 6239
rect 7481 6205 7515 6239
rect 10768 6205 10802 6239
rect 10977 6205 11011 6239
rect 9321 6137 9355 6171
rect 9873 6137 9907 6171
rect 4629 6069 4663 6103
rect 8033 6069 8067 6103
rect 12633 6069 12667 6103
rect 4537 5865 4571 5899
rect 4905 5865 4939 5899
rect 5779 5865 5813 5899
rect 9229 5865 9263 5899
rect 7021 5797 7055 5831
rect 9873 5797 9907 5831
rect 10425 5797 10459 5831
rect 5549 5729 5583 5763
rect 7297 5729 7331 5763
rect 7849 5729 7883 5763
rect 8033 5661 8067 5695
rect 9781 5661 9815 5695
rect 8493 5525 8527 5559
rect 4537 5321 4571 5355
rect 6193 5321 6227 5355
rect 6469 5321 6503 5355
rect 4997 5185 5031 5219
rect 8125 5321 8159 5355
rect 8217 5321 8251 5355
rect 9781 5321 9815 5355
rect 10057 5321 10091 5355
rect 6929 5185 6963 5219
rect 7205 5185 7239 5219
rect 7941 5185 7975 5219
rect 6469 5117 6503 5151
rect 8125 5117 8159 5151
rect 8401 5117 8435 5151
rect 8953 5117 8987 5151
rect 5318 5049 5352 5083
rect 7021 5049 7055 5083
rect 4813 4981 4847 5015
rect 5917 4981 5951 5015
rect 6653 4981 6687 5015
rect 8493 4981 8527 5015
rect 5457 4777 5491 4811
rect 6929 4777 6963 4811
rect 7297 4777 7331 4811
rect 8585 4777 8619 4811
rect 9781 4777 9815 4811
rect 10701 4777 10735 4811
rect 6101 4709 6135 4743
rect 6653 4709 6687 4743
rect 7665 4709 7699 4743
rect 4629 4641 4663 4675
rect 4905 4641 4939 4675
rect 9689 4641 9723 4675
rect 10241 4641 10275 4675
rect 5089 4573 5123 4607
rect 6009 4573 6043 4607
rect 7573 4573 7607 4607
rect 7849 4573 7883 4607
rect 3709 4233 3743 4267
rect 4307 4233 4341 4267
rect 6561 4233 6595 4267
rect 9689 4233 9723 4267
rect 10977 4233 11011 4267
rect 4077 4165 4111 4199
rect 4997 4165 5031 4199
rect 6193 4165 6227 4199
rect 7481 4165 7515 4199
rect 3065 4097 3099 4131
rect 3295 4097 3329 4131
rect 8217 4097 8251 4131
rect 10057 4097 10091 4131
rect 10333 4097 10367 4131
rect 4236 4029 4270 4063
rect 5273 3961 5307 3995
rect 5365 3961 5399 3995
rect 5917 3961 5951 3995
rect 8538 3961 8572 3995
rect 10149 3961 10183 3995
rect 4721 3893 4755 3927
rect 6837 3893 6871 3927
rect 8125 3893 8159 3927
rect 9137 3893 9171 3927
rect 5733 3689 5767 3723
rect 6285 3689 6319 3723
rect 6837 3689 6871 3723
rect 7297 3689 7331 3723
rect 7757 3689 7791 3723
rect 8769 3689 8803 3723
rect 10701 3689 10735 3723
rect 8125 3621 8159 3655
rect 9873 3621 9907 3655
rect 4629 3553 4663 3587
rect 4905 3553 4939 3587
rect 7849 3553 7883 3587
rect 5089 3485 5123 3519
rect 5917 3485 5951 3519
rect 9045 3485 9079 3519
rect 9781 3485 9815 3519
rect 11253 3485 11287 3519
rect 10333 3417 10367 3451
rect 5457 3349 5491 3383
rect 4537 3145 4571 3179
rect 5917 3145 5951 3179
rect 6561 3145 6595 3179
rect 9505 3145 9539 3179
rect 11345 3145 11379 3179
rect 7021 3077 7055 3111
rect 4997 3009 5031 3043
rect 8217 3009 8251 3043
rect 9873 3009 9907 3043
rect 10057 3009 10091 3043
rect 3341 2941 3375 2975
rect 3709 2941 3743 2975
rect 3985 2941 4019 2975
rect 4169 2941 4203 2975
rect 6837 2941 6871 2975
rect 7389 2941 7423 2975
rect 12516 2941 12550 2975
rect 12909 2941 12943 2975
rect 5318 2873 5352 2907
rect 6193 2873 6227 2907
rect 8538 2873 8572 2907
rect 10149 2873 10183 2907
rect 10701 2873 10735 2907
rect 4813 2805 4847 2839
rect 8033 2805 8067 2839
rect 9137 2805 9171 2839
rect 10977 2805 11011 2839
rect 12587 2805 12621 2839
rect 3525 2601 3559 2635
rect 5089 2601 5123 2635
rect 7849 2601 7883 2635
rect 10425 2601 10459 2635
rect 3893 2533 3927 2567
rect 5457 2533 5491 2567
rect 6377 2533 6411 2567
rect 7205 2533 7239 2567
rect 4169 2465 4203 2499
rect 6929 2465 6963 2499
rect 8493 2465 8527 2499
rect 8744 2465 8778 2499
rect 9137 2465 9171 2499
rect 9781 2465 9815 2499
rect 10885 2465 10919 2499
rect 12700 2465 12734 2499
rect 13093 2465 13127 2499
rect 5365 2397 5399 2431
rect 11437 2397 11471 2431
rect 4813 2329 4847 2363
rect 5917 2329 5951 2363
rect 12771 2329 12805 2363
rect 4353 2261 4387 2295
rect 6653 2261 6687 2295
rect 8125 2261 8159 2295
rect 8815 2261 8849 2295
rect 9965 2261 9999 2295
rect 11069 2261 11103 2295
<< metal1 >>
rect 566 39584 572 39636
rect 624 39624 630 39636
rect 1210 39624 1216 39636
rect 624 39596 1216 39624
rect 624 39584 630 39596
rect 1210 39584 1216 39596
rect 1268 39584 1274 39636
rect 2774 39584 2780 39636
rect 2832 39624 2838 39636
rect 3510 39624 3516 39636
rect 2832 39596 3516 39624
rect 2832 39584 2838 39596
rect 3510 39584 3516 39596
rect 3568 39584 3574 39636
rect 13814 39584 13820 39636
rect 13872 39624 13878 39636
rect 15378 39624 15384 39636
rect 13872 39596 15384 39624
rect 13872 39584 13878 39596
rect 15378 39584 15384 39596
rect 15436 39584 15442 39636
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 10042 35816 10048 35828
rect 10003 35788 10048 35816
rect 10042 35776 10048 35788
rect 10100 35776 10106 35828
rect 5534 35572 5540 35624
rect 5592 35612 5598 35624
rect 6892 35615 6950 35621
rect 6892 35612 6904 35615
rect 5592 35584 6904 35612
rect 5592 35572 5598 35584
rect 6892 35581 6904 35584
rect 6938 35612 6950 35615
rect 7285 35615 7343 35621
rect 7285 35612 7297 35615
rect 6938 35584 7297 35612
rect 6938 35581 6950 35584
rect 6892 35575 6950 35581
rect 7285 35581 7297 35584
rect 7331 35581 7343 35615
rect 7285 35575 7343 35581
rect 8941 35615 8999 35621
rect 8941 35581 8953 35615
rect 8987 35612 8999 35615
rect 9306 35612 9312 35624
rect 8987 35584 9312 35612
rect 8987 35581 8999 35584
rect 8941 35575 8999 35581
rect 9306 35572 9312 35584
rect 9364 35612 9370 35624
rect 9804 35615 9862 35621
rect 9804 35612 9816 35615
rect 9364 35584 9816 35612
rect 9364 35572 9370 35584
rect 9804 35581 9816 35584
rect 9850 35612 9862 35615
rect 10229 35615 10287 35621
rect 10229 35612 10241 35615
rect 9850 35584 10241 35612
rect 9850 35581 9862 35584
rect 9804 35575 9862 35581
rect 10229 35581 10241 35584
rect 10275 35581 10287 35615
rect 10229 35575 10287 35581
rect 5350 35504 5356 35556
rect 5408 35544 5414 35556
rect 6730 35544 6736 35556
rect 5408 35516 6736 35544
rect 5408 35504 5414 35516
rect 6730 35504 6736 35516
rect 6788 35504 6794 35556
rect 8113 35547 8171 35553
rect 8113 35513 8125 35547
rect 8159 35544 8171 35547
rect 8294 35544 8300 35556
rect 8159 35516 8300 35544
rect 8159 35513 8171 35516
rect 8113 35507 8171 35513
rect 8294 35504 8300 35516
rect 8352 35504 8358 35556
rect 8386 35504 8392 35556
rect 8444 35544 8450 35556
rect 8444 35516 8489 35544
rect 8444 35504 8450 35516
rect 6822 35436 6828 35488
rect 6880 35476 6886 35488
rect 6963 35479 7021 35485
rect 6963 35476 6975 35479
rect 6880 35448 6975 35476
rect 6880 35436 6886 35448
rect 6963 35445 6975 35448
rect 7009 35445 7021 35479
rect 6963 35439 7021 35445
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 6822 35272 6828 35284
rect 6783 35244 6828 35272
rect 6822 35232 6828 35244
rect 6880 35232 6886 35284
rect 8294 35232 8300 35284
rect 8352 35272 8358 35284
rect 8481 35275 8539 35281
rect 8481 35272 8493 35275
rect 8352 35244 8493 35272
rect 8352 35232 8358 35244
rect 8481 35241 8493 35244
rect 8527 35241 8539 35275
rect 8481 35235 8539 35241
rect 9861 35275 9919 35281
rect 9861 35241 9873 35275
rect 9907 35272 9919 35275
rect 10502 35272 10508 35284
rect 9907 35244 10508 35272
rect 9907 35241 9919 35244
rect 9861 35235 9919 35241
rect 10502 35232 10508 35244
rect 10560 35232 10566 35284
rect 7006 35164 7012 35216
rect 7064 35204 7070 35216
rect 7101 35207 7159 35213
rect 7101 35204 7113 35207
rect 7064 35176 7113 35204
rect 7064 35164 7070 35176
rect 7101 35173 7113 35176
rect 7147 35173 7159 35207
rect 7101 35167 7159 35173
rect 5956 35139 6014 35145
rect 5956 35105 5968 35139
rect 6002 35136 6014 35139
rect 6178 35136 6184 35148
rect 6002 35108 6184 35136
rect 6002 35105 6014 35108
rect 5956 35099 6014 35105
rect 6178 35096 6184 35108
rect 6236 35096 6242 35148
rect 9674 35136 9680 35148
rect 9635 35108 9680 35136
rect 9674 35096 9680 35108
rect 9732 35096 9738 35148
rect 6043 35071 6101 35077
rect 6043 35037 6055 35071
rect 6089 35068 6101 35071
rect 6457 35071 6515 35077
rect 6457 35068 6469 35071
rect 6089 35040 6469 35068
rect 6089 35037 6101 35040
rect 6043 35031 6101 35037
rect 6457 35037 6469 35040
rect 6503 35068 6515 35071
rect 7009 35071 7067 35077
rect 7009 35068 7021 35071
rect 6503 35040 7021 35068
rect 6503 35037 6515 35040
rect 6457 35031 6515 35037
rect 7009 35037 7021 35040
rect 7055 35037 7067 35071
rect 7009 35031 7067 35037
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35068 7711 35071
rect 9766 35068 9772 35080
rect 7699 35040 9772 35068
rect 7699 35037 7711 35040
rect 7653 35031 7711 35037
rect 9766 35028 9772 35040
rect 9824 35028 9830 35080
rect 8294 34932 8300 34944
rect 8255 34904 8300 34932
rect 8294 34892 8300 34904
rect 8352 34892 8358 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 5534 34728 5540 34740
rect 5495 34700 5540 34728
rect 5534 34688 5540 34700
rect 5592 34688 5598 34740
rect 5718 34688 5724 34740
rect 5776 34728 5782 34740
rect 6178 34728 6184 34740
rect 5776 34700 6184 34728
rect 5776 34688 5782 34700
rect 6178 34688 6184 34700
rect 6236 34688 6242 34740
rect 6730 34688 6736 34740
rect 6788 34728 6794 34740
rect 9674 34728 9680 34740
rect 6788 34700 9680 34728
rect 6788 34688 6794 34700
rect 9674 34688 9680 34700
rect 9732 34688 9738 34740
rect 9950 34688 9956 34740
rect 10008 34728 10014 34740
rect 10229 34731 10287 34737
rect 10229 34728 10241 34731
rect 10008 34700 10241 34728
rect 10008 34688 10014 34700
rect 10229 34697 10241 34700
rect 10275 34697 10287 34731
rect 10229 34691 10287 34697
rect 12621 34731 12679 34737
rect 12621 34697 12633 34731
rect 12667 34728 12679 34731
rect 12802 34728 12808 34740
rect 12667 34700 12808 34728
rect 12667 34697 12679 34700
rect 12621 34691 12679 34697
rect 12802 34688 12808 34700
rect 12860 34688 12866 34740
rect 5813 34663 5871 34669
rect 5813 34629 5825 34663
rect 5859 34660 5871 34663
rect 7098 34660 7104 34672
rect 5859 34632 7104 34660
rect 5859 34629 5871 34632
rect 5813 34623 5871 34629
rect 7098 34620 7104 34632
rect 7156 34620 7162 34672
rect 7558 34660 7564 34672
rect 7519 34632 7564 34660
rect 7558 34620 7564 34632
rect 7616 34660 7622 34672
rect 7616 34632 8616 34660
rect 7616 34620 7622 34632
rect 8588 34604 8616 34632
rect 6822 34552 6828 34604
rect 6880 34592 6886 34604
rect 7009 34595 7067 34601
rect 7009 34592 7021 34595
rect 6880 34564 7021 34592
rect 6880 34552 6886 34564
rect 7009 34561 7021 34564
rect 7055 34561 7067 34595
rect 8570 34592 8576 34604
rect 8483 34564 8576 34592
rect 7009 34555 7067 34561
rect 8570 34552 8576 34564
rect 8628 34552 8634 34604
rect 9217 34595 9275 34601
rect 9217 34561 9229 34595
rect 9263 34592 9275 34595
rect 9306 34592 9312 34604
rect 9263 34564 9312 34592
rect 9263 34561 9275 34564
rect 9217 34555 9275 34561
rect 9306 34552 9312 34564
rect 9364 34552 9370 34604
rect 5534 34484 5540 34536
rect 5592 34524 5598 34536
rect 5629 34527 5687 34533
rect 5629 34524 5641 34527
rect 5592 34496 5641 34524
rect 5592 34484 5598 34496
rect 5629 34493 5641 34496
rect 5675 34524 5687 34527
rect 5994 34524 6000 34536
rect 5675 34496 6000 34524
rect 5675 34493 5687 34496
rect 5629 34487 5687 34493
rect 5994 34484 6000 34496
rect 6052 34484 6058 34536
rect 10042 34524 10048 34536
rect 10003 34496 10048 34524
rect 10042 34484 10048 34496
rect 10100 34524 10106 34536
rect 10597 34527 10655 34533
rect 10597 34524 10609 34527
rect 10100 34496 10609 34524
rect 10100 34484 10106 34496
rect 10597 34493 10609 34496
rect 10643 34493 10655 34527
rect 10597 34487 10655 34493
rect 11238 34484 11244 34536
rect 11296 34524 11302 34536
rect 12437 34527 12495 34533
rect 12437 34524 12449 34527
rect 11296 34496 12449 34524
rect 11296 34484 11302 34496
rect 12437 34493 12449 34496
rect 12483 34524 12495 34527
rect 12989 34527 13047 34533
rect 12989 34524 13001 34527
rect 12483 34496 13001 34524
rect 12483 34493 12495 34496
rect 12437 34487 12495 34493
rect 12989 34493 13001 34496
rect 13035 34493 13047 34527
rect 12989 34487 13047 34493
rect 6641 34459 6699 34465
rect 6641 34425 6653 34459
rect 6687 34456 6699 34459
rect 7006 34456 7012 34468
rect 6687 34428 7012 34456
rect 6687 34425 6699 34428
rect 6641 34419 6699 34425
rect 7006 34416 7012 34428
rect 7064 34456 7070 34468
rect 7101 34459 7159 34465
rect 7101 34456 7113 34459
rect 7064 34428 7113 34456
rect 7064 34416 7070 34428
rect 7101 34425 7113 34428
rect 7147 34425 7159 34459
rect 7101 34419 7159 34425
rect 8662 34416 8668 34468
rect 8720 34456 8726 34468
rect 8720 34428 8765 34456
rect 8720 34416 8726 34428
rect 7926 34388 7932 34400
rect 7887 34360 7932 34388
rect 7926 34348 7932 34360
rect 7984 34348 7990 34400
rect 8389 34391 8447 34397
rect 8389 34357 8401 34391
rect 8435 34388 8447 34391
rect 8680 34388 8708 34416
rect 8435 34360 8708 34388
rect 8435 34357 8447 34360
rect 8389 34351 8447 34357
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 8294 34184 8300 34196
rect 8255 34156 8300 34184
rect 8294 34144 8300 34156
rect 8352 34144 8358 34196
rect 8570 34184 8576 34196
rect 8531 34156 8576 34184
rect 8570 34144 8576 34156
rect 8628 34144 8634 34196
rect 7466 34076 7472 34128
rect 7524 34116 7530 34128
rect 7698 34119 7756 34125
rect 7698 34116 7710 34119
rect 7524 34088 7710 34116
rect 7524 34076 7530 34088
rect 7698 34085 7710 34088
rect 7744 34085 7756 34119
rect 7698 34079 7756 34085
rect 9582 34076 9588 34128
rect 9640 34116 9646 34128
rect 9861 34119 9919 34125
rect 9861 34116 9873 34119
rect 9640 34088 9873 34116
rect 9640 34076 9646 34088
rect 9861 34085 9873 34088
rect 9907 34085 9919 34119
rect 9861 34079 9919 34085
rect 6086 34048 6092 34060
rect 6047 34020 6092 34048
rect 6086 34008 6092 34020
rect 6144 34008 6150 34060
rect 6270 34048 6276 34060
rect 6231 34020 6276 34048
rect 6270 34008 6276 34020
rect 6328 34008 6334 34060
rect 6549 34051 6607 34057
rect 6549 34017 6561 34051
rect 6595 34048 6607 34051
rect 7377 34051 7435 34057
rect 7377 34048 7389 34051
rect 6595 34020 7389 34048
rect 6595 34017 6607 34020
rect 6549 34011 6607 34017
rect 7377 34017 7389 34020
rect 7423 34048 7435 34051
rect 7926 34048 7932 34060
rect 7423 34020 7932 34048
rect 7423 34017 7435 34020
rect 7377 34011 7435 34017
rect 7926 34008 7932 34020
rect 7984 34008 7990 34060
rect 4798 33980 4804 33992
rect 4759 33952 4804 33980
rect 4798 33940 4804 33952
rect 4856 33940 4862 33992
rect 9766 33980 9772 33992
rect 9727 33952 9772 33980
rect 9766 33940 9772 33952
rect 9824 33940 9830 33992
rect 10045 33983 10103 33989
rect 10045 33949 10057 33983
rect 10091 33949 10103 33983
rect 10045 33943 10103 33949
rect 9306 33872 9312 33924
rect 9364 33912 9370 33924
rect 10060 33912 10088 33943
rect 9364 33884 10088 33912
rect 9364 33872 9370 33884
rect 7006 33844 7012 33856
rect 6967 33816 7012 33844
rect 7006 33804 7012 33816
rect 7064 33804 7070 33856
rect 8386 33804 8392 33856
rect 8444 33844 8450 33856
rect 10042 33844 10048 33856
rect 8444 33816 10048 33844
rect 8444 33804 8450 33816
rect 10042 33804 10048 33816
rect 10100 33804 10106 33856
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 6270 33640 6276 33652
rect 4126 33612 6276 33640
rect 4126 33584 4154 33612
rect 6270 33600 6276 33612
rect 6328 33600 6334 33652
rect 7006 33600 7012 33652
rect 7064 33640 7070 33652
rect 7745 33643 7803 33649
rect 7745 33640 7757 33643
rect 7064 33612 7757 33640
rect 7064 33600 7070 33612
rect 7745 33609 7757 33612
rect 7791 33609 7803 33643
rect 7745 33603 7803 33609
rect 8662 33600 8668 33652
rect 8720 33640 8726 33652
rect 9493 33643 9551 33649
rect 9493 33640 9505 33643
rect 8720 33612 9505 33640
rect 8720 33600 8726 33612
rect 9493 33609 9505 33612
rect 9539 33609 9551 33643
rect 9493 33603 9551 33609
rect 9766 33600 9772 33652
rect 9824 33640 9830 33652
rect 10137 33643 10195 33649
rect 10137 33640 10149 33643
rect 9824 33612 10149 33640
rect 9824 33600 9830 33612
rect 10137 33609 10149 33612
rect 10183 33609 10195 33643
rect 10137 33603 10195 33609
rect 4062 33532 4068 33584
rect 4120 33544 4154 33584
rect 4525 33575 4583 33581
rect 4120 33532 4126 33544
rect 4525 33541 4537 33575
rect 4571 33572 4583 33575
rect 4571 33544 5120 33572
rect 4571 33541 4583 33544
rect 4525 33535 4583 33541
rect 3970 33328 3976 33380
rect 4028 33368 4034 33380
rect 4540 33368 4568 33535
rect 5092 33445 5120 33544
rect 9306 33532 9312 33584
rect 9364 33572 9370 33584
rect 9784 33572 9812 33600
rect 9364 33544 9812 33572
rect 9364 33532 9370 33544
rect 6564 33476 7144 33504
rect 6564 33445 6592 33476
rect 4801 33439 4859 33445
rect 4801 33405 4813 33439
rect 4847 33405 4859 33439
rect 4801 33399 4859 33405
rect 5077 33439 5135 33445
rect 5077 33405 5089 33439
rect 5123 33405 5135 33439
rect 6549 33439 6607 33445
rect 6549 33436 6561 33439
rect 5077 33399 5135 33405
rect 5321 33408 6561 33436
rect 4028 33340 4568 33368
rect 4028 33328 4034 33340
rect 4614 33328 4620 33380
rect 4672 33368 4678 33380
rect 4816 33368 4844 33399
rect 4672 33340 4844 33368
rect 4672 33328 4678 33340
rect 4706 33300 4712 33312
rect 4667 33272 4712 33300
rect 4706 33260 4712 33272
rect 4764 33260 4770 33312
rect 4816 33300 4844 33340
rect 4982 33328 4988 33380
rect 5040 33368 5046 33380
rect 5321 33368 5349 33408
rect 6549 33405 6561 33408
rect 6595 33405 6607 33439
rect 6549 33399 6607 33405
rect 6638 33396 6644 33448
rect 6696 33436 6702 33448
rect 6825 33439 6883 33445
rect 6825 33436 6837 33439
rect 6696 33408 6837 33436
rect 6696 33396 6702 33408
rect 6825 33405 6837 33408
rect 6871 33405 6883 33439
rect 7116 33436 7144 33476
rect 8570 33436 8576 33448
rect 7116 33408 7189 33436
rect 8531 33408 8576 33436
rect 6825 33399 6883 33405
rect 5040 33340 5349 33368
rect 5905 33371 5963 33377
rect 5040 33328 5046 33340
rect 5905 33337 5917 33371
rect 5951 33368 5963 33371
rect 6270 33368 6276 33380
rect 5951 33340 6276 33368
rect 5951 33337 5963 33340
rect 5905 33331 5963 33337
rect 6270 33328 6276 33340
rect 6328 33368 6334 33380
rect 6914 33368 6920 33380
rect 6328 33340 6920 33368
rect 6328 33328 6334 33340
rect 6914 33328 6920 33340
rect 6972 33328 6978 33380
rect 7161 33377 7189 33408
rect 8570 33396 8576 33408
rect 8628 33396 8634 33448
rect 7147 33371 7205 33377
rect 7147 33337 7159 33371
rect 7193 33368 7205 33371
rect 7466 33368 7472 33380
rect 7193 33340 7472 33368
rect 7193 33337 7205 33340
rect 7147 33331 7205 33337
rect 7466 33328 7472 33340
rect 7524 33368 7530 33380
rect 8021 33371 8079 33377
rect 8021 33368 8033 33371
rect 7524 33340 8033 33368
rect 7524 33328 7530 33340
rect 8021 33337 8033 33340
rect 8067 33368 8079 33371
rect 8389 33371 8447 33377
rect 8389 33368 8401 33371
rect 8067 33340 8401 33368
rect 8067 33337 8079 33340
rect 8021 33331 8079 33337
rect 8389 33337 8401 33340
rect 8435 33368 8447 33371
rect 8894 33371 8952 33377
rect 8894 33368 8906 33371
rect 8435 33340 8906 33368
rect 8435 33337 8447 33340
rect 8389 33331 8447 33337
rect 8894 33337 8906 33340
rect 8940 33337 8952 33371
rect 8894 33331 8952 33337
rect 6086 33300 6092 33312
rect 4816 33272 6092 33300
rect 6086 33260 6092 33272
rect 6144 33300 6150 33312
rect 6181 33303 6239 33309
rect 6181 33300 6193 33303
rect 6144 33272 6193 33300
rect 6144 33260 6150 33272
rect 6181 33269 6193 33272
rect 6227 33300 6239 33303
rect 8662 33300 8668 33312
rect 6227 33272 8668 33300
rect 6227 33269 6239 33272
rect 6181 33263 6239 33269
rect 8662 33260 8668 33272
rect 8720 33260 8726 33312
rect 9582 33260 9588 33312
rect 9640 33300 9646 33312
rect 9769 33303 9827 33309
rect 9769 33300 9781 33303
rect 9640 33272 9781 33300
rect 9640 33260 9646 33272
rect 9769 33269 9781 33272
rect 9815 33269 9827 33303
rect 9769 33263 9827 33269
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 4614 33096 4620 33108
rect 4575 33068 4620 33096
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 7466 33096 7472 33108
rect 7427 33068 7472 33096
rect 7466 33056 7472 33068
rect 7524 33056 7530 33108
rect 8021 33099 8079 33105
rect 8021 33065 8033 33099
rect 8067 33096 8079 33099
rect 9582 33096 9588 33108
rect 8067 33068 9588 33096
rect 8067 33065 8079 33068
rect 8021 33059 8079 33065
rect 9582 33056 9588 33068
rect 9640 33056 9646 33108
rect 4982 32988 4988 33040
rect 5040 33028 5046 33040
rect 5122 33031 5180 33037
rect 5122 33028 5134 33031
rect 5040 33000 5134 33028
rect 5040 32988 5046 33000
rect 5122 32997 5134 33000
rect 5168 32997 5180 33031
rect 5122 32991 5180 32997
rect 4798 32892 4804 32904
rect 4759 32864 4804 32892
rect 4798 32852 4804 32864
rect 4856 32852 4862 32904
rect 7098 32892 7104 32904
rect 7059 32864 7104 32892
rect 7098 32852 7104 32864
rect 7156 32852 7162 32904
rect 4338 32784 4344 32836
rect 4396 32824 4402 32836
rect 8570 32824 8576 32836
rect 4396 32796 8576 32824
rect 4396 32784 4402 32796
rect 8570 32784 8576 32796
rect 8628 32784 8634 32836
rect 5350 32716 5356 32768
rect 5408 32756 5414 32768
rect 5721 32759 5779 32765
rect 5721 32756 5733 32759
rect 5408 32728 5733 32756
rect 5408 32716 5414 32728
rect 5721 32725 5733 32728
rect 5767 32756 5779 32759
rect 5997 32759 6055 32765
rect 5997 32756 6009 32759
rect 5767 32728 6009 32756
rect 5767 32725 5779 32728
rect 5721 32719 5779 32725
rect 5997 32725 6009 32728
rect 6043 32725 6055 32759
rect 5997 32719 6055 32725
rect 6549 32759 6607 32765
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 6638 32756 6644 32768
rect 6595 32728 6644 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 6638 32716 6644 32728
rect 6696 32716 6702 32768
rect 6914 32756 6920 32768
rect 6875 32728 6920 32756
rect 6914 32716 6920 32728
rect 6972 32716 6978 32768
rect 10042 32756 10048 32768
rect 10003 32728 10048 32756
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 7466 32512 7472 32564
rect 7524 32552 7530 32564
rect 7837 32555 7895 32561
rect 7837 32552 7849 32555
rect 7524 32524 7849 32552
rect 7524 32512 7530 32524
rect 7837 32521 7849 32524
rect 7883 32521 7895 32555
rect 7837 32515 7895 32521
rect 4154 32444 4160 32496
rect 4212 32484 4218 32496
rect 6549 32487 6607 32493
rect 6549 32484 6561 32487
rect 4212 32456 6561 32484
rect 4212 32444 4218 32456
rect 6549 32453 6561 32456
rect 6595 32484 6607 32487
rect 6595 32456 6868 32484
rect 6595 32453 6607 32456
rect 6549 32447 6607 32453
rect 4338 32416 4344 32428
rect 4299 32388 4344 32416
rect 4338 32376 4344 32388
rect 4396 32376 4402 32428
rect 4890 32376 4896 32428
rect 4948 32416 4954 32428
rect 5261 32419 5319 32425
rect 5261 32416 5273 32419
rect 4948 32388 5273 32416
rect 4948 32376 4954 32388
rect 5261 32385 5273 32388
rect 5307 32416 5319 32419
rect 6181 32419 6239 32425
rect 6181 32416 6193 32419
rect 5307 32388 6193 32416
rect 5307 32385 5319 32388
rect 5261 32379 5319 32385
rect 6181 32385 6193 32388
rect 6227 32385 6239 32419
rect 6181 32379 6239 32385
rect 3513 32351 3571 32357
rect 3513 32317 3525 32351
rect 3559 32348 3571 32351
rect 3605 32351 3663 32357
rect 3605 32348 3617 32351
rect 3559 32320 3617 32348
rect 3559 32317 3571 32320
rect 3513 32311 3571 32317
rect 3605 32317 3617 32320
rect 3651 32317 3663 32351
rect 4062 32348 4068 32360
rect 4023 32320 4068 32348
rect 3605 32311 3663 32317
rect 3620 32280 3648 32311
rect 4062 32308 4068 32320
rect 4120 32308 4126 32360
rect 6840 32357 6868 32456
rect 6914 32376 6920 32428
rect 6972 32416 6978 32428
rect 6972 32388 10088 32416
rect 6972 32376 6978 32388
rect 7392 32357 7420 32388
rect 10060 32360 10088 32388
rect 6825 32351 6883 32357
rect 6825 32317 6837 32351
rect 6871 32317 6883 32351
rect 6825 32311 6883 32317
rect 7377 32351 7435 32357
rect 7377 32317 7389 32351
rect 7423 32317 7435 32351
rect 8662 32348 8668 32360
rect 8623 32320 8668 32348
rect 7377 32311 7435 32317
rect 8662 32308 8668 32320
rect 8720 32308 8726 32360
rect 8849 32351 8907 32357
rect 8849 32317 8861 32351
rect 8895 32317 8907 32351
rect 8849 32311 8907 32317
rect 4338 32280 4344 32292
rect 3620 32252 4344 32280
rect 4338 32240 4344 32252
rect 4396 32240 4402 32292
rect 5350 32240 5356 32292
rect 5408 32280 5414 32292
rect 5905 32283 5963 32289
rect 5408 32252 5453 32280
rect 5408 32240 5414 32252
rect 5905 32249 5917 32283
rect 5951 32280 5963 32283
rect 7006 32280 7012 32292
rect 5951 32252 7012 32280
rect 5951 32249 5963 32252
rect 5905 32243 5963 32249
rect 7006 32240 7012 32252
rect 7064 32240 7070 32292
rect 8297 32283 8355 32289
rect 8297 32249 8309 32283
rect 8343 32280 8355 32283
rect 8864 32280 8892 32311
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 9953 32351 10011 32357
rect 9953 32348 9965 32351
rect 9732 32320 9965 32348
rect 9732 32308 9738 32320
rect 9953 32317 9965 32320
rect 9999 32317 10011 32351
rect 9953 32311 10011 32317
rect 10042 32308 10048 32360
rect 10100 32348 10106 32360
rect 10413 32351 10471 32357
rect 10413 32348 10425 32351
rect 10100 32320 10425 32348
rect 10100 32308 10106 32320
rect 10413 32317 10425 32320
rect 10459 32317 10471 32351
rect 10413 32311 10471 32317
rect 10226 32280 10232 32292
rect 8343 32252 10232 32280
rect 8343 32249 8355 32252
rect 8297 32243 8355 32249
rect 10226 32240 10232 32252
rect 10284 32240 10290 32292
rect 4893 32215 4951 32221
rect 4893 32181 4905 32215
rect 4939 32212 4951 32215
rect 4982 32212 4988 32224
rect 4939 32184 4988 32212
rect 4939 32181 4951 32184
rect 4893 32175 4951 32181
rect 4982 32172 4988 32184
rect 5040 32172 5046 32224
rect 6638 32172 6644 32224
rect 6696 32212 6702 32224
rect 6917 32215 6975 32221
rect 6917 32212 6929 32215
rect 6696 32184 6929 32212
rect 6696 32172 6702 32184
rect 6917 32181 6929 32184
rect 6963 32181 6975 32215
rect 8478 32212 8484 32224
rect 8439 32184 8484 32212
rect 6917 32175 6975 32181
rect 8478 32172 8484 32184
rect 8536 32172 8542 32224
rect 9674 32172 9680 32224
rect 9732 32212 9738 32224
rect 9769 32215 9827 32221
rect 9769 32212 9781 32215
rect 9732 32184 9781 32212
rect 9732 32172 9738 32184
rect 9769 32181 9781 32184
rect 9815 32181 9827 32215
rect 10042 32212 10048 32224
rect 10003 32184 10048 32212
rect 9769 32175 9827 32181
rect 10042 32172 10048 32184
rect 10100 32172 10106 32224
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 3418 31968 3424 32020
rect 3476 32008 3482 32020
rect 3697 32011 3755 32017
rect 3697 32008 3709 32011
rect 3476 31980 3709 32008
rect 3476 31968 3482 31980
rect 3697 31977 3709 31980
rect 3743 32008 3755 32011
rect 4062 32008 4068 32020
rect 3743 31980 4068 32008
rect 3743 31977 3755 31980
rect 3697 31971 3755 31977
rect 4062 31968 4068 31980
rect 4120 31968 4126 32020
rect 4798 32008 4804 32020
rect 4759 31980 4804 32008
rect 4798 31968 4804 31980
rect 4856 31968 4862 32020
rect 9766 32008 9772 32020
rect 9727 31980 9772 32008
rect 9766 31968 9772 31980
rect 9824 31968 9830 32020
rect 11379 32011 11437 32017
rect 11379 31977 11391 32011
rect 11425 32008 11437 32011
rect 13998 32008 14004 32020
rect 11425 31980 14004 32008
rect 11425 31977 11437 31980
rect 11379 31971 11437 31977
rect 13998 31968 14004 31980
rect 14056 31968 14062 32020
rect 4982 31900 4988 31952
rect 5040 31940 5046 31952
rect 5306 31943 5364 31949
rect 5306 31940 5318 31943
rect 5040 31912 5318 31940
rect 5040 31900 5046 31912
rect 5306 31909 5318 31912
rect 5352 31909 5364 31943
rect 6914 31940 6920 31952
rect 6875 31912 6920 31940
rect 5306 31903 5364 31909
rect 6914 31900 6920 31912
rect 6972 31900 6978 31952
rect 7098 31900 7104 31952
rect 7156 31940 7162 31952
rect 7837 31943 7895 31949
rect 7837 31940 7849 31943
rect 7156 31912 7849 31940
rect 7156 31900 7162 31912
rect 7837 31909 7849 31912
rect 7883 31940 7895 31943
rect 10042 31940 10048 31952
rect 7883 31912 10048 31940
rect 7883 31909 7895 31912
rect 7837 31903 7895 31909
rect 10042 31900 10048 31912
rect 10100 31900 10106 31952
rect 9674 31872 9680 31884
rect 9635 31844 9680 31872
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10226 31872 10232 31884
rect 10139 31844 10232 31872
rect 10226 31832 10232 31844
rect 10284 31872 10290 31884
rect 10962 31872 10968 31884
rect 10284 31844 10968 31872
rect 10284 31832 10290 31844
rect 10962 31832 10968 31844
rect 11020 31832 11026 31884
rect 11308 31875 11366 31881
rect 11308 31841 11320 31875
rect 11354 31872 11366 31875
rect 11422 31872 11428 31884
rect 11354 31844 11428 31872
rect 11354 31841 11366 31844
rect 11308 31835 11366 31841
rect 11422 31832 11428 31844
rect 11480 31832 11486 31884
rect 4614 31764 4620 31816
rect 4672 31804 4678 31816
rect 4985 31807 5043 31813
rect 4985 31804 4997 31807
rect 4672 31776 4997 31804
rect 4672 31764 4678 31776
rect 4985 31773 4997 31776
rect 5031 31773 5043 31807
rect 6822 31804 6828 31816
rect 6783 31776 6828 31804
rect 4985 31767 5043 31773
rect 6822 31764 6828 31776
rect 6880 31764 6886 31816
rect 7006 31764 7012 31816
rect 7064 31804 7070 31816
rect 7101 31807 7159 31813
rect 7101 31804 7113 31807
rect 7064 31776 7113 31804
rect 7064 31764 7070 31776
rect 7101 31773 7113 31776
rect 7147 31773 7159 31807
rect 7101 31767 7159 31773
rect 5902 31668 5908 31680
rect 5863 31640 5908 31668
rect 5902 31628 5908 31640
rect 5960 31628 5966 31680
rect 8481 31671 8539 31677
rect 8481 31637 8493 31671
rect 8527 31668 8539 31671
rect 8662 31668 8668 31680
rect 8527 31640 8668 31668
rect 8527 31637 8539 31640
rect 8481 31631 8539 31637
rect 8662 31628 8668 31640
rect 8720 31668 8726 31680
rect 9490 31668 9496 31680
rect 8720 31640 9496 31668
rect 8720 31628 8726 31640
rect 9490 31628 9496 31640
rect 9548 31628 9554 31680
rect 10134 31628 10140 31680
rect 10192 31668 10198 31680
rect 10689 31671 10747 31677
rect 10689 31668 10701 31671
rect 10192 31640 10701 31668
rect 10192 31628 10198 31640
rect 10689 31637 10701 31640
rect 10735 31637 10747 31671
rect 10689 31631 10747 31637
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 6822 31464 6828 31476
rect 5684 31436 6828 31464
rect 5684 31424 5690 31436
rect 6822 31424 6828 31436
rect 6880 31464 6886 31476
rect 7377 31467 7435 31473
rect 7377 31464 7389 31467
rect 6880 31436 7389 31464
rect 6880 31424 6886 31436
rect 7377 31433 7389 31436
rect 7423 31433 7435 31467
rect 11422 31464 11428 31476
rect 11383 31436 11428 31464
rect 7377 31427 7435 31433
rect 11422 31424 11428 31436
rect 11480 31424 11486 31476
rect 5813 31399 5871 31405
rect 5813 31365 5825 31399
rect 5859 31396 5871 31399
rect 6914 31396 6920 31408
rect 5859 31368 6920 31396
rect 5859 31365 5871 31368
rect 5813 31359 5871 31365
rect 6914 31356 6920 31368
rect 6972 31396 6978 31408
rect 7009 31399 7067 31405
rect 7009 31396 7021 31399
rect 6972 31368 7021 31396
rect 6972 31356 6978 31368
rect 7009 31365 7021 31368
rect 7055 31365 7067 31399
rect 7009 31359 7067 31365
rect 10410 31356 10416 31408
rect 10468 31396 10474 31408
rect 10689 31399 10747 31405
rect 10689 31396 10701 31399
rect 10468 31368 10701 31396
rect 10468 31356 10474 31368
rect 10689 31365 10701 31368
rect 10735 31396 10747 31399
rect 11440 31396 11468 31424
rect 10735 31368 11468 31396
rect 10735 31365 10747 31368
rect 10689 31359 10747 31365
rect 4801 31331 4859 31337
rect 4801 31297 4813 31331
rect 4847 31328 4859 31331
rect 4982 31328 4988 31340
rect 4847 31300 4988 31328
rect 4847 31297 4859 31300
rect 4801 31291 4859 31297
rect 4982 31288 4988 31300
rect 5040 31288 5046 31340
rect 7837 31331 7895 31337
rect 7837 31297 7849 31331
rect 7883 31328 7895 31331
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 7883 31300 8309 31328
rect 7883 31297 7895 31300
rect 7837 31291 7895 31297
rect 8297 31297 8309 31300
rect 8343 31328 8355 31331
rect 9766 31328 9772 31340
rect 8343 31300 9772 31328
rect 8343 31297 8355 31300
rect 8297 31291 8355 31297
rect 9766 31288 9772 31300
rect 9824 31288 9830 31340
rect 10134 31328 10140 31340
rect 10095 31300 10140 31328
rect 10134 31288 10140 31300
rect 10192 31288 10198 31340
rect 3605 31263 3663 31269
rect 3605 31229 3617 31263
rect 3651 31229 3663 31263
rect 3605 31223 3663 31229
rect 3881 31263 3939 31269
rect 3881 31229 3893 31263
rect 3927 31260 3939 31263
rect 3970 31260 3976 31272
rect 3927 31232 3976 31260
rect 3927 31229 3939 31232
rect 3881 31223 3939 31229
rect 3237 31195 3295 31201
rect 3237 31161 3249 31195
rect 3283 31192 3295 31195
rect 3620 31192 3648 31223
rect 3970 31220 3976 31232
rect 4028 31220 4034 31272
rect 4065 31263 4123 31269
rect 4065 31229 4077 31263
rect 4111 31260 4123 31263
rect 4893 31263 4951 31269
rect 4893 31260 4905 31263
rect 4111 31232 4905 31260
rect 4111 31229 4123 31232
rect 4065 31223 4123 31229
rect 4893 31229 4905 31232
rect 4939 31260 4951 31263
rect 6089 31263 6147 31269
rect 6089 31260 6101 31263
rect 4939 31232 6101 31260
rect 4939 31229 4951 31232
rect 4893 31223 4951 31229
rect 6089 31229 6101 31232
rect 6135 31229 6147 31263
rect 9674 31260 9680 31272
rect 6089 31223 6147 31229
rect 8220 31232 9680 31260
rect 3283 31164 4844 31192
rect 3283 31161 3295 31164
rect 3237 31155 3295 31161
rect 4433 31127 4491 31133
rect 4433 31093 4445 31127
rect 4479 31124 4491 31127
rect 4614 31124 4620 31136
rect 4479 31096 4620 31124
rect 4479 31093 4491 31096
rect 4433 31087 4491 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 4816 31124 4844 31164
rect 4982 31152 4988 31204
rect 5040 31192 5046 31204
rect 5214 31195 5272 31201
rect 5214 31192 5226 31195
rect 5040 31164 5226 31192
rect 5040 31152 5046 31164
rect 5214 31161 5226 31164
rect 5260 31161 5272 31195
rect 8220 31192 8248 31232
rect 9674 31220 9680 31232
rect 9732 31220 9738 31272
rect 5214 31155 5272 31161
rect 5552 31164 8248 31192
rect 8618 31195 8676 31201
rect 5552 31136 5580 31164
rect 8618 31161 8630 31195
rect 8664 31161 8676 31195
rect 8618 31155 8676 31161
rect 5534 31124 5540 31136
rect 4816 31096 5540 31124
rect 5534 31084 5540 31096
rect 5592 31084 5598 31136
rect 8110 31124 8116 31136
rect 8071 31096 8116 31124
rect 8110 31084 8116 31096
rect 8168 31124 8174 31136
rect 8633 31124 8661 31155
rect 10226 31152 10232 31204
rect 10284 31192 10290 31204
rect 10284 31164 10329 31192
rect 10284 31152 10290 31164
rect 8168 31096 8661 31124
rect 9217 31127 9275 31133
rect 8168 31084 8174 31096
rect 9217 31093 9229 31127
rect 9263 31124 9275 31127
rect 9582 31124 9588 31136
rect 9263 31096 9588 31124
rect 9263 31093 9275 31096
rect 9217 31087 9275 31093
rect 9582 31084 9588 31096
rect 9640 31084 9646 31136
rect 10962 31084 10968 31136
rect 11020 31124 11026 31136
rect 11057 31127 11115 31133
rect 11057 31124 11069 31127
rect 11020 31096 11069 31124
rect 11020 31084 11026 31096
rect 11057 31093 11069 31096
rect 11103 31093 11115 31127
rect 11057 31087 11115 31093
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 3421 30923 3479 30929
rect 3421 30889 3433 30923
rect 3467 30920 3479 30923
rect 3970 30920 3976 30932
rect 3467 30892 3976 30920
rect 3467 30889 3479 30892
rect 3421 30883 3479 30889
rect 3970 30880 3976 30892
rect 4028 30880 4034 30932
rect 5368 30892 6224 30920
rect 4246 30812 4252 30864
rect 4304 30852 4310 30864
rect 4479 30855 4537 30861
rect 4479 30852 4491 30855
rect 4304 30824 4491 30852
rect 4304 30812 4310 30824
rect 4479 30821 4491 30824
rect 4525 30821 4537 30855
rect 4479 30815 4537 30821
rect 3970 30744 3976 30796
rect 4028 30784 4034 30796
rect 4392 30787 4450 30793
rect 4392 30784 4404 30787
rect 4028 30756 4404 30784
rect 4028 30744 4034 30756
rect 4392 30753 4404 30756
rect 4438 30784 4450 30787
rect 5368 30784 5396 30892
rect 5629 30855 5687 30861
rect 5629 30821 5641 30855
rect 5675 30852 5687 30855
rect 5902 30852 5908 30864
rect 5675 30824 5908 30852
rect 5675 30821 5687 30824
rect 5629 30815 5687 30821
rect 5902 30812 5908 30824
rect 5960 30812 5966 30864
rect 6196 30861 6224 30892
rect 8110 30880 8116 30932
rect 8168 30920 8174 30932
rect 8205 30923 8263 30929
rect 8205 30920 8217 30923
rect 8168 30892 8217 30920
rect 8168 30880 8174 30892
rect 8205 30889 8217 30892
rect 8251 30889 8263 30923
rect 8205 30883 8263 30889
rect 8757 30923 8815 30929
rect 8757 30889 8769 30923
rect 8803 30920 8815 30923
rect 10226 30920 10232 30932
rect 8803 30892 10232 30920
rect 8803 30889 8815 30892
rect 8757 30883 8815 30889
rect 10226 30880 10232 30892
rect 10284 30920 10290 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10284 30892 10701 30920
rect 10284 30880 10290 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 6181 30855 6239 30861
rect 6181 30821 6193 30855
rect 6227 30852 6239 30855
rect 7006 30852 7012 30864
rect 6227 30824 7012 30852
rect 6227 30821 6239 30824
rect 6181 30815 6239 30821
rect 7006 30812 7012 30824
rect 7064 30812 7070 30864
rect 9858 30852 9864 30864
rect 9819 30824 9864 30852
rect 9858 30812 9864 30824
rect 9916 30812 9922 30864
rect 10410 30852 10416 30864
rect 10371 30824 10416 30852
rect 10410 30812 10416 30824
rect 10468 30812 10474 30864
rect 4438 30756 5396 30784
rect 4438 30753 4450 30756
rect 4392 30747 4450 30753
rect 5350 30676 5356 30728
rect 5408 30716 5414 30728
rect 5537 30719 5595 30725
rect 5537 30716 5549 30719
rect 5408 30688 5549 30716
rect 5408 30676 5414 30688
rect 5537 30685 5549 30688
rect 5583 30685 5595 30719
rect 7834 30716 7840 30728
rect 7795 30688 7840 30716
rect 5537 30679 5595 30685
rect 7834 30676 7840 30688
rect 7892 30676 7898 30728
rect 9766 30716 9772 30728
rect 9679 30688 9772 30716
rect 9766 30676 9772 30688
rect 9824 30716 9830 30728
rect 11241 30719 11299 30725
rect 11241 30716 11253 30719
rect 9824 30688 11253 30716
rect 9824 30676 9830 30688
rect 11241 30685 11253 30688
rect 11287 30685 11299 30719
rect 11241 30679 11299 30685
rect 4982 30580 4988 30592
rect 4943 30552 4988 30580
rect 4982 30540 4988 30552
rect 5040 30540 5046 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 3881 30379 3939 30385
rect 3881 30345 3893 30379
rect 3927 30376 3939 30379
rect 3970 30376 3976 30388
rect 3927 30348 3976 30376
rect 3927 30345 3939 30348
rect 3881 30339 3939 30345
rect 3970 30336 3976 30348
rect 4028 30336 4034 30388
rect 4062 30336 4068 30388
rect 4120 30376 4126 30388
rect 5813 30379 5871 30385
rect 4120 30336 4154 30376
rect 5813 30345 5825 30379
rect 5859 30376 5871 30379
rect 5902 30376 5908 30388
rect 5859 30348 5908 30376
rect 5859 30345 5871 30348
rect 5813 30339 5871 30345
rect 5902 30336 5908 30348
rect 5960 30336 5966 30388
rect 9766 30376 9772 30388
rect 9727 30348 9772 30376
rect 9766 30336 9772 30348
rect 9824 30336 9830 30388
rect 9858 30336 9864 30388
rect 9916 30376 9922 30388
rect 11425 30379 11483 30385
rect 11425 30376 11437 30379
rect 9916 30348 11437 30376
rect 9916 30336 9922 30348
rect 11425 30345 11437 30348
rect 11471 30345 11483 30379
rect 11425 30339 11483 30345
rect 4126 30104 4154 30336
rect 4982 30268 4988 30320
rect 5040 30308 5046 30320
rect 7745 30311 7803 30317
rect 7745 30308 7757 30311
rect 5040 30280 7757 30308
rect 5040 30268 5046 30280
rect 7745 30277 7757 30280
rect 7791 30308 7803 30311
rect 8110 30308 8116 30320
rect 7791 30280 8116 30308
rect 7791 30277 7803 30280
rect 7745 30271 7803 30277
rect 8110 30268 8116 30280
rect 8168 30268 8174 30320
rect 9217 30311 9275 30317
rect 9217 30277 9229 30311
rect 9263 30308 9275 30311
rect 9876 30308 9904 30336
rect 9263 30280 9904 30308
rect 9263 30277 9275 30280
rect 9217 30271 9275 30277
rect 7006 30240 7012 30252
rect 4724 30212 7012 30240
rect 4338 30132 4344 30184
rect 4396 30172 4402 30184
rect 4724 30181 4752 30212
rect 7006 30200 7012 30212
rect 7064 30200 7070 30252
rect 8297 30243 8355 30249
rect 8297 30209 8309 30243
rect 8343 30240 8355 30243
rect 8478 30240 8484 30252
rect 8343 30212 8484 30240
rect 8343 30209 8355 30212
rect 8297 30203 8355 30209
rect 8478 30200 8484 30212
rect 8536 30200 8542 30252
rect 10410 30240 10416 30252
rect 10371 30212 10416 30240
rect 10410 30200 10416 30212
rect 10468 30200 10474 30252
rect 4617 30175 4675 30181
rect 4617 30172 4629 30175
rect 4396 30144 4629 30172
rect 4396 30132 4402 30144
rect 4617 30141 4629 30144
rect 4663 30172 4675 30175
rect 4709 30175 4767 30181
rect 4709 30172 4721 30175
rect 4663 30144 4721 30172
rect 4663 30141 4675 30144
rect 4617 30135 4675 30141
rect 4709 30141 4721 30144
rect 4755 30141 4767 30175
rect 5169 30175 5227 30181
rect 5169 30172 5181 30175
rect 4709 30135 4767 30141
rect 4816 30144 5181 30172
rect 4249 30107 4307 30113
rect 4249 30104 4261 30107
rect 4126 30076 4261 30104
rect 4249 30073 4261 30076
rect 4295 30104 4307 30107
rect 4430 30104 4436 30116
rect 4295 30076 4436 30104
rect 4295 30073 4307 30076
rect 4249 30067 4307 30073
rect 4430 30064 4436 30076
rect 4488 30104 4494 30116
rect 4816 30104 4844 30144
rect 5169 30141 5181 30144
rect 5215 30141 5227 30175
rect 5169 30135 5227 30141
rect 6730 30132 6736 30184
rect 6788 30172 6794 30184
rect 6860 30175 6918 30181
rect 6860 30172 6872 30175
rect 6788 30144 6872 30172
rect 6788 30132 6794 30144
rect 6860 30141 6872 30144
rect 6906 30172 6918 30175
rect 7285 30175 7343 30181
rect 7285 30172 7297 30175
rect 6906 30144 7297 30172
rect 6906 30141 6918 30144
rect 6860 30135 6918 30141
rect 7285 30141 7297 30144
rect 7331 30141 7343 30175
rect 7285 30135 7343 30141
rect 4488 30076 4844 30104
rect 4488 30064 4494 30076
rect 8110 30064 8116 30116
rect 8168 30104 8174 30116
rect 8618 30107 8676 30113
rect 8618 30104 8630 30107
rect 8168 30076 8630 30104
rect 8168 30064 8174 30076
rect 8618 30073 8630 30076
rect 8664 30073 8676 30107
rect 10134 30104 10140 30116
rect 10095 30076 10140 30104
rect 8618 30067 8676 30073
rect 10134 30064 10140 30076
rect 10192 30064 10198 30116
rect 10229 30107 10287 30113
rect 10229 30073 10241 30107
rect 10275 30104 10287 30107
rect 11057 30107 11115 30113
rect 11057 30104 11069 30107
rect 10275 30076 11069 30104
rect 10275 30073 10287 30076
rect 10229 30067 10287 30073
rect 11057 30073 11069 30076
rect 11103 30073 11115 30107
rect 11057 30067 11115 30073
rect 4614 29996 4620 30048
rect 4672 30036 4678 30048
rect 4801 30039 4859 30045
rect 4801 30036 4813 30039
rect 4672 30008 4813 30036
rect 4672 29996 4678 30008
rect 4801 30005 4813 30008
rect 4847 30005 4859 30039
rect 4801 29999 4859 30005
rect 5350 29996 5356 30048
rect 5408 30036 5414 30048
rect 6089 30039 6147 30045
rect 6089 30036 6101 30039
rect 5408 30008 6101 30036
rect 5408 29996 5414 30008
rect 6089 30005 6101 30008
rect 6135 30005 6147 30039
rect 6089 29999 6147 30005
rect 6822 29996 6828 30048
rect 6880 30036 6886 30048
rect 6963 30039 7021 30045
rect 6963 30036 6975 30039
rect 6880 30008 6975 30036
rect 6880 29996 6886 30008
rect 6963 30005 6975 30008
rect 7009 30005 7021 30039
rect 6963 29999 7021 30005
rect 9582 29996 9588 30048
rect 9640 30036 9646 30048
rect 10244 30036 10272 30067
rect 9640 30008 10272 30036
rect 9640 29996 9646 30008
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 4154 29792 4160 29844
rect 4212 29832 4218 29844
rect 8389 29835 8447 29841
rect 4212 29804 4257 29832
rect 4212 29792 4218 29804
rect 8389 29801 8401 29835
rect 8435 29832 8447 29835
rect 8478 29832 8484 29844
rect 8435 29804 8484 29832
rect 8435 29801 8447 29804
rect 8389 29795 8447 29801
rect 8478 29792 8484 29804
rect 8536 29792 8542 29844
rect 9769 29835 9827 29841
rect 9769 29832 9781 29835
rect 8634 29804 9781 29832
rect 6822 29764 6828 29776
rect 6783 29736 6828 29764
rect 6822 29724 6828 29736
rect 6880 29764 6886 29776
rect 7009 29767 7067 29773
rect 7009 29764 7021 29767
rect 6880 29736 7021 29764
rect 6880 29724 6886 29736
rect 7009 29733 7021 29736
rect 7055 29733 7067 29767
rect 7009 29727 7067 29733
rect 7098 29724 7104 29776
rect 7156 29764 7162 29776
rect 7156 29736 7201 29764
rect 7156 29724 7162 29736
rect 7834 29724 7840 29776
rect 7892 29764 7898 29776
rect 8021 29767 8079 29773
rect 8021 29764 8033 29767
rect 7892 29736 8033 29764
rect 7892 29724 7898 29736
rect 8021 29733 8033 29736
rect 8067 29764 8079 29767
rect 8634 29764 8662 29804
rect 9769 29801 9781 29804
rect 9815 29801 9827 29835
rect 9769 29795 9827 29801
rect 10134 29792 10140 29844
rect 10192 29832 10198 29844
rect 10689 29835 10747 29841
rect 10689 29832 10701 29835
rect 10192 29804 10701 29832
rect 10192 29792 10198 29804
rect 10689 29801 10701 29804
rect 10735 29801 10747 29835
rect 10689 29795 10747 29801
rect 8067 29736 8662 29764
rect 8067 29733 8079 29736
rect 8021 29727 8079 29733
rect 4062 29696 4068 29708
rect 4023 29668 4068 29696
rect 4062 29656 4068 29668
rect 4120 29656 4126 29708
rect 4430 29656 4436 29708
rect 4488 29696 4494 29708
rect 4525 29699 4583 29705
rect 4525 29696 4537 29699
rect 4488 29668 4537 29696
rect 4488 29656 4494 29668
rect 4525 29665 4537 29668
rect 4571 29665 4583 29699
rect 4525 29659 4583 29665
rect 4614 29656 4620 29708
rect 4672 29696 4678 29708
rect 5902 29696 5908 29708
rect 5960 29705 5966 29708
rect 5960 29699 5998 29705
rect 4672 29668 5908 29696
rect 4672 29656 4678 29668
rect 5902 29656 5908 29668
rect 5986 29665 5998 29699
rect 5960 29659 5998 29665
rect 8548 29699 8606 29705
rect 8548 29665 8560 29699
rect 8594 29696 8606 29699
rect 8662 29696 8668 29708
rect 8594 29668 8668 29696
rect 8594 29665 8606 29668
rect 8548 29659 8606 29665
rect 5960 29656 5966 29659
rect 8662 29656 8668 29668
rect 8720 29656 8726 29708
rect 9674 29696 9680 29708
rect 9635 29668 9680 29696
rect 9674 29656 9680 29668
rect 9732 29656 9738 29708
rect 9858 29656 9864 29708
rect 9916 29696 9922 29708
rect 10137 29699 10195 29705
rect 10137 29696 10149 29699
rect 9916 29668 10149 29696
rect 9916 29656 9922 29668
rect 10137 29665 10149 29668
rect 10183 29696 10195 29699
rect 10962 29696 10968 29708
rect 10183 29668 10968 29696
rect 10183 29665 10195 29668
rect 10137 29659 10195 29665
rect 10962 29656 10968 29668
rect 11020 29656 11026 29708
rect 7653 29631 7711 29637
rect 7653 29597 7665 29631
rect 7699 29628 7711 29631
rect 9306 29628 9312 29640
rect 7699 29600 9312 29628
rect 7699 29597 7711 29600
rect 7653 29591 7711 29597
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 6043 29495 6101 29501
rect 6043 29461 6055 29495
rect 6089 29492 6101 29495
rect 6914 29492 6920 29504
rect 6089 29464 6920 29492
rect 6089 29461 6101 29464
rect 6043 29455 6101 29461
rect 6914 29452 6920 29464
rect 6972 29452 6978 29504
rect 8478 29452 8484 29504
rect 8536 29492 8542 29504
rect 8619 29495 8677 29501
rect 8619 29492 8631 29495
rect 8536 29464 8631 29492
rect 8536 29452 8542 29464
rect 8619 29461 8631 29464
rect 8665 29492 8677 29495
rect 8941 29495 8999 29501
rect 8941 29492 8953 29495
rect 8665 29464 8953 29492
rect 8665 29461 8677 29464
rect 8619 29455 8677 29461
rect 8941 29461 8953 29464
rect 8987 29461 8999 29495
rect 8941 29455 8999 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 5902 29288 5908 29300
rect 5863 29260 5908 29288
rect 5902 29248 5908 29260
rect 5960 29248 5966 29300
rect 7006 29180 7012 29232
rect 7064 29220 7070 29232
rect 9674 29220 9680 29232
rect 7064 29192 9680 29220
rect 7064 29180 7070 29192
rect 9674 29180 9680 29192
rect 9732 29180 9738 29232
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29152 3387 29155
rect 4154 29152 4160 29164
rect 3375 29124 4160 29152
rect 3375 29121 3387 29124
rect 3329 29115 3387 29121
rect 4154 29112 4160 29124
rect 4212 29152 4218 29164
rect 6914 29152 6920 29164
rect 4212 29124 4257 29152
rect 6875 29124 6920 29152
rect 4212 29112 4218 29124
rect 6914 29112 6920 29124
rect 6972 29112 6978 29164
rect 7558 29152 7564 29164
rect 7519 29124 7564 29152
rect 7558 29112 7564 29124
rect 7616 29152 7622 29164
rect 8294 29152 8300 29164
rect 7616 29124 8300 29152
rect 7616 29112 7622 29124
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 8478 29152 8484 29164
rect 8439 29124 8484 29152
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 9125 29155 9183 29161
rect 9125 29121 9137 29155
rect 9171 29152 9183 29155
rect 9306 29152 9312 29164
rect 9171 29124 9312 29152
rect 9171 29121 9183 29124
rect 9125 29115 9183 29121
rect 9306 29112 9312 29124
rect 9364 29112 9370 29164
rect 4065 29019 4123 29025
rect 4065 28985 4077 29019
rect 4111 29016 4123 29019
rect 4478 29019 4536 29025
rect 4478 29016 4490 29019
rect 4111 28988 4490 29016
rect 4111 28985 4123 28988
rect 4065 28979 4123 28985
rect 4478 28985 4490 28988
rect 4524 29016 4536 29019
rect 4982 29016 4988 29028
rect 4524 28988 4988 29016
rect 4524 28985 4536 28988
rect 4478 28979 4536 28985
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 7009 29019 7067 29025
rect 7009 28985 7021 29019
rect 7055 28985 7067 29019
rect 7009 28979 7067 28985
rect 3697 28951 3755 28957
rect 3697 28917 3709 28951
rect 3743 28948 3755 28951
rect 3878 28948 3884 28960
rect 3743 28920 3884 28948
rect 3743 28917 3755 28920
rect 3697 28911 3755 28917
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 5074 28948 5080 28960
rect 5035 28920 5080 28948
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 6641 28951 6699 28957
rect 6641 28917 6653 28951
rect 6687 28948 6699 28951
rect 7024 28948 7052 28979
rect 8110 28976 8116 29028
rect 8168 29016 8174 29028
rect 8573 29019 8631 29025
rect 8573 29016 8585 29019
rect 8168 28988 8585 29016
rect 8168 28976 8174 28988
rect 8573 28985 8585 28988
rect 8619 28985 8631 29019
rect 8573 28979 8631 28985
rect 7098 28948 7104 28960
rect 6687 28920 7104 28948
rect 6687 28917 6699 28920
rect 6641 28911 6699 28917
rect 7098 28908 7104 28920
rect 7156 28948 7162 28960
rect 7837 28951 7895 28957
rect 7837 28948 7849 28951
rect 7156 28920 7849 28948
rect 7156 28908 7162 28920
rect 7837 28917 7849 28920
rect 7883 28917 7895 28951
rect 7837 28911 7895 28917
rect 8297 28951 8355 28957
rect 8297 28917 8309 28951
rect 8343 28948 8355 28951
rect 8662 28948 8668 28960
rect 8343 28920 8668 28948
rect 8343 28917 8355 28920
rect 8297 28911 8355 28917
rect 8662 28908 8668 28920
rect 8720 28948 8726 28960
rect 9582 28948 9588 28960
rect 8720 28920 9588 28948
rect 8720 28908 8726 28920
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 9858 28908 9864 28960
rect 9916 28948 9922 28960
rect 10045 28951 10103 28957
rect 10045 28948 10057 28951
rect 9916 28920 10057 28948
rect 9916 28908 9922 28920
rect 10045 28917 10057 28920
rect 10091 28917 10103 28951
rect 10045 28911 10103 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 1578 28744 1584 28756
rect 1539 28716 1584 28744
rect 1578 28704 1584 28716
rect 1636 28704 1642 28756
rect 4341 28747 4399 28753
rect 4341 28713 4353 28747
rect 4387 28744 4399 28747
rect 4430 28744 4436 28756
rect 4387 28716 4436 28744
rect 4387 28713 4399 28716
rect 4341 28707 4399 28713
rect 4430 28704 4436 28716
rect 4488 28704 4494 28756
rect 4982 28704 4988 28756
rect 5040 28744 5046 28756
rect 6178 28744 6184 28756
rect 5040 28716 6184 28744
rect 5040 28704 5046 28716
rect 6178 28704 6184 28716
rect 6236 28744 6242 28756
rect 6236 28716 6545 28744
rect 6236 28704 6242 28716
rect 4801 28679 4859 28685
rect 4801 28645 4813 28679
rect 4847 28676 4859 28679
rect 5074 28676 5080 28688
rect 4847 28648 5080 28676
rect 4847 28645 4859 28648
rect 4801 28639 4859 28645
rect 5074 28636 5080 28648
rect 5132 28636 5138 28688
rect 6517 28685 6545 28716
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 7377 28747 7435 28753
rect 7377 28744 7389 28747
rect 6972 28716 7389 28744
rect 6972 28704 6978 28716
rect 7377 28713 7389 28716
rect 7423 28713 7435 28747
rect 7377 28707 7435 28713
rect 6502 28679 6560 28685
rect 6502 28645 6514 28679
rect 6548 28645 6560 28679
rect 8110 28676 8116 28688
rect 8071 28648 8116 28676
rect 6502 28639 6560 28645
rect 8110 28636 8116 28648
rect 8168 28676 8174 28688
rect 8941 28679 8999 28685
rect 8941 28676 8953 28679
rect 8168 28648 8953 28676
rect 8168 28636 8174 28648
rect 8941 28645 8953 28648
rect 8987 28645 8999 28679
rect 8941 28639 8999 28645
rect 1394 28608 1400 28620
rect 1355 28580 1400 28608
rect 1394 28568 1400 28580
rect 1452 28568 1458 28620
rect 2682 28568 2688 28620
rect 2740 28608 2746 28620
rect 2996 28611 3054 28617
rect 2996 28608 3008 28611
rect 2740 28580 3008 28608
rect 2740 28568 2746 28580
rect 2996 28577 3008 28580
rect 3042 28577 3054 28611
rect 7098 28608 7104 28620
rect 7059 28580 7104 28608
rect 2996 28571 3054 28577
rect 3011 28472 3039 28571
rect 7098 28568 7104 28580
rect 7156 28568 7162 28620
rect 9766 28617 9772 28620
rect 9744 28611 9772 28617
rect 9744 28608 9756 28611
rect 9679 28580 9756 28608
rect 9744 28577 9756 28580
rect 9824 28608 9830 28620
rect 11054 28608 11060 28620
rect 9824 28580 11060 28608
rect 9744 28571 9772 28577
rect 9766 28568 9772 28571
rect 9824 28568 9830 28580
rect 11054 28568 11060 28580
rect 11112 28568 11118 28620
rect 3099 28543 3157 28549
rect 3099 28509 3111 28543
rect 3145 28540 3157 28543
rect 4338 28540 4344 28552
rect 3145 28512 4344 28540
rect 3145 28509 3157 28512
rect 3099 28503 3157 28509
rect 4338 28500 4344 28512
rect 4396 28540 4402 28552
rect 4709 28543 4767 28549
rect 4709 28540 4721 28543
rect 4396 28512 4721 28540
rect 4396 28500 4402 28512
rect 4709 28509 4721 28512
rect 4755 28509 4767 28543
rect 5350 28540 5356 28552
rect 5311 28512 5356 28540
rect 4709 28503 4767 28509
rect 5350 28500 5356 28512
rect 5408 28500 5414 28552
rect 6086 28500 6092 28552
rect 6144 28540 6150 28552
rect 6181 28543 6239 28549
rect 6181 28540 6193 28543
rect 6144 28512 6193 28540
rect 6144 28500 6150 28512
rect 6181 28509 6193 28512
rect 6227 28509 6239 28543
rect 8021 28543 8079 28549
rect 8021 28540 8033 28543
rect 6181 28503 6239 28509
rect 7760 28512 8033 28540
rect 6730 28472 6736 28484
rect 3011 28444 6736 28472
rect 6730 28432 6736 28444
rect 6788 28432 6794 28484
rect 7760 28416 7788 28512
rect 8021 28509 8033 28512
rect 8067 28509 8079 28543
rect 8294 28540 8300 28552
rect 8255 28512 8300 28540
rect 8021 28503 8079 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 3970 28364 3976 28416
rect 4028 28404 4034 28416
rect 4430 28404 4436 28416
rect 4028 28376 4436 28404
rect 4028 28364 4034 28376
rect 4430 28364 4436 28376
rect 4488 28364 4494 28416
rect 4982 28364 4988 28416
rect 5040 28404 5046 28416
rect 5629 28407 5687 28413
rect 5629 28404 5641 28407
rect 5040 28376 5641 28404
rect 5040 28364 5046 28376
rect 5629 28373 5641 28376
rect 5675 28373 5687 28407
rect 7742 28404 7748 28416
rect 7703 28376 7748 28404
rect 5629 28367 5687 28373
rect 7742 28364 7748 28376
rect 7800 28364 7806 28416
rect 9815 28407 9873 28413
rect 9815 28373 9827 28407
rect 9861 28404 9873 28407
rect 9950 28404 9956 28416
rect 9861 28376 9956 28404
rect 9861 28373 9873 28376
rect 9815 28367 9873 28373
rect 9950 28364 9956 28376
rect 10008 28404 10014 28416
rect 10137 28407 10195 28413
rect 10137 28404 10149 28407
rect 10008 28376 10149 28404
rect 10008 28364 10014 28376
rect 10137 28373 10149 28376
rect 10183 28373 10195 28407
rect 10137 28367 10195 28373
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 4801 28203 4859 28209
rect 4801 28169 4813 28203
rect 4847 28200 4859 28203
rect 5074 28200 5080 28212
rect 4847 28172 5080 28200
rect 4847 28169 4859 28172
rect 4801 28163 4859 28169
rect 5074 28160 5080 28172
rect 5132 28160 5138 28212
rect 6178 28200 6184 28212
rect 6139 28172 6184 28200
rect 6178 28160 6184 28172
rect 6236 28160 6242 28212
rect 6963 28203 7021 28209
rect 6963 28169 6975 28203
rect 7009 28200 7021 28203
rect 7742 28200 7748 28212
rect 7009 28172 7748 28200
rect 7009 28169 7021 28172
rect 6963 28163 7021 28169
rect 7742 28160 7748 28172
rect 7800 28160 7806 28212
rect 9766 28200 9772 28212
rect 9727 28172 9772 28200
rect 9766 28160 9772 28172
rect 9824 28160 9830 28212
rect 3421 28135 3479 28141
rect 3421 28132 3433 28135
rect 2935 28104 3433 28132
rect 1394 27956 1400 28008
rect 1452 27996 1458 28008
rect 2935 28005 2963 28104
rect 3421 28101 3433 28104
rect 3467 28132 3479 28135
rect 4614 28132 4620 28144
rect 3467 28104 4620 28132
rect 3467 28101 3479 28104
rect 3421 28095 3479 28101
rect 4614 28092 4620 28104
rect 4672 28092 4678 28144
rect 6196 28132 6224 28160
rect 7929 28135 7987 28141
rect 7929 28132 7941 28135
rect 6196 28104 7941 28132
rect 7929 28101 7941 28104
rect 7975 28101 7987 28135
rect 7929 28095 7987 28101
rect 3007 28067 3065 28073
rect 3007 28033 3019 28067
rect 3053 28064 3065 28067
rect 4982 28064 4988 28076
rect 3053 28036 4988 28064
rect 3053 28033 3065 28036
rect 3007 28027 3065 28033
rect 4982 28024 4988 28036
rect 5040 28024 5046 28076
rect 5626 28064 5632 28076
rect 5587 28036 5632 28064
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 1673 27999 1731 28005
rect 1673 27996 1685 27999
rect 1452 27968 1685 27996
rect 1452 27956 1458 27968
rect 1673 27965 1685 27968
rect 1719 27996 1731 27999
rect 2920 27999 2978 28005
rect 2920 27996 2932 27999
rect 1719 27968 2932 27996
rect 1719 27965 1731 27968
rect 1673 27959 1731 27965
rect 2920 27965 2932 27968
rect 2966 27965 2978 27999
rect 2920 27959 2978 27965
rect 3948 27999 4006 28005
rect 3948 27965 3960 27999
rect 3994 27965 4006 27999
rect 3948 27959 4006 27965
rect 6860 27999 6918 28005
rect 6860 27965 6872 27999
rect 6906 27965 6918 27999
rect 6860 27959 6918 27965
rect 2590 27888 2596 27940
rect 2648 27928 2654 27940
rect 3963 27928 3991 27959
rect 4341 27931 4399 27937
rect 4341 27928 4353 27931
rect 2648 27900 4353 27928
rect 2648 27888 2654 27900
rect 4341 27897 4353 27900
rect 4387 27897 4399 27931
rect 4341 27891 4399 27897
rect 3694 27860 3700 27872
rect 3655 27832 3700 27860
rect 3694 27820 3700 27832
rect 3752 27820 3758 27872
rect 4019 27863 4077 27869
rect 4019 27829 4031 27863
rect 4065 27860 4077 27863
rect 4246 27860 4252 27872
rect 4065 27832 4252 27860
rect 4065 27829 4077 27832
rect 4019 27823 4077 27829
rect 4246 27820 4252 27832
rect 4304 27820 4310 27872
rect 4356 27860 4384 27891
rect 5074 27888 5080 27940
rect 5132 27928 5138 27940
rect 5132 27900 5177 27928
rect 5132 27888 5138 27900
rect 6086 27888 6092 27940
rect 6144 27928 6150 27940
rect 6549 27931 6607 27937
rect 6549 27928 6561 27931
rect 6144 27900 6561 27928
rect 6144 27888 6150 27900
rect 6549 27897 6561 27900
rect 6595 27897 6607 27931
rect 6549 27891 6607 27897
rect 6875 27860 6903 27959
rect 7944 27928 7972 28095
rect 9950 28064 9956 28076
rect 9911 28036 9956 28064
rect 9950 28024 9956 28036
rect 10008 28024 10014 28076
rect 10134 28024 10140 28076
rect 10192 28064 10198 28076
rect 10229 28067 10287 28073
rect 10229 28064 10241 28067
rect 10192 28036 10241 28064
rect 10192 28024 10198 28036
rect 10229 28033 10241 28036
rect 10275 28033 10287 28067
rect 10229 28027 10287 28033
rect 8113 27999 8171 28005
rect 8113 27965 8125 27999
rect 8159 27996 8171 27999
rect 8754 27996 8760 28008
rect 8159 27968 8760 27996
rect 8159 27965 8171 27968
rect 8113 27959 8171 27965
rect 8754 27956 8760 27968
rect 8812 27956 8818 28008
rect 8434 27931 8492 27937
rect 8434 27928 8446 27931
rect 7944 27900 8446 27928
rect 8434 27897 8446 27900
rect 8480 27897 8492 27931
rect 9401 27931 9459 27937
rect 9401 27928 9413 27931
rect 8434 27891 8492 27897
rect 9048 27900 9413 27928
rect 9048 27869 9076 27900
rect 9401 27897 9413 27900
rect 9447 27928 9459 27931
rect 10042 27928 10048 27940
rect 9447 27900 10048 27928
rect 9447 27897 9459 27900
rect 9401 27891 9459 27897
rect 10042 27888 10048 27900
rect 10100 27888 10106 27940
rect 7285 27863 7343 27869
rect 7285 27860 7297 27863
rect 4356 27832 7297 27860
rect 7285 27829 7297 27832
rect 7331 27829 7343 27863
rect 7285 27823 7343 27829
rect 9033 27863 9091 27869
rect 9033 27829 9045 27863
rect 9079 27829 9091 27863
rect 9033 27823 9091 27829
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3513 27659 3571 27665
rect 3513 27625 3525 27659
rect 3559 27656 3571 27659
rect 3970 27656 3976 27668
rect 3559 27628 3976 27656
rect 3559 27625 3571 27628
rect 3513 27619 3571 27625
rect 3970 27616 3976 27628
rect 4028 27616 4034 27668
rect 4338 27656 4344 27668
rect 4299 27628 4344 27656
rect 4338 27616 4344 27628
rect 4396 27616 4402 27668
rect 4709 27659 4767 27665
rect 4709 27625 4721 27659
rect 4755 27656 4767 27659
rect 5074 27656 5080 27668
rect 4755 27628 5080 27656
rect 4755 27625 4767 27628
rect 4709 27619 4767 27625
rect 5074 27616 5080 27628
rect 5132 27616 5138 27668
rect 7285 27659 7343 27665
rect 7285 27625 7297 27659
rect 7331 27656 7343 27659
rect 7929 27659 7987 27665
rect 7929 27656 7941 27659
rect 7331 27628 7941 27656
rect 7331 27625 7343 27628
rect 7285 27619 7343 27625
rect 7929 27625 7941 27628
rect 7975 27656 7987 27659
rect 8110 27656 8116 27668
rect 7975 27628 8116 27656
rect 7975 27625 7987 27628
rect 7929 27619 7987 27625
rect 8110 27616 8116 27628
rect 8168 27616 8174 27668
rect 11514 27616 11520 27668
rect 11572 27656 11578 27668
rect 11609 27659 11667 27665
rect 11609 27656 11621 27659
rect 11572 27628 11621 27656
rect 11572 27616 11578 27628
rect 11609 27625 11621 27628
rect 11655 27625 11667 27659
rect 11609 27619 11667 27625
rect 4062 27548 4068 27600
rect 4120 27588 4126 27600
rect 4982 27588 4988 27600
rect 4120 27560 4988 27588
rect 4120 27548 4126 27560
rect 4982 27548 4988 27560
rect 5040 27548 5046 27600
rect 5537 27591 5595 27597
rect 5537 27557 5549 27591
rect 5583 27588 5595 27591
rect 6086 27588 6092 27600
rect 5583 27560 6092 27588
rect 5583 27557 5595 27560
rect 5537 27551 5595 27557
rect 6086 27548 6092 27560
rect 6144 27548 6150 27600
rect 6178 27548 6184 27600
rect 6236 27588 6242 27600
rect 6686 27591 6744 27597
rect 6686 27588 6698 27591
rect 6236 27560 6698 27588
rect 6236 27548 6242 27560
rect 6686 27557 6698 27560
rect 6732 27557 6744 27591
rect 6686 27551 6744 27557
rect 8205 27591 8263 27597
rect 8205 27557 8217 27591
rect 8251 27588 8263 27591
rect 8386 27588 8392 27600
rect 8251 27560 8392 27588
rect 8251 27557 8263 27560
rect 8205 27551 8263 27557
rect 8386 27548 8392 27560
rect 8444 27548 8450 27600
rect 9861 27591 9919 27597
rect 9861 27557 9873 27591
rect 9907 27588 9919 27591
rect 10042 27588 10048 27600
rect 9907 27560 10048 27588
rect 9907 27557 9919 27560
rect 9861 27551 9919 27557
rect 10042 27548 10048 27560
rect 10100 27588 10106 27600
rect 11054 27588 11060 27600
rect 10100 27560 11060 27588
rect 10100 27548 10106 27560
rect 11054 27548 11060 27560
rect 11112 27548 11118 27600
rect 4798 27520 4804 27532
rect 4759 27492 4804 27520
rect 4798 27480 4804 27492
rect 4856 27480 4862 27532
rect 5258 27520 5264 27532
rect 5219 27492 5264 27520
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 11422 27520 11428 27532
rect 11383 27492 11428 27520
rect 11422 27480 11428 27492
rect 11480 27480 11486 27532
rect 4706 27412 4712 27464
rect 4764 27452 4770 27464
rect 6365 27455 6423 27461
rect 6365 27452 6377 27455
rect 4764 27424 6377 27452
rect 4764 27412 4770 27424
rect 6365 27421 6377 27424
rect 6411 27452 6423 27455
rect 7926 27452 7932 27464
rect 6411 27424 7932 27452
rect 6411 27421 6423 27424
rect 6365 27415 6423 27421
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 8435 27455 8493 27461
rect 8435 27421 8447 27455
rect 8481 27452 8493 27455
rect 9398 27452 9404 27464
rect 8481 27424 9404 27452
rect 8481 27421 8493 27424
rect 8435 27415 8493 27421
rect 9398 27412 9404 27424
rect 9456 27452 9462 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9456 27424 9781 27452
rect 9456 27412 9462 27424
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 10226 27452 10232 27464
rect 10187 27424 10232 27452
rect 9769 27415 9827 27421
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 2682 27344 2688 27396
rect 2740 27384 2746 27396
rect 3694 27384 3700 27396
rect 2740 27356 3700 27384
rect 2740 27344 2746 27356
rect 3694 27344 3700 27356
rect 3752 27344 3758 27396
rect 4430 27344 4436 27396
rect 4488 27384 4494 27396
rect 5994 27384 6000 27396
rect 4488 27356 6000 27384
rect 4488 27344 4494 27356
rect 5994 27344 6000 27356
rect 6052 27344 6058 27396
rect 8754 27384 8760 27396
rect 8667 27356 8760 27384
rect 8754 27344 8760 27356
rect 8812 27384 8818 27396
rect 9950 27384 9956 27396
rect 8812 27356 9956 27384
rect 8812 27344 8818 27356
rect 9950 27344 9956 27356
rect 10008 27344 10014 27396
rect 5810 27316 5816 27328
rect 5771 27288 5816 27316
rect 5810 27276 5816 27288
rect 5868 27276 5874 27328
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 9125 27319 9183 27325
rect 9125 27316 9137 27319
rect 8904 27288 9137 27316
rect 8904 27276 8910 27288
rect 9125 27285 9137 27288
rect 9171 27285 9183 27319
rect 9125 27279 9183 27285
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 3142 27072 3148 27124
rect 3200 27112 3206 27124
rect 4430 27112 4436 27124
rect 3200 27084 4436 27112
rect 3200 27072 3206 27084
rect 4430 27072 4436 27084
rect 4488 27072 4494 27124
rect 4525 27115 4583 27121
rect 4525 27081 4537 27115
rect 4571 27112 4583 27115
rect 5258 27112 5264 27124
rect 4571 27084 5264 27112
rect 4571 27081 4583 27084
rect 4525 27075 4583 27081
rect 3418 27004 3424 27056
rect 3476 27044 3482 27056
rect 4540 27044 4568 27075
rect 5258 27072 5264 27084
rect 5316 27072 5322 27124
rect 5442 27072 5448 27124
rect 5500 27112 5506 27124
rect 6178 27112 6184 27124
rect 5500 27084 6184 27112
rect 5500 27072 5506 27084
rect 6178 27072 6184 27084
rect 6236 27112 6242 27124
rect 6365 27115 6423 27121
rect 6365 27112 6377 27115
rect 6236 27084 6377 27112
rect 6236 27072 6242 27084
rect 6365 27081 6377 27084
rect 6411 27081 6423 27115
rect 7926 27112 7932 27124
rect 7887 27084 7932 27112
rect 6365 27075 6423 27081
rect 7926 27072 7932 27084
rect 7984 27072 7990 27124
rect 8386 27112 8392 27124
rect 8347 27084 8392 27112
rect 8386 27072 8392 27084
rect 8444 27072 8450 27124
rect 11054 27112 11060 27124
rect 11015 27084 11060 27112
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 3476 27016 4568 27044
rect 3476 27004 3482 27016
rect 4798 27004 4804 27056
rect 4856 27044 4862 27056
rect 4893 27047 4951 27053
rect 4893 27044 4905 27047
rect 4856 27016 4905 27044
rect 4856 27004 4862 27016
rect 4893 27013 4905 27016
rect 4939 27044 4951 27047
rect 4939 27016 6132 27044
rect 4939 27013 4951 27016
rect 4893 27007 4951 27013
rect 4246 26936 4252 26988
rect 4304 26976 4310 26988
rect 5077 26979 5135 26985
rect 5077 26976 5089 26979
rect 4304 26948 5089 26976
rect 4304 26936 4310 26948
rect 5077 26945 5089 26948
rect 5123 26976 5135 26979
rect 5810 26976 5816 26988
rect 5123 26948 5816 26976
rect 5123 26945 5135 26948
rect 5077 26939 5135 26945
rect 5810 26936 5816 26948
rect 5868 26936 5874 26988
rect 6104 26976 6132 27016
rect 7742 27004 7748 27056
rect 7800 27044 7806 27056
rect 8404 27044 8432 27072
rect 9309 27047 9367 27053
rect 9309 27044 9321 27047
rect 7800 27016 8432 27044
rect 8496 27016 9321 27044
rect 7800 27004 7806 27016
rect 8496 26976 8524 27016
rect 9309 27013 9321 27016
rect 9355 27013 9367 27047
rect 9309 27007 9367 27013
rect 6104 26948 8524 26976
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26976 8631 26979
rect 8846 26976 8852 26988
rect 8619 26948 8852 26976
rect 8619 26945 8631 26948
rect 8573 26939 8631 26945
rect 8846 26936 8852 26948
rect 8904 26936 8910 26988
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26976 9275 26979
rect 10226 26976 10232 26988
rect 9263 26948 10232 26976
rect 9263 26945 9275 26948
rect 9217 26939 9275 26945
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 3697 26911 3755 26917
rect 3697 26877 3709 26911
rect 3743 26877 3755 26911
rect 3970 26908 3976 26920
rect 3931 26880 3976 26908
rect 3697 26871 3755 26877
rect 3329 26843 3387 26849
rect 3329 26809 3341 26843
rect 3375 26840 3387 26843
rect 3712 26840 3740 26871
rect 3970 26868 3976 26880
rect 4028 26868 4034 26920
rect 6914 26908 6920 26920
rect 6875 26880 6920 26908
rect 6914 26868 6920 26880
rect 6972 26868 6978 26920
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26877 7435 26911
rect 7377 26871 7435 26877
rect 9309 26911 9367 26917
rect 9309 26877 9321 26911
rect 9355 26908 9367 26911
rect 9953 26911 10011 26917
rect 9953 26908 9965 26911
rect 9355 26880 9965 26908
rect 9355 26877 9367 26880
rect 9309 26871 9367 26877
rect 9953 26877 9965 26880
rect 9999 26908 10011 26911
rect 10045 26911 10103 26917
rect 10045 26908 10057 26911
rect 9999 26880 10057 26908
rect 9999 26877 10011 26880
rect 9953 26871 10011 26877
rect 10045 26877 10057 26880
rect 10091 26877 10103 26911
rect 10045 26871 10103 26877
rect 10505 26911 10563 26917
rect 10505 26877 10517 26911
rect 10551 26877 10563 26911
rect 10505 26871 10563 26877
rect 3375 26812 3740 26840
rect 3375 26809 3387 26812
rect 3329 26803 3387 26809
rect 3712 26772 3740 26812
rect 4157 26843 4215 26849
rect 4157 26809 4169 26843
rect 4203 26840 4215 26843
rect 4338 26840 4344 26852
rect 4203 26812 4344 26840
rect 4203 26809 4215 26812
rect 4157 26803 4215 26809
rect 4338 26800 4344 26812
rect 4396 26800 4402 26852
rect 5166 26800 5172 26852
rect 5224 26840 5230 26852
rect 5224 26812 5269 26840
rect 5224 26800 5230 26812
rect 5350 26800 5356 26852
rect 5408 26840 5414 26852
rect 5721 26843 5779 26849
rect 5721 26840 5733 26843
rect 5408 26812 5733 26840
rect 5408 26800 5414 26812
rect 5721 26809 5733 26812
rect 5767 26840 5779 26843
rect 6638 26840 6644 26852
rect 5767 26812 6644 26840
rect 5767 26809 5779 26812
rect 5721 26803 5779 26809
rect 6638 26800 6644 26812
rect 6696 26800 6702 26852
rect 4798 26772 4804 26784
rect 3712 26744 4804 26772
rect 4798 26732 4804 26744
rect 4856 26732 4862 26784
rect 5258 26732 5264 26784
rect 5316 26772 5322 26784
rect 5994 26772 6000 26784
rect 5316 26744 6000 26772
rect 5316 26732 5322 26744
rect 5994 26732 6000 26744
rect 6052 26772 6058 26784
rect 7392 26772 7420 26871
rect 7650 26840 7656 26852
rect 7611 26812 7656 26840
rect 7650 26800 7656 26812
rect 7708 26800 7714 26852
rect 8662 26840 8668 26852
rect 8623 26812 8668 26840
rect 8662 26800 8668 26812
rect 8720 26800 8726 26852
rect 9858 26840 9864 26852
rect 9508 26812 9864 26840
rect 9508 26781 9536 26812
rect 9858 26800 9864 26812
rect 9916 26840 9922 26852
rect 10520 26840 10548 26871
rect 9916 26812 10548 26840
rect 9916 26800 9922 26812
rect 9493 26775 9551 26781
rect 9493 26772 9505 26775
rect 6052 26744 9505 26772
rect 6052 26732 6058 26744
rect 9493 26741 9505 26744
rect 9539 26741 9551 26775
rect 9493 26735 9551 26741
rect 9950 26732 9956 26784
rect 10008 26772 10014 26784
rect 10137 26775 10195 26781
rect 10137 26772 10149 26775
rect 10008 26744 10149 26772
rect 10008 26732 10014 26744
rect 10137 26741 10149 26744
rect 10183 26741 10195 26775
rect 11422 26772 11428 26784
rect 11383 26744 11428 26772
rect 10137 26735 10195 26741
rect 11422 26732 11428 26744
rect 11480 26732 11486 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 3418 26568 3424 26580
rect 3379 26540 3424 26568
rect 3418 26528 3424 26540
rect 3476 26568 3482 26580
rect 3970 26568 3976 26580
rect 3476 26540 3976 26568
rect 3476 26528 3482 26540
rect 3970 26528 3976 26540
rect 4028 26528 4034 26580
rect 4246 26528 4252 26580
rect 4304 26568 4310 26580
rect 6914 26568 6920 26580
rect 4304 26540 6920 26568
rect 4304 26528 4310 26540
rect 6914 26528 6920 26540
rect 6972 26568 6978 26580
rect 7101 26571 7159 26577
rect 7101 26568 7113 26571
rect 6972 26540 7113 26568
rect 6972 26528 6978 26540
rect 7101 26537 7113 26540
rect 7147 26537 7159 26571
rect 7101 26531 7159 26537
rect 8662 26528 8668 26580
rect 8720 26568 8726 26580
rect 8757 26571 8815 26577
rect 8757 26568 8769 26571
rect 8720 26540 8769 26568
rect 8720 26528 8726 26540
rect 8757 26537 8769 26540
rect 8803 26568 8815 26571
rect 9033 26571 9091 26577
rect 9033 26568 9045 26571
rect 8803 26540 9045 26568
rect 8803 26537 8815 26540
rect 8757 26531 8815 26537
rect 9033 26537 9045 26540
rect 9079 26537 9091 26571
rect 9398 26568 9404 26580
rect 9359 26540 9404 26568
rect 9033 26531 9091 26537
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 4522 26460 4528 26512
rect 4580 26500 4586 26512
rect 4703 26503 4761 26509
rect 4703 26500 4715 26503
rect 4580 26472 4715 26500
rect 4580 26460 4586 26472
rect 4703 26469 4715 26472
rect 4749 26500 4761 26503
rect 5442 26500 5448 26512
rect 4749 26472 5448 26500
rect 4749 26469 4761 26472
rect 4703 26463 4761 26469
rect 5442 26460 5448 26472
rect 5500 26460 5506 26512
rect 6270 26500 6276 26512
rect 6231 26472 6276 26500
rect 6270 26460 6276 26472
rect 6328 26460 6334 26512
rect 7926 26460 7932 26512
rect 7984 26500 7990 26512
rect 8158 26503 8216 26509
rect 8158 26500 8170 26503
rect 7984 26472 8170 26500
rect 7984 26460 7990 26472
rect 8158 26469 8170 26472
rect 8204 26469 8216 26503
rect 9858 26500 9864 26512
rect 9819 26472 9864 26500
rect 8158 26463 8216 26469
rect 9858 26460 9864 26472
rect 9916 26460 9922 26512
rect 10226 26460 10232 26512
rect 10284 26500 10290 26512
rect 10413 26503 10471 26509
rect 10413 26500 10425 26503
rect 10284 26472 10425 26500
rect 10284 26460 10290 26472
rect 10413 26469 10425 26472
rect 10459 26469 10471 26503
rect 11422 26500 11428 26512
rect 10413 26463 10471 26469
rect 11307 26472 11428 26500
rect 1949 26435 2007 26441
rect 1949 26401 1961 26435
rect 1995 26432 2007 26435
rect 2038 26432 2044 26444
rect 1995 26404 2044 26432
rect 1995 26401 2007 26404
rect 1949 26395 2007 26401
rect 2038 26392 2044 26404
rect 2096 26392 2102 26444
rect 2961 26435 3019 26441
rect 2961 26401 2973 26435
rect 3007 26432 3019 26435
rect 3050 26432 3056 26444
rect 3007 26404 3056 26432
rect 3007 26401 3019 26404
rect 2961 26395 3019 26401
rect 3050 26392 3056 26404
rect 3108 26392 3114 26444
rect 11307 26441 11335 26472
rect 11422 26460 11428 26472
rect 11480 26460 11486 26512
rect 11292 26435 11350 26441
rect 11292 26401 11304 26435
rect 11338 26401 11350 26435
rect 11292 26395 11350 26401
rect 4338 26364 4344 26376
rect 4299 26336 4344 26364
rect 4338 26324 4344 26336
rect 4396 26324 4402 26376
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6638 26364 6644 26376
rect 6599 26336 6644 26364
rect 6181 26327 6239 26333
rect 2087 26299 2145 26305
rect 2087 26265 2099 26299
rect 2133 26296 2145 26299
rect 6196 26296 6224 26327
rect 6638 26324 6644 26336
rect 6696 26324 6702 26376
rect 7834 26364 7840 26376
rect 7795 26336 7840 26364
rect 7834 26324 7840 26336
rect 7892 26324 7898 26376
rect 9769 26367 9827 26373
rect 9769 26333 9781 26367
rect 9815 26364 9827 26367
rect 10870 26364 10876 26376
rect 9815 26336 10876 26364
rect 9815 26333 9827 26336
rect 9769 26327 9827 26333
rect 10870 26324 10876 26336
rect 10928 26364 10934 26376
rect 11379 26367 11437 26373
rect 11379 26364 11391 26367
rect 10928 26336 11391 26364
rect 10928 26324 10934 26336
rect 11379 26333 11391 26336
rect 11425 26333 11437 26367
rect 11379 26327 11437 26333
rect 6454 26296 6460 26308
rect 2133 26268 6460 26296
rect 2133 26265 2145 26268
rect 2087 26259 2145 26265
rect 6454 26256 6460 26268
rect 6512 26256 6518 26308
rect 3099 26231 3157 26237
rect 3099 26197 3111 26231
rect 3145 26228 3157 26231
rect 3326 26228 3332 26240
rect 3145 26200 3332 26228
rect 3145 26197 3157 26200
rect 3099 26191 3157 26197
rect 3326 26188 3332 26200
rect 3384 26188 3390 26240
rect 5166 26188 5172 26240
rect 5224 26228 5230 26240
rect 5261 26231 5319 26237
rect 5261 26228 5273 26231
rect 5224 26200 5273 26228
rect 5224 26188 5230 26200
rect 5261 26197 5273 26200
rect 5307 26228 5319 26231
rect 5537 26231 5595 26237
rect 5537 26228 5549 26231
rect 5307 26200 5549 26228
rect 5307 26197 5319 26200
rect 5261 26191 5319 26197
rect 5537 26197 5549 26200
rect 5583 26197 5595 26231
rect 5537 26191 5595 26197
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 2593 26027 2651 26033
rect 2593 25993 2605 26027
rect 2639 26024 2651 26027
rect 4522 26024 4528 26036
rect 2639 25996 4451 26024
rect 4483 25996 4528 26024
rect 2639 25993 2651 25996
rect 2593 25987 2651 25993
rect 2038 25956 2044 25968
rect 1951 25928 2044 25956
rect 2038 25916 2044 25928
rect 2096 25956 2102 25968
rect 4249 25959 4307 25965
rect 4249 25956 4261 25959
rect 2096 25928 4261 25956
rect 2096 25916 2102 25928
rect 4249 25925 4261 25928
rect 4295 25925 4307 25959
rect 4423 25956 4451 25996
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 4614 25984 4620 26036
rect 4672 26024 4678 26036
rect 5718 26024 5724 26036
rect 4672 25996 5724 26024
rect 4672 25984 4678 25996
rect 5718 25984 5724 25996
rect 5776 25984 5782 26036
rect 6181 26027 6239 26033
rect 6181 25993 6193 26027
rect 6227 26024 6239 26027
rect 6270 26024 6276 26036
rect 6227 25996 6276 26024
rect 6227 25993 6239 25996
rect 6181 25987 6239 25993
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 6454 26024 6460 26036
rect 6415 25996 6460 26024
rect 6454 25984 6460 25996
rect 6512 25984 6518 26036
rect 8662 25984 8668 26036
rect 8720 26024 8726 26036
rect 9677 26027 9735 26033
rect 9677 26024 9689 26027
rect 8720 25996 9689 26024
rect 8720 25984 8726 25996
rect 9677 25993 9689 25996
rect 9723 26024 9735 26027
rect 10042 26024 10048 26036
rect 9723 25996 10048 26024
rect 9723 25993 9735 25996
rect 9677 25987 9735 25993
rect 10042 25984 10048 25996
rect 10100 25984 10106 26036
rect 10870 26024 10876 26036
rect 10831 25996 10876 26024
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 5258 25956 5264 25968
rect 4423 25928 5264 25956
rect 4249 25919 4307 25925
rect 5258 25916 5264 25928
rect 5316 25916 5322 25968
rect 5626 25956 5632 25968
rect 5587 25928 5632 25956
rect 5626 25916 5632 25928
rect 5684 25916 5690 25968
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 2958 25888 2964 25900
rect 1820 25860 2964 25888
rect 1820 25848 1826 25860
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 3326 25848 3332 25900
rect 3384 25888 3390 25900
rect 3384 25860 4936 25888
rect 3384 25848 3390 25860
rect 2406 25820 2412 25832
rect 2367 25792 2412 25820
rect 2406 25780 2412 25792
rect 2464 25780 2470 25832
rect 3697 25823 3755 25829
rect 3697 25789 3709 25823
rect 3743 25789 3755 25823
rect 3878 25820 3884 25832
rect 3839 25792 3884 25820
rect 3697 25783 3755 25789
rect 3712 25752 3740 25783
rect 3878 25780 3884 25792
rect 3936 25780 3942 25832
rect 4157 25823 4215 25829
rect 4157 25789 4169 25823
rect 4203 25820 4215 25823
rect 4706 25820 4712 25832
rect 4203 25792 4712 25820
rect 4203 25789 4215 25792
rect 4157 25783 4215 25789
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 3970 25752 3976 25764
rect 3712 25724 3976 25752
rect 3970 25712 3976 25724
rect 4028 25752 4034 25764
rect 4908 25752 4936 25860
rect 7650 25848 7656 25900
rect 7708 25888 7714 25900
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7708 25860 8125 25888
rect 7708 25848 7714 25860
rect 8113 25857 8125 25860
rect 8159 25888 8171 25891
rect 8938 25888 8944 25900
rect 8159 25860 8944 25888
rect 8159 25857 8171 25860
rect 8113 25851 8171 25857
rect 8938 25848 8944 25860
rect 8996 25848 9002 25900
rect 10134 25848 10140 25900
rect 10192 25888 10198 25900
rect 10229 25891 10287 25897
rect 10229 25888 10241 25891
rect 10192 25860 10241 25888
rect 10192 25848 10198 25860
rect 10229 25857 10241 25860
rect 10275 25857 10287 25891
rect 10229 25851 10287 25857
rect 5810 25780 5816 25832
rect 5868 25820 5874 25832
rect 6860 25823 6918 25829
rect 6860 25820 6872 25823
rect 5868 25792 6872 25820
rect 5868 25780 5874 25792
rect 6860 25789 6872 25792
rect 6906 25820 6918 25823
rect 7285 25823 7343 25829
rect 7285 25820 7297 25823
rect 6906 25792 7297 25820
rect 6906 25789 6918 25792
rect 6860 25783 6918 25789
rect 7285 25789 7297 25792
rect 7331 25789 7343 25823
rect 7285 25783 7343 25789
rect 5074 25752 5080 25764
rect 4028 25724 4154 25752
rect 4908 25724 5080 25752
rect 4028 25712 4034 25724
rect 3050 25684 3056 25696
rect 3011 25656 3056 25684
rect 3050 25644 3056 25656
rect 3108 25644 3114 25696
rect 4126 25684 4154 25724
rect 5074 25712 5080 25724
rect 5132 25712 5138 25764
rect 5166 25712 5172 25764
rect 5224 25752 5230 25764
rect 8434 25755 8492 25761
rect 5224 25724 5269 25752
rect 5224 25712 5230 25724
rect 8434 25721 8446 25755
rect 8480 25721 8492 25755
rect 9950 25752 9956 25764
rect 9911 25724 9956 25752
rect 8434 25715 8492 25721
rect 4246 25684 4252 25696
rect 4126 25656 4252 25684
rect 4246 25644 4252 25656
rect 4304 25644 4310 25696
rect 4341 25687 4399 25693
rect 4341 25653 4353 25687
rect 4387 25684 4399 25687
rect 4706 25684 4712 25696
rect 4387 25656 4712 25684
rect 4387 25653 4399 25656
rect 4341 25647 4399 25653
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 4893 25687 4951 25693
rect 4893 25653 4905 25687
rect 4939 25684 4951 25687
rect 5184 25684 5212 25712
rect 4939 25656 5212 25684
rect 6963 25687 7021 25693
rect 4939 25653 4951 25656
rect 4893 25647 4951 25653
rect 6963 25653 6975 25687
rect 7009 25684 7021 25687
rect 7190 25684 7196 25696
rect 7009 25656 7196 25684
rect 7009 25653 7021 25656
rect 6963 25647 7021 25653
rect 7190 25644 7196 25656
rect 7248 25644 7254 25696
rect 7926 25684 7932 25696
rect 7887 25656 7932 25684
rect 7926 25644 7932 25656
rect 7984 25684 7990 25696
rect 8449 25684 8477 25715
rect 9950 25712 9956 25724
rect 10008 25712 10014 25764
rect 10042 25712 10048 25764
rect 10100 25752 10106 25764
rect 10100 25724 10145 25752
rect 10100 25712 10106 25724
rect 7984 25656 8477 25684
rect 9033 25687 9091 25693
rect 7984 25644 7990 25656
rect 9033 25653 9045 25687
rect 9079 25684 9091 25687
rect 9398 25684 9404 25696
rect 9079 25656 9404 25684
rect 9079 25653 9091 25656
rect 9033 25647 9091 25653
rect 9398 25644 9404 25656
rect 9456 25644 9462 25696
rect 11333 25687 11391 25693
rect 11333 25653 11345 25687
rect 11379 25684 11391 25687
rect 11422 25684 11428 25696
rect 11379 25656 11428 25684
rect 11379 25653 11391 25656
rect 11333 25647 11391 25653
rect 11422 25644 11428 25656
rect 11480 25684 11486 25696
rect 12158 25684 12164 25696
rect 11480 25656 12164 25684
rect 11480 25644 11486 25656
rect 12158 25644 12164 25656
rect 12216 25644 12222 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 3145 25483 3203 25489
rect 3145 25449 3157 25483
rect 3191 25480 3203 25483
rect 3878 25480 3884 25492
rect 3191 25452 3884 25480
rect 3191 25449 3203 25452
rect 3145 25443 3203 25449
rect 3878 25440 3884 25452
rect 3936 25440 3942 25492
rect 4338 25480 4344 25492
rect 4299 25452 4344 25480
rect 4338 25440 4344 25452
rect 4396 25440 4402 25492
rect 5074 25440 5080 25492
rect 5132 25480 5138 25492
rect 5813 25483 5871 25489
rect 5813 25480 5825 25483
rect 5132 25452 5825 25480
rect 5132 25440 5138 25452
rect 5813 25449 5825 25452
rect 5859 25449 5871 25483
rect 5813 25443 5871 25449
rect 8619 25483 8677 25489
rect 8619 25449 8631 25483
rect 8665 25480 8677 25483
rect 8846 25480 8852 25492
rect 8665 25452 8852 25480
rect 8665 25449 8677 25452
rect 8619 25443 8677 25449
rect 8846 25440 8852 25452
rect 8904 25440 8910 25492
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 8996 25452 9041 25480
rect 8996 25440 9002 25452
rect 9950 25440 9956 25492
rect 10008 25480 10014 25492
rect 10689 25483 10747 25489
rect 10689 25480 10701 25483
rect 10008 25452 10701 25480
rect 10008 25440 10014 25452
rect 10689 25449 10701 25452
rect 10735 25480 10747 25483
rect 11379 25483 11437 25489
rect 11379 25480 11391 25483
rect 10735 25452 11391 25480
rect 10735 25449 10747 25452
rect 10689 25443 10747 25449
rect 11379 25449 11391 25452
rect 11425 25449 11437 25483
rect 11379 25443 11437 25449
rect 4522 25372 4528 25424
rect 4580 25412 4586 25424
rect 4938 25415 4996 25421
rect 4938 25412 4950 25415
rect 4580 25384 4950 25412
rect 4580 25372 4586 25384
rect 4938 25381 4950 25384
rect 4984 25381 4996 25415
rect 4938 25375 4996 25381
rect 7653 25415 7711 25421
rect 7653 25381 7665 25415
rect 7699 25412 7711 25415
rect 7834 25412 7840 25424
rect 7699 25384 7840 25412
rect 7699 25381 7711 25384
rect 7653 25375 7711 25381
rect 7834 25372 7840 25384
rect 7892 25412 7898 25424
rect 8297 25415 8355 25421
rect 8297 25412 8309 25415
rect 7892 25384 8309 25412
rect 7892 25372 7898 25384
rect 8297 25381 8309 25384
rect 8343 25381 8355 25415
rect 8297 25375 8355 25381
rect 9398 25372 9404 25424
rect 9456 25412 9462 25424
rect 9858 25412 9864 25424
rect 9456 25384 9864 25412
rect 9456 25372 9462 25384
rect 9858 25372 9864 25384
rect 9916 25412 9922 25424
rect 10410 25412 10416 25424
rect 9916 25384 10416 25412
rect 9916 25372 9922 25384
rect 10410 25372 10416 25384
rect 10468 25372 10474 25424
rect 2961 25347 3019 25353
rect 2961 25313 2973 25347
rect 3007 25344 3019 25347
rect 3234 25344 3240 25356
rect 3007 25316 3240 25344
rect 3007 25313 3019 25316
rect 2961 25307 3019 25313
rect 3234 25304 3240 25316
rect 3292 25304 3298 25356
rect 5258 25304 5264 25356
rect 5316 25344 5322 25356
rect 5537 25347 5595 25353
rect 5537 25344 5549 25347
rect 5316 25316 5549 25344
rect 5316 25304 5322 25316
rect 5537 25313 5549 25316
rect 5583 25344 5595 25347
rect 6178 25344 6184 25356
rect 5583 25316 6184 25344
rect 5583 25313 5595 25316
rect 5537 25307 5595 25313
rect 6178 25304 6184 25316
rect 6236 25304 6242 25356
rect 6914 25344 6920 25356
rect 6875 25316 6920 25344
rect 6914 25304 6920 25316
rect 6972 25304 6978 25356
rect 7377 25347 7435 25353
rect 7377 25313 7389 25347
rect 7423 25313 7435 25347
rect 7377 25307 7435 25313
rect 3513 25279 3571 25285
rect 3513 25245 3525 25279
rect 3559 25276 3571 25279
rect 3970 25276 3976 25288
rect 3559 25248 3976 25276
rect 3559 25245 3571 25248
rect 3513 25239 3571 25245
rect 3970 25236 3976 25248
rect 4028 25236 4034 25288
rect 4614 25276 4620 25288
rect 4575 25248 4620 25276
rect 4614 25236 4620 25248
rect 4672 25236 4678 25288
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 4764 25248 5028 25276
rect 4764 25236 4770 25248
rect 2406 25168 2412 25220
rect 2464 25208 2470 25220
rect 2501 25211 2559 25217
rect 2501 25208 2513 25211
rect 2464 25180 2513 25208
rect 2464 25168 2470 25180
rect 2501 25177 2513 25180
rect 2547 25208 2559 25211
rect 4890 25208 4896 25220
rect 2547 25180 4896 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 4890 25168 4896 25180
rect 4948 25168 4954 25220
rect 5000 25208 5028 25248
rect 5994 25236 6000 25288
rect 6052 25276 6058 25288
rect 7392 25276 7420 25307
rect 8386 25304 8392 25356
rect 8444 25344 8450 25356
rect 8516 25347 8574 25353
rect 8516 25344 8528 25347
rect 8444 25316 8528 25344
rect 8444 25304 8450 25316
rect 8516 25313 8528 25316
rect 8562 25313 8574 25347
rect 11238 25344 11244 25356
rect 11199 25316 11244 25344
rect 8516 25307 8574 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 9766 25276 9772 25288
rect 6052 25248 7420 25276
rect 9727 25248 9772 25276
rect 6052 25236 6058 25248
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 10134 25276 10140 25288
rect 10095 25248 10140 25276
rect 10134 25236 10140 25248
rect 10192 25236 10198 25288
rect 6730 25208 6736 25220
rect 5000 25180 6736 25208
rect 6730 25168 6736 25180
rect 6788 25208 6794 25220
rect 10502 25208 10508 25220
rect 6788 25180 10508 25208
rect 6788 25168 6794 25180
rect 10502 25168 10508 25180
rect 10560 25168 10566 25220
rect 6822 25140 6828 25152
rect 6783 25112 6828 25140
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 7098 25100 7104 25152
rect 7156 25140 7162 25152
rect 7926 25140 7932 25152
rect 7156 25112 7932 25140
rect 7156 25100 7162 25112
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4212 24908 4257 24936
rect 4212 24896 4218 24908
rect 4522 24896 4528 24948
rect 4580 24936 4586 24948
rect 9766 24945 9772 24948
rect 4893 24939 4951 24945
rect 4893 24936 4905 24939
rect 4580 24908 4905 24936
rect 4580 24896 4586 24908
rect 4893 24905 4905 24908
rect 4939 24905 4951 24939
rect 4893 24899 4951 24905
rect 9493 24939 9551 24945
rect 9493 24905 9505 24939
rect 9539 24936 9551 24939
rect 9723 24939 9772 24945
rect 9723 24936 9735 24939
rect 9539 24908 9735 24936
rect 9539 24905 9551 24908
rect 9493 24899 9551 24905
rect 9723 24905 9735 24908
rect 9769 24905 9772 24939
rect 9723 24899 9772 24905
rect 9766 24896 9772 24899
rect 9824 24896 9830 24948
rect 10410 24936 10416 24948
rect 10371 24908 10416 24936
rect 10410 24896 10416 24908
rect 10468 24896 10474 24948
rect 11238 24936 11244 24948
rect 11199 24908 11244 24936
rect 11238 24896 11244 24908
rect 11296 24896 11302 24948
rect 3145 24871 3203 24877
rect 3145 24837 3157 24871
rect 3191 24868 3203 24871
rect 4062 24868 4068 24880
rect 3191 24840 4068 24868
rect 3191 24837 3203 24840
rect 3145 24831 3203 24837
rect 4062 24828 4068 24840
rect 4120 24868 4126 24880
rect 4430 24868 4436 24880
rect 4120 24840 4436 24868
rect 4120 24828 4126 24840
rect 4430 24828 4436 24840
rect 4488 24828 4494 24880
rect 4617 24871 4675 24877
rect 4617 24837 4629 24871
rect 4663 24868 4675 24871
rect 5810 24868 5816 24880
rect 4663 24840 5816 24868
rect 4663 24837 4675 24840
rect 4617 24831 4675 24837
rect 2961 24735 3019 24741
rect 2961 24701 2973 24735
rect 3007 24732 3019 24735
rect 3878 24732 3884 24744
rect 3007 24704 3884 24732
rect 3007 24701 3019 24704
rect 2961 24695 3019 24701
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 4062 24732 4068 24744
rect 4019 24704 4068 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 4062 24692 4068 24704
rect 4120 24732 4126 24744
rect 4632 24732 4660 24831
rect 5810 24828 5816 24840
rect 5868 24828 5874 24880
rect 5994 24828 6000 24880
rect 6052 24868 6058 24880
rect 6181 24871 6239 24877
rect 6181 24868 6193 24871
rect 6052 24840 6193 24868
rect 6052 24828 6058 24840
rect 6181 24837 6193 24840
rect 6227 24837 6239 24871
rect 6181 24831 6239 24837
rect 9125 24871 9183 24877
rect 9125 24837 9137 24871
rect 9171 24868 9183 24871
rect 11256 24868 11284 24896
rect 9171 24840 11284 24868
rect 9171 24837 9183 24840
rect 9125 24831 9183 24837
rect 5626 24800 5632 24812
rect 5587 24772 5632 24800
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 6880 24772 7113 24800
rect 6880 24760 6886 24772
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 4120 24704 4660 24732
rect 4120 24692 4126 24704
rect 8478 24692 8484 24744
rect 8536 24732 8542 24744
rect 8624 24735 8682 24741
rect 8624 24732 8636 24735
rect 8536 24704 8636 24732
rect 8536 24692 8542 24704
rect 8624 24701 8636 24704
rect 8670 24732 8682 24735
rect 9140 24732 9168 24831
rect 8670 24704 9168 24732
rect 9652 24735 9710 24741
rect 8670 24701 8682 24704
rect 8624 24695 8682 24701
rect 9652 24701 9664 24735
rect 9698 24732 9710 24735
rect 10042 24732 10048 24744
rect 9698 24704 10048 24732
rect 9698 24701 9710 24704
rect 9652 24695 9710 24701
rect 10042 24692 10048 24704
rect 10100 24692 10106 24744
rect 2222 24624 2228 24676
rect 2280 24664 2286 24676
rect 5166 24664 5172 24676
rect 2280 24636 5172 24664
rect 2280 24624 2286 24636
rect 5166 24624 5172 24636
rect 5224 24624 5230 24676
rect 5258 24624 5264 24676
rect 5316 24664 5322 24676
rect 5316 24636 5361 24664
rect 5316 24624 5322 24636
rect 5534 24624 5540 24676
rect 5592 24664 5598 24676
rect 5994 24664 6000 24676
rect 5592 24636 6000 24664
rect 5592 24624 5598 24636
rect 5994 24624 6000 24636
rect 6052 24624 6058 24676
rect 7193 24667 7251 24673
rect 7193 24633 7205 24667
rect 7239 24633 7251 24667
rect 7742 24664 7748 24676
rect 7703 24636 7748 24664
rect 7193 24627 7251 24633
rect 3234 24556 3240 24608
rect 3292 24596 3298 24608
rect 3421 24599 3479 24605
rect 3421 24596 3433 24599
rect 3292 24568 3433 24596
rect 3292 24556 3298 24568
rect 3421 24565 3433 24568
rect 3467 24565 3479 24599
rect 3878 24596 3884 24608
rect 3839 24568 3884 24596
rect 3421 24559 3479 24565
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 4982 24556 4988 24608
rect 5040 24596 5046 24608
rect 5350 24596 5356 24608
rect 5040 24568 5356 24596
rect 5040 24556 5046 24568
rect 5350 24556 5356 24568
rect 5408 24596 5414 24608
rect 6549 24599 6607 24605
rect 6549 24596 6561 24599
rect 5408 24568 6561 24596
rect 5408 24556 5414 24568
rect 6549 24565 6561 24568
rect 6595 24596 6607 24599
rect 6914 24596 6920 24608
rect 6595 24568 6920 24596
rect 6595 24565 6607 24568
rect 6549 24559 6607 24565
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 7208 24596 7236 24627
rect 7742 24624 7748 24636
rect 7800 24624 7806 24676
rect 7926 24624 7932 24676
rect 7984 24664 7990 24676
rect 8386 24664 8392 24676
rect 7984 24636 8392 24664
rect 7984 24624 7990 24636
rect 8386 24624 8392 24636
rect 8444 24624 8450 24676
rect 8711 24667 8769 24673
rect 8711 24633 8723 24667
rect 8757 24664 8769 24667
rect 9306 24664 9312 24676
rect 8757 24636 9312 24664
rect 8757 24633 8769 24636
rect 8711 24627 8769 24633
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 8018 24596 8024 24608
rect 7208 24568 8024 24596
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 2498 24352 2504 24404
rect 2556 24392 2562 24404
rect 3099 24395 3157 24401
rect 3099 24392 3111 24395
rect 2556 24364 3111 24392
rect 2556 24352 2562 24364
rect 3099 24361 3111 24364
rect 3145 24361 3157 24395
rect 3099 24355 3157 24361
rect 3881 24395 3939 24401
rect 3881 24361 3893 24395
rect 3927 24392 3939 24395
rect 4433 24395 4491 24401
rect 4433 24392 4445 24395
rect 3927 24364 4445 24392
rect 3927 24361 3939 24364
rect 3881 24355 3939 24361
rect 4433 24361 4445 24364
rect 4479 24392 4491 24395
rect 4614 24392 4620 24404
rect 4479 24364 4620 24392
rect 4479 24361 4491 24364
rect 4433 24355 4491 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 5258 24352 5264 24404
rect 5316 24392 5322 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 5316 24364 5733 24392
rect 5316 24352 5322 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 6411 24395 6469 24401
rect 6411 24361 6423 24395
rect 6457 24392 6469 24395
rect 6822 24392 6828 24404
rect 6457 24364 6828 24392
rect 6457 24361 6469 24364
rect 6411 24355 6469 24361
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 2087 24327 2145 24333
rect 2087 24293 2099 24327
rect 2133 24293 2145 24327
rect 2087 24287 2145 24293
rect 2102 24256 2130 24287
rect 5166 24284 5172 24336
rect 5224 24324 5230 24336
rect 6089 24327 6147 24333
rect 6089 24324 6101 24327
rect 5224 24296 6101 24324
rect 5224 24284 5230 24296
rect 6089 24293 6101 24296
rect 6135 24293 6147 24327
rect 6089 24287 6147 24293
rect 7469 24327 7527 24333
rect 7469 24293 7481 24327
rect 7515 24324 7527 24327
rect 8018 24324 8024 24336
rect 7515 24296 8024 24324
rect 7515 24293 7527 24296
rect 7469 24287 7527 24293
rect 8018 24284 8024 24296
rect 8076 24284 8082 24336
rect 2222 24256 2228 24268
rect 2102 24228 2228 24256
rect 2222 24216 2228 24228
rect 2280 24216 2286 24268
rect 2866 24216 2872 24268
rect 2924 24256 2930 24268
rect 2996 24259 3054 24265
rect 2996 24256 3008 24259
rect 2924 24228 3008 24256
rect 2924 24216 2930 24228
rect 2996 24225 3008 24228
rect 3042 24225 3054 24259
rect 2996 24219 3054 24225
rect 3970 24216 3976 24268
rect 4028 24256 4034 24268
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 4028 24228 4629 24256
rect 4028 24216 4034 24228
rect 4617 24225 4629 24228
rect 4663 24256 4675 24259
rect 4706 24256 4712 24268
rect 4663 24228 4712 24256
rect 4663 24225 4675 24228
rect 4617 24219 4675 24225
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 4801 24259 4859 24265
rect 4801 24225 4813 24259
rect 4847 24225 4859 24259
rect 4801 24219 4859 24225
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 2038 24188 2044 24200
rect 1903 24160 2044 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 4430 24148 4436 24200
rect 4488 24188 4494 24200
rect 4816 24188 4844 24219
rect 5902 24216 5908 24268
rect 5960 24256 5966 24268
rect 6270 24256 6276 24268
rect 6328 24265 6334 24268
rect 6328 24259 6366 24265
rect 5960 24228 6276 24256
rect 5960 24216 5966 24228
rect 6270 24216 6276 24228
rect 6354 24225 6366 24259
rect 6328 24219 6366 24225
rect 6328 24216 6334 24219
rect 4488 24160 4844 24188
rect 7377 24191 7435 24197
rect 4488 24148 4494 24160
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 7834 24188 7840 24200
rect 7423 24160 7840 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 7834 24148 7840 24160
rect 7892 24148 7898 24200
rect 8021 24191 8079 24197
rect 8021 24157 8033 24191
rect 8067 24188 8079 24191
rect 8846 24188 8852 24200
rect 8067 24160 8852 24188
rect 8067 24157 8079 24160
rect 8021 24151 8079 24157
rect 8846 24148 8852 24160
rect 8904 24148 8910 24200
rect 4522 24080 4528 24132
rect 4580 24120 4586 24132
rect 6825 24123 6883 24129
rect 6825 24120 6837 24123
rect 4580 24092 6837 24120
rect 4580 24080 4586 24092
rect 6825 24089 6837 24092
rect 6871 24120 6883 24123
rect 7098 24120 7104 24132
rect 6871 24092 7104 24120
rect 6871 24089 6883 24092
rect 6825 24083 6883 24089
rect 7098 24080 7104 24092
rect 7156 24080 7162 24132
rect 1673 24055 1731 24061
rect 1673 24021 1685 24055
rect 1719 24052 1731 24055
rect 1762 24052 1768 24064
rect 1719 24024 1768 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 3418 24052 3424 24064
rect 3379 24024 3424 24052
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 5445 24055 5503 24061
rect 5445 24021 5457 24055
rect 5491 24052 5503 24055
rect 5626 24052 5632 24064
rect 5491 24024 5632 24052
rect 5491 24021 5503 24024
rect 5445 24015 5503 24021
rect 5626 24012 5632 24024
rect 5684 24012 5690 24064
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1535 23851 1593 23857
rect 1535 23817 1547 23851
rect 1581 23848 1593 23851
rect 1670 23848 1676 23860
rect 1581 23820 1676 23848
rect 1581 23817 1593 23820
rect 1535 23811 1593 23817
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 4985 23851 5043 23857
rect 4985 23848 4997 23851
rect 4856 23820 4997 23848
rect 4856 23808 4862 23820
rect 4985 23817 4997 23820
rect 5031 23817 5043 23851
rect 4985 23811 5043 23817
rect 3510 23780 3516 23792
rect 3471 23752 3516 23780
rect 3510 23740 3516 23752
rect 3568 23740 3574 23792
rect 3252 23684 3740 23712
rect 1464 23647 1522 23653
rect 1464 23613 1476 23647
rect 1510 23644 1522 23647
rect 1762 23644 1768 23656
rect 1510 23616 1768 23644
rect 1510 23613 1522 23616
rect 1464 23607 1522 23613
rect 1762 23604 1768 23616
rect 1820 23644 1826 23656
rect 2498 23644 2504 23656
rect 1820 23616 2504 23644
rect 1820 23604 1826 23616
rect 2498 23604 2504 23616
rect 2556 23604 2562 23656
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 3050 23468 3056 23520
rect 3108 23508 3114 23520
rect 3252 23517 3280 23684
rect 3418 23644 3424 23656
rect 3379 23616 3424 23644
rect 3418 23604 3424 23616
rect 3476 23604 3482 23656
rect 3712 23653 3740 23684
rect 4522 23672 4528 23724
rect 4580 23712 4586 23724
rect 4798 23712 4804 23724
rect 4580 23684 4804 23712
rect 4580 23672 4586 23684
rect 4798 23672 4804 23684
rect 4856 23672 4862 23724
rect 3697 23647 3755 23653
rect 3697 23613 3709 23647
rect 3743 23613 3755 23647
rect 5000 23644 5028 23811
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 6270 23848 6276 23860
rect 5592 23820 6276 23848
rect 5592 23808 5598 23820
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 13633 23851 13691 23857
rect 13633 23817 13645 23851
rect 13679 23848 13691 23851
rect 15470 23848 15476 23860
rect 13679 23820 15476 23848
rect 13679 23817 13691 23820
rect 13633 23811 13691 23817
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 7834 23740 7840 23792
rect 7892 23780 7898 23792
rect 10275 23783 10333 23789
rect 10275 23780 10287 23783
rect 7892 23752 10287 23780
rect 7892 23740 7898 23752
rect 10275 23749 10287 23752
rect 10321 23749 10333 23783
rect 10275 23743 10333 23749
rect 8662 23712 8668 23724
rect 8623 23684 8668 23712
rect 8662 23672 8668 23684
rect 8720 23672 8726 23724
rect 8846 23672 8852 23724
rect 8904 23712 8910 23724
rect 8941 23715 8999 23721
rect 8941 23712 8953 23715
rect 8904 23684 8953 23712
rect 8904 23672 8910 23684
rect 8941 23681 8953 23684
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 5074 23644 5080 23656
rect 4987 23616 5080 23644
rect 3697 23607 3755 23613
rect 5074 23604 5080 23616
rect 5132 23644 5138 23656
rect 5169 23647 5227 23653
rect 5169 23644 5181 23647
rect 5132 23616 5181 23644
rect 5132 23604 5138 23616
rect 5169 23613 5181 23616
rect 5215 23613 5227 23647
rect 5626 23644 5632 23656
rect 5587 23616 5632 23644
rect 5169 23607 5227 23613
rect 5626 23604 5632 23616
rect 5684 23604 5690 23656
rect 6822 23644 6828 23656
rect 6783 23616 6828 23644
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23644 7803 23647
rect 8202 23644 8208 23656
rect 7791 23616 8208 23644
rect 7791 23613 7803 23616
rect 7745 23607 7803 23613
rect 8202 23604 8208 23616
rect 8260 23604 8266 23656
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10172 23647 10230 23653
rect 10172 23644 10184 23647
rect 10100 23616 10184 23644
rect 10100 23604 10106 23616
rect 10172 23613 10184 23616
rect 10218 23644 10230 23647
rect 10594 23644 10600 23656
rect 10218 23616 10600 23644
rect 10218 23613 10230 23616
rect 10172 23607 10230 23613
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 13078 23604 13084 23656
rect 13136 23644 13142 23656
rect 13449 23647 13507 23653
rect 13449 23644 13461 23647
rect 13136 23616 13461 23644
rect 13136 23604 13142 23616
rect 13449 23613 13461 23616
rect 13495 23644 13507 23647
rect 14001 23647 14059 23653
rect 14001 23644 14013 23647
rect 13495 23616 14013 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 14001 23613 14013 23616
rect 14047 23613 14059 23647
rect 14001 23607 14059 23613
rect 3436 23576 3464 23604
rect 4246 23576 4252 23588
rect 3436 23548 4252 23576
rect 4246 23536 4252 23548
rect 4304 23536 4310 23588
rect 5905 23579 5963 23585
rect 5905 23545 5917 23579
rect 5951 23576 5963 23579
rect 6178 23576 6184 23588
rect 5951 23548 6184 23576
rect 5951 23545 5963 23548
rect 5905 23539 5963 23545
rect 6178 23536 6184 23548
rect 6236 23536 6242 23588
rect 8386 23536 8392 23588
rect 8444 23576 8450 23588
rect 8481 23579 8539 23585
rect 8481 23576 8493 23579
rect 8444 23548 8493 23576
rect 8444 23536 8450 23548
rect 8481 23545 8493 23548
rect 8527 23576 8539 23579
rect 8757 23579 8815 23585
rect 8757 23576 8769 23579
rect 8527 23548 8769 23576
rect 8527 23545 8539 23548
rect 8481 23539 8539 23545
rect 8757 23545 8769 23548
rect 8803 23545 8815 23579
rect 8757 23539 8815 23545
rect 3237 23511 3295 23517
rect 3237 23508 3249 23511
rect 3108 23480 3249 23508
rect 3108 23468 3114 23480
rect 3237 23477 3249 23480
rect 3283 23477 3295 23511
rect 3237 23471 3295 23477
rect 3418 23468 3424 23520
rect 3476 23508 3482 23520
rect 3881 23511 3939 23517
rect 3881 23508 3893 23511
rect 3476 23480 3893 23508
rect 3476 23468 3482 23480
rect 3881 23477 3893 23480
rect 3927 23477 3939 23511
rect 3881 23471 3939 23477
rect 4525 23511 4583 23517
rect 4525 23477 4537 23511
rect 4571 23508 4583 23511
rect 4706 23508 4712 23520
rect 4571 23480 4712 23508
rect 4571 23477 4583 23480
rect 4525 23471 4583 23477
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 7193 23511 7251 23517
rect 7193 23508 7205 23511
rect 7156 23480 7205 23508
rect 7156 23468 7162 23480
rect 7193 23477 7205 23480
rect 7239 23477 7251 23511
rect 8018 23508 8024 23520
rect 7979 23480 8024 23508
rect 7193 23471 7251 23477
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 4430 23304 4436 23316
rect 4391 23276 4436 23304
rect 4430 23264 4436 23276
rect 4488 23264 4494 23316
rect 7834 23304 7840 23316
rect 7795 23276 7840 23304
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 1670 23236 1676 23248
rect 1412 23208 1676 23236
rect 1412 23177 1440 23208
rect 1670 23196 1676 23208
rect 1728 23236 1734 23248
rect 4982 23236 4988 23248
rect 1728 23208 4988 23236
rect 1728 23196 1734 23208
rect 4982 23196 4988 23208
rect 5040 23236 5046 23248
rect 5534 23236 5540 23248
rect 5040 23208 5540 23236
rect 5040 23196 5046 23208
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 6638 23245 6644 23248
rect 6635 23236 6644 23245
rect 6551 23208 6644 23236
rect 6635 23199 6644 23208
rect 6696 23236 6702 23248
rect 7098 23236 7104 23248
rect 6696 23208 7104 23236
rect 6638 23196 6644 23199
rect 6696 23196 6702 23208
rect 7098 23196 7104 23208
rect 7156 23196 7162 23248
rect 8202 23236 8208 23248
rect 8163 23208 8208 23236
rect 8202 23196 8208 23208
rect 8260 23196 8266 23248
rect 8757 23239 8815 23245
rect 8757 23205 8769 23239
rect 8803 23236 8815 23239
rect 8846 23236 8852 23248
rect 8803 23208 8852 23236
rect 8803 23205 8815 23208
rect 8757 23199 8815 23205
rect 8846 23196 8852 23208
rect 8904 23196 8910 23248
rect 9306 23196 9312 23248
rect 9364 23236 9370 23248
rect 9766 23236 9772 23248
rect 9364 23208 9772 23236
rect 9364 23196 9370 23208
rect 9766 23196 9772 23208
rect 9824 23196 9830 23248
rect 9858 23196 9864 23248
rect 9916 23236 9922 23248
rect 9916 23208 9961 23236
rect 9916 23196 9922 23208
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23137 1455 23171
rect 1397 23131 1455 23137
rect 3028 23171 3086 23177
rect 3028 23137 3040 23171
rect 3074 23168 3086 23171
rect 3142 23168 3148 23180
rect 3074 23140 3148 23168
rect 3074 23137 3086 23140
rect 3028 23131 3086 23137
rect 3142 23128 3148 23140
rect 3200 23128 3206 23180
rect 4706 23168 4712 23180
rect 4667 23140 4712 23168
rect 4706 23128 4712 23140
rect 4764 23128 4770 23180
rect 5261 23171 5319 23177
rect 5261 23137 5273 23171
rect 5307 23168 5319 23171
rect 5626 23168 5632 23180
rect 5307 23140 5632 23168
rect 5307 23137 5319 23140
rect 5261 23131 5319 23137
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 7190 23128 7196 23180
rect 7248 23128 7254 23180
rect 7282 23128 7288 23180
rect 7340 23168 7346 23180
rect 7926 23168 7932 23180
rect 7340 23140 7932 23168
rect 7340 23128 7346 23140
rect 7926 23128 7932 23140
rect 7984 23128 7990 23180
rect 5442 23100 5448 23112
rect 5403 23072 5448 23100
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6273 23103 6331 23109
rect 6273 23100 6285 23103
rect 6236 23072 6285 23100
rect 6236 23060 6242 23072
rect 6273 23069 6285 23072
rect 6319 23069 6331 23103
rect 7208 23100 7236 23128
rect 8110 23100 8116 23112
rect 7208 23072 8116 23100
rect 6273 23063 6331 23069
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 10045 23103 10103 23109
rect 10045 23100 10057 23103
rect 9048 23072 10057 23100
rect 3099 23035 3157 23041
rect 3099 23001 3111 23035
rect 3145 23032 3157 23035
rect 6730 23032 6736 23044
rect 3145 23004 6736 23032
rect 3145 23001 3157 23004
rect 3099 22995 3157 23001
rect 6730 22992 6736 23004
rect 6788 22992 6794 23044
rect 7193 23035 7251 23041
rect 7193 23001 7205 23035
rect 7239 23032 7251 23035
rect 8018 23032 8024 23044
rect 7239 23004 8024 23032
rect 7239 23001 7251 23004
rect 7193 22995 7251 23001
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 2958 22924 2964 22976
rect 3016 22964 3022 22976
rect 3421 22967 3479 22973
rect 3421 22964 3433 22967
rect 3016 22936 3433 22964
rect 3016 22924 3022 22936
rect 3421 22933 3433 22936
rect 3467 22964 3479 22967
rect 3510 22964 3516 22976
rect 3467 22936 3516 22964
rect 3467 22933 3479 22936
rect 3421 22927 3479 22933
rect 3510 22924 3516 22936
rect 3568 22924 3574 22976
rect 3881 22967 3939 22973
rect 3881 22933 3893 22967
rect 3927 22964 3939 22967
rect 4338 22964 4344 22976
rect 3927 22936 4344 22964
rect 3927 22933 3939 22936
rect 3881 22927 3939 22933
rect 4338 22924 4344 22936
rect 4396 22924 4402 22976
rect 5902 22924 5908 22976
rect 5960 22964 5966 22976
rect 6822 22964 6828 22976
rect 5960 22936 6828 22964
rect 5960 22924 5966 22936
rect 6822 22924 6828 22936
rect 6880 22964 6886 22976
rect 7469 22967 7527 22973
rect 7469 22964 7481 22967
rect 6880 22936 7481 22964
rect 6880 22924 6886 22936
rect 7469 22933 7481 22936
rect 7515 22933 7527 22967
rect 7469 22927 7527 22933
rect 8570 22924 8576 22976
rect 8628 22964 8634 22976
rect 9048 22973 9076 23072
rect 10045 23069 10057 23072
rect 10091 23069 10103 23103
rect 10045 23063 10103 23069
rect 9033 22967 9091 22973
rect 9033 22964 9045 22967
rect 8628 22936 9045 22964
rect 8628 22924 8634 22936
rect 9033 22933 9045 22936
rect 9079 22933 9091 22967
rect 9033 22927 9091 22933
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 1670 22760 1676 22772
rect 1631 22732 1676 22760
rect 1670 22720 1676 22732
rect 1728 22720 1734 22772
rect 2685 22763 2743 22769
rect 2685 22729 2697 22763
rect 2731 22760 2743 22763
rect 4062 22760 4068 22772
rect 2731 22732 4068 22760
rect 2731 22729 2743 22732
rect 2685 22723 2743 22729
rect 2200 22559 2258 22565
rect 2200 22525 2212 22559
rect 2246 22556 2258 22559
rect 2700 22556 2728 22723
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 4706 22760 4712 22772
rect 4667 22732 4712 22760
rect 4706 22720 4712 22732
rect 4764 22720 4770 22772
rect 6273 22763 6331 22769
rect 6273 22729 6285 22763
rect 6319 22760 6331 22763
rect 6638 22760 6644 22772
rect 6319 22732 6644 22760
rect 6319 22729 6331 22732
rect 6273 22723 6331 22729
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8386 22760 8392 22772
rect 7975 22732 8392 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 9824 22732 10149 22760
rect 9824 22720 9830 22732
rect 10137 22729 10149 22732
rect 10183 22729 10195 22763
rect 10137 22723 10195 22729
rect 2958 22584 2964 22636
rect 3016 22624 3022 22636
rect 3237 22627 3295 22633
rect 3237 22624 3249 22627
rect 3016 22596 3249 22624
rect 3016 22584 3022 22596
rect 3237 22593 3249 22596
rect 3283 22593 3295 22627
rect 3237 22587 3295 22593
rect 3881 22627 3939 22633
rect 3881 22593 3893 22627
rect 3927 22624 3939 22627
rect 3970 22624 3976 22636
rect 3927 22596 3976 22624
rect 3927 22593 3939 22596
rect 3881 22587 3939 22593
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 5442 22584 5448 22636
rect 5500 22624 5506 22636
rect 7009 22627 7067 22633
rect 7009 22624 7021 22627
rect 5500 22596 7021 22624
rect 5500 22584 5506 22596
rect 7009 22593 7021 22596
rect 7055 22624 7067 22627
rect 7466 22624 7472 22636
rect 7055 22596 7472 22624
rect 7055 22593 7067 22596
rect 7009 22587 7067 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 8404 22624 8432 22720
rect 8662 22652 8668 22704
rect 8720 22692 8726 22704
rect 10459 22695 10517 22701
rect 10459 22692 10471 22695
rect 8720 22664 10471 22692
rect 8720 22652 8726 22664
rect 10459 22661 10471 22664
rect 10505 22661 10517 22695
rect 10459 22655 10517 22661
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 8404 22596 9781 22624
rect 9769 22593 9781 22596
rect 9815 22624 9827 22627
rect 9858 22624 9864 22636
rect 9815 22596 9864 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 9858 22584 9864 22596
rect 9916 22584 9922 22636
rect 2246 22528 2728 22556
rect 3145 22559 3203 22565
rect 2246 22525 2258 22528
rect 2200 22519 2258 22525
rect 3145 22525 3157 22559
rect 3191 22525 3203 22559
rect 3145 22519 3203 22525
rect 3160 22488 3188 22519
rect 3326 22516 3332 22568
rect 3384 22556 3390 22568
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 3384 22528 3433 22556
rect 3384 22516 3390 22528
rect 3421 22525 3433 22528
rect 3467 22556 3479 22559
rect 4157 22559 4215 22565
rect 4157 22556 4169 22559
rect 3467 22528 4169 22556
rect 3467 22525 3479 22528
rect 3421 22519 3479 22525
rect 4157 22525 4169 22528
rect 4203 22525 4215 22559
rect 5166 22556 5172 22568
rect 5127 22528 5172 22556
rect 4157 22519 4215 22525
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 5626 22556 5632 22568
rect 5587 22528 5632 22556
rect 5626 22516 5632 22528
rect 5684 22516 5690 22568
rect 5902 22556 5908 22568
rect 5863 22528 5908 22556
rect 5902 22516 5908 22528
rect 5960 22516 5966 22568
rect 9582 22516 9588 22568
rect 9640 22556 9646 22568
rect 10388 22559 10446 22565
rect 10388 22556 10400 22559
rect 9640 22528 10400 22556
rect 9640 22516 9646 22528
rect 10388 22525 10400 22528
rect 10434 22556 10446 22559
rect 10778 22556 10784 22568
rect 10434 22528 10784 22556
rect 10434 22525 10446 22528
rect 10388 22519 10446 22525
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 4338 22488 4344 22500
rect 3160 22460 4344 22488
rect 4338 22448 4344 22460
rect 4396 22448 4402 22500
rect 7098 22448 7104 22500
rect 7156 22488 7162 22500
rect 7330 22491 7388 22497
rect 7330 22488 7342 22491
rect 7156 22460 7342 22488
rect 7156 22448 7162 22460
rect 7330 22457 7342 22460
rect 7376 22457 7388 22491
rect 7330 22451 7388 22457
rect 7926 22448 7932 22500
rect 7984 22488 7990 22500
rect 8570 22488 8576 22500
rect 7984 22460 8576 22488
rect 7984 22448 7990 22460
rect 8570 22448 8576 22460
rect 8628 22488 8634 22500
rect 8849 22491 8907 22497
rect 8849 22488 8861 22491
rect 8628 22460 8861 22488
rect 8628 22448 8634 22460
rect 8849 22457 8861 22460
rect 8895 22457 8907 22491
rect 8849 22451 8907 22457
rect 8941 22491 8999 22497
rect 8941 22457 8953 22491
rect 8987 22457 8999 22491
rect 9490 22488 9496 22500
rect 9451 22460 9496 22488
rect 8941 22451 8999 22457
rect 2271 22423 2329 22429
rect 2271 22389 2283 22423
rect 2317 22420 2329 22423
rect 2774 22420 2780 22432
rect 2317 22392 2780 22420
rect 2317 22389 2329 22392
rect 2271 22383 2329 22389
rect 2774 22380 2780 22392
rect 2832 22380 2838 22432
rect 2958 22420 2964 22432
rect 2919 22392 2964 22420
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 3970 22380 3976 22432
rect 4028 22420 4034 22432
rect 4706 22420 4712 22432
rect 4028 22392 4712 22420
rect 4028 22380 4034 22392
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 6638 22380 6644 22432
rect 6696 22420 6702 22432
rect 8202 22420 8208 22432
rect 6696 22392 8208 22420
rect 6696 22380 6702 22392
rect 8202 22380 8208 22392
rect 8260 22380 8266 22432
rect 8662 22420 8668 22432
rect 8623 22392 8668 22420
rect 8662 22380 8668 22392
rect 8720 22420 8726 22432
rect 8956 22420 8984 22451
rect 9490 22448 9496 22460
rect 9548 22448 9554 22500
rect 8720 22392 8984 22420
rect 8720 22380 8726 22392
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6273 22219 6331 22225
rect 6273 22216 6285 22219
rect 6236 22188 6285 22216
rect 6236 22176 6242 22188
rect 6273 22185 6285 22188
rect 6319 22185 6331 22219
rect 7466 22216 7472 22228
rect 7427 22188 7472 22216
rect 6273 22179 6331 22185
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 8110 22176 8116 22228
rect 8168 22216 8174 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 8168 22188 9045 22216
rect 8168 22176 8174 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 11379 22219 11437 22225
rect 11379 22185 11391 22219
rect 11425 22216 11437 22219
rect 13814 22216 13820 22228
rect 11425 22188 13820 22216
rect 11425 22185 11437 22188
rect 11379 22179 11437 22185
rect 13814 22176 13820 22188
rect 13872 22176 13878 22228
rect 3145 22151 3203 22157
rect 3145 22117 3157 22151
rect 3191 22148 3203 22151
rect 3326 22148 3332 22160
rect 3191 22120 3332 22148
rect 3191 22117 3203 22120
rect 3145 22111 3203 22117
rect 3326 22108 3332 22120
rect 3384 22108 3390 22160
rect 3881 22151 3939 22157
rect 3881 22117 3893 22151
rect 3927 22148 3939 22151
rect 3927 22120 4746 22148
rect 3927 22117 3939 22120
rect 3881 22111 3939 22117
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 3050 22080 3056 22092
rect 1443 22052 2963 22080
rect 3011 22052 3056 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 2317 22015 2375 22021
rect 2317 21981 2329 22015
rect 2363 22012 2375 22015
rect 2406 22012 2412 22024
rect 2363 21984 2412 22012
rect 2363 21981 2375 21984
rect 2317 21975 2375 21981
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2935 22012 2963 22052
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 4062 22040 4068 22092
rect 4120 22080 4126 22092
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 4120 22052 4169 22080
rect 4120 22040 4126 22052
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 4157 22043 4215 22049
rect 4433 22083 4491 22089
rect 4433 22049 4445 22083
rect 4479 22080 4491 22083
rect 4614 22080 4620 22092
rect 4479 22052 4620 22080
rect 4479 22049 4491 22052
rect 4433 22043 4491 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 4718 22080 4746 22120
rect 6546 22108 6552 22160
rect 6604 22148 6610 22160
rect 6641 22151 6699 22157
rect 6641 22148 6653 22151
rect 6604 22120 6653 22148
rect 6604 22108 6610 22120
rect 6641 22117 6653 22120
rect 6687 22117 6699 22151
rect 6641 22111 6699 22117
rect 7193 22151 7251 22157
rect 7193 22117 7205 22151
rect 7239 22148 7251 22151
rect 7926 22148 7932 22160
rect 7239 22120 7932 22148
rect 7239 22117 7251 22120
rect 7193 22111 7251 22117
rect 7926 22108 7932 22120
rect 7984 22108 7990 22160
rect 8202 22148 8208 22160
rect 8163 22120 8208 22148
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 9858 22148 9864 22160
rect 9819 22120 9864 22148
rect 9858 22108 9864 22120
rect 9916 22108 9922 22160
rect 5626 22080 5632 22092
rect 4718 22052 5632 22080
rect 5626 22040 5632 22052
rect 5684 22040 5690 22092
rect 11238 22080 11244 22092
rect 11199 22052 11244 22080
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 4893 22015 4951 22021
rect 2935 21984 4844 22012
rect 106 21904 112 21956
rect 164 21944 170 21956
rect 3142 21944 3148 21956
rect 164 21916 3148 21944
rect 164 21904 170 21916
rect 3142 21904 3148 21916
rect 3200 21944 3206 21956
rect 3421 21947 3479 21953
rect 3421 21944 3433 21947
rect 3200 21916 3433 21944
rect 3200 21904 3206 21916
rect 3421 21913 3433 21916
rect 3467 21913 3479 21947
rect 3421 21907 3479 21913
rect 4154 21904 4160 21956
rect 4212 21944 4218 21956
rect 4249 21947 4307 21953
rect 4249 21944 4261 21947
rect 4212 21916 4261 21944
rect 4212 21904 4218 21916
rect 4249 21913 4261 21916
rect 4295 21913 4307 21947
rect 4816 21944 4844 21984
rect 4893 21981 4905 22015
rect 4939 22012 4951 22015
rect 6362 22012 6368 22024
rect 4939 21984 6368 22012
rect 4939 21981 4951 21984
rect 4893 21975 4951 21981
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 22012 6607 22015
rect 6730 22012 6736 22024
rect 6595 21984 6736 22012
rect 6595 21981 6607 21984
rect 6549 21975 6607 21981
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 8113 22015 8171 22021
rect 8113 21981 8125 22015
rect 8159 22012 8171 22015
rect 8846 22012 8852 22024
rect 8159 21984 8852 22012
rect 8159 21981 8171 21984
rect 8113 21975 8171 21981
rect 8846 21972 8852 21984
rect 8904 21972 8910 22024
rect 9769 22015 9827 22021
rect 9769 21981 9781 22015
rect 9815 21981 9827 22015
rect 10042 22012 10048 22024
rect 10003 21984 10048 22012
rect 9769 21975 9827 21981
rect 8665 21947 8723 21953
rect 4816 21916 7972 21944
rect 4249 21907 4307 21913
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 1857 21879 1915 21885
rect 1857 21876 1869 21879
rect 1452 21848 1869 21876
rect 1452 21836 1458 21848
rect 1857 21845 1869 21848
rect 1903 21845 1915 21879
rect 1857 21839 1915 21845
rect 2314 21836 2320 21888
rect 2372 21876 2378 21888
rect 5166 21876 5172 21888
rect 2372 21848 5172 21876
rect 2372 21836 2378 21848
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 5626 21876 5632 21888
rect 5587 21848 5632 21876
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 7834 21876 7840 21888
rect 7795 21848 7840 21876
rect 7834 21836 7840 21848
rect 7892 21836 7898 21888
rect 7944 21876 7972 21916
rect 8665 21913 8677 21947
rect 8711 21944 8723 21947
rect 8754 21944 8760 21956
rect 8711 21916 8760 21944
rect 8711 21913 8723 21916
rect 8665 21907 8723 21913
rect 8754 21904 8760 21916
rect 8812 21944 8818 21956
rect 9490 21944 9496 21956
rect 8812 21916 9496 21944
rect 8812 21904 8818 21916
rect 9490 21904 9496 21916
rect 9548 21904 9554 21956
rect 9784 21876 9812 21975
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 9950 21876 9956 21888
rect 7944 21848 9956 21876
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 2593 21675 2651 21681
rect 2593 21641 2605 21675
rect 2639 21672 2651 21675
rect 3050 21672 3056 21684
rect 2639 21644 3056 21672
rect 2639 21641 2651 21644
rect 2593 21635 2651 21641
rect 3050 21632 3056 21644
rect 3108 21632 3114 21684
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 4798 21672 4804 21684
rect 4212 21644 4660 21672
rect 4759 21644 4804 21672
rect 4212 21632 4218 21644
rect 4632 21604 4660 21644
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 7285 21675 7343 21681
rect 7285 21641 7297 21675
rect 7331 21672 7343 21675
rect 8202 21672 8208 21684
rect 7331 21644 8208 21672
rect 7331 21641 7343 21644
rect 7285 21635 7343 21641
rect 8202 21632 8208 21644
rect 8260 21672 8266 21684
rect 8665 21675 8723 21681
rect 8665 21672 8677 21675
rect 8260 21644 8677 21672
rect 8260 21632 8266 21644
rect 8665 21641 8677 21644
rect 8711 21641 8723 21675
rect 8665 21635 8723 21641
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 8941 21675 8999 21681
rect 8941 21672 8953 21675
rect 8904 21644 8953 21672
rect 8904 21632 8910 21644
rect 8941 21641 8953 21644
rect 8987 21641 8999 21675
rect 9950 21672 9956 21684
rect 9911 21644 9956 21672
rect 8941 21635 8999 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 4706 21604 4712 21616
rect 4632 21576 4712 21604
rect 4706 21564 4712 21576
rect 4764 21564 4770 21616
rect 2038 21496 2044 21548
rect 2096 21536 2102 21548
rect 4816 21536 4844 21632
rect 5813 21607 5871 21613
rect 5813 21573 5825 21607
rect 5859 21604 5871 21607
rect 9858 21604 9864 21616
rect 5859 21576 9864 21604
rect 5859 21573 5871 21576
rect 5813 21567 5871 21573
rect 9858 21564 9864 21576
rect 9916 21604 9922 21616
rect 10321 21607 10379 21613
rect 10321 21604 10333 21607
rect 9916 21576 10333 21604
rect 9916 21564 9922 21576
rect 10321 21573 10333 21576
rect 10367 21573 10379 21607
rect 10321 21567 10379 21573
rect 2096 21508 4660 21536
rect 2096 21496 2102 21508
rect 1210 21428 1216 21480
rect 1268 21468 1274 21480
rect 1581 21471 1639 21477
rect 1581 21468 1593 21471
rect 1268 21440 1593 21468
rect 1268 21428 1274 21440
rect 1581 21437 1593 21440
rect 1627 21468 1639 21471
rect 1854 21468 1860 21480
rect 1627 21440 1860 21468
rect 1627 21437 1639 21440
rect 1581 21431 1639 21437
rect 1854 21428 1860 21440
rect 1912 21428 1918 21480
rect 3050 21468 3056 21480
rect 3011 21440 3056 21468
rect 3050 21428 3056 21440
rect 3108 21428 3114 21480
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21437 3203 21471
rect 3326 21468 3332 21480
rect 3287 21440 3332 21468
rect 3145 21431 3203 21437
rect 2222 21400 2228 21412
rect 2183 21372 2228 21400
rect 2222 21360 2228 21372
rect 2280 21360 2286 21412
rect 3160 21400 3188 21431
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 2976 21372 3188 21400
rect 3789 21403 3847 21409
rect 2976 21344 3004 21372
rect 3789 21369 3801 21403
rect 3835 21400 3847 21403
rect 4062 21400 4068 21412
rect 3835 21372 4068 21400
rect 3835 21369 3847 21372
rect 3789 21363 3847 21369
rect 4062 21360 4068 21372
rect 4120 21400 4126 21412
rect 4430 21400 4436 21412
rect 4120 21372 4436 21400
rect 4120 21360 4126 21372
rect 4430 21360 4436 21372
rect 4488 21360 4494 21412
rect 2958 21332 2964 21344
rect 2919 21304 2964 21332
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 4632 21332 4660 21508
rect 4724 21508 4844 21536
rect 4724 21400 4752 21508
rect 6362 21496 6368 21548
rect 6420 21536 6426 21548
rect 10965 21539 11023 21545
rect 10965 21536 10977 21539
rect 6420 21508 10977 21536
rect 6420 21496 6426 21508
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 4856 21440 4905 21468
rect 4856 21428 4862 21440
rect 4893 21437 4905 21440
rect 4939 21468 4951 21471
rect 6089 21471 6147 21477
rect 6089 21468 6101 21471
rect 4939 21440 6101 21468
rect 4939 21437 4951 21440
rect 4893 21431 4951 21437
rect 6089 21437 6101 21440
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 7745 21471 7803 21477
rect 7745 21468 7757 21471
rect 6972 21440 7757 21468
rect 6972 21428 6978 21440
rect 7745 21437 7757 21440
rect 7791 21468 7803 21471
rect 7834 21468 7840 21480
rect 7791 21440 7840 21468
rect 7791 21437 7803 21440
rect 7745 21431 7803 21437
rect 7834 21428 7840 21440
rect 7892 21428 7898 21480
rect 10520 21477 10548 21508
rect 10965 21505 10977 21508
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 10505 21471 10563 21477
rect 10505 21437 10517 21471
rect 10551 21437 10563 21471
rect 10505 21431 10563 21437
rect 5214 21403 5272 21409
rect 5214 21400 5226 21403
rect 4724 21372 5226 21400
rect 5214 21369 5226 21372
rect 5260 21369 5272 21403
rect 5214 21363 5272 21369
rect 7098 21360 7104 21412
rect 7156 21400 7162 21412
rect 8110 21409 8116 21412
rect 7561 21403 7619 21409
rect 7561 21400 7573 21403
rect 7156 21372 7573 21400
rect 7156 21360 7162 21372
rect 7561 21369 7573 21372
rect 7607 21400 7619 21403
rect 8066 21403 8116 21409
rect 8066 21400 8078 21403
rect 7607 21372 8078 21400
rect 7607 21369 7619 21372
rect 7561 21363 7619 21369
rect 8066 21369 8078 21372
rect 8112 21369 8116 21403
rect 8066 21363 8116 21369
rect 8110 21360 8116 21363
rect 8168 21360 8174 21412
rect 10318 21360 10324 21412
rect 10376 21400 10382 21412
rect 11238 21400 11244 21412
rect 10376 21372 11244 21400
rect 10376 21360 10382 21372
rect 11238 21360 11244 21372
rect 11296 21400 11302 21412
rect 11333 21403 11391 21409
rect 11333 21400 11345 21403
rect 11296 21372 11345 21400
rect 11296 21360 11302 21372
rect 11333 21369 11345 21372
rect 11379 21369 11391 21403
rect 11333 21363 11391 21369
rect 5810 21332 5816 21344
rect 4632 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 9490 21332 9496 21344
rect 9451 21304 9496 21332
rect 9490 21292 9496 21304
rect 9548 21292 9554 21344
rect 9582 21292 9588 21344
rect 9640 21332 9646 21344
rect 10689 21335 10747 21341
rect 10689 21332 10701 21335
rect 9640 21304 10701 21332
rect 9640 21292 9646 21304
rect 10689 21301 10701 21304
rect 10735 21301 10747 21335
rect 10689 21295 10747 21301
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 1854 21128 1860 21140
rect 1815 21100 1860 21128
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 2222 21128 2228 21140
rect 2183 21100 2228 21128
rect 2222 21088 2228 21100
rect 2280 21128 2286 21140
rect 2280 21100 2728 21128
rect 2280 21088 2286 21100
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 2406 20992 2412 21004
rect 2367 20964 2412 20992
rect 2406 20952 2412 20964
rect 2464 20952 2470 21004
rect 2700 21001 2728 21100
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 3421 21131 3479 21137
rect 3421 21128 3433 21131
rect 3384 21100 3433 21128
rect 3384 21088 3390 21100
rect 3421 21097 3433 21100
rect 3467 21097 3479 21131
rect 4890 21128 4896 21140
rect 4851 21100 4896 21128
rect 3421 21091 3479 21097
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 7193 21131 7251 21137
rect 7193 21128 7205 21131
rect 6788 21100 7205 21128
rect 6788 21088 6794 21100
rect 7193 21097 7205 21100
rect 7239 21097 7251 21131
rect 8110 21128 8116 21140
rect 8071 21100 8116 21128
rect 7193 21091 7251 21097
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 8662 21128 8668 21140
rect 8623 21100 8668 21128
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 3145 21063 3203 21069
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 3234 21060 3240 21072
rect 3191 21032 3240 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 6914 21060 6920 21072
rect 6875 21032 6920 21060
rect 6914 21020 6920 21032
rect 6972 21020 6978 21072
rect 9490 21020 9496 21072
rect 9548 21060 9554 21072
rect 9769 21063 9827 21069
rect 9769 21060 9781 21063
rect 9548 21032 9781 21060
rect 9548 21020 9554 21032
rect 9769 21029 9781 21032
rect 9815 21029 9827 21063
rect 9769 21023 9827 21029
rect 9858 21020 9864 21072
rect 9916 21060 9922 21072
rect 9916 21032 9961 21060
rect 9916 21020 9922 21032
rect 2685 20995 2743 21001
rect 2685 20961 2697 20995
rect 2731 20961 2743 20995
rect 2685 20955 2743 20961
rect 2424 20924 2452 20952
rect 1596 20896 2452 20924
rect 2700 20924 2728 20955
rect 3050 20952 3056 21004
rect 3108 20992 3114 21004
rect 3789 20995 3847 21001
rect 3789 20992 3801 20995
rect 3108 20964 3801 20992
rect 3108 20952 3114 20964
rect 3789 20961 3801 20964
rect 3835 20961 3847 20995
rect 4430 20992 4436 21004
rect 4391 20964 4436 20992
rect 3789 20955 3847 20961
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20992 4767 20995
rect 6178 20992 6184 21004
rect 4755 20964 5580 20992
rect 6139 20964 6184 20992
rect 4755 20961 4767 20964
rect 4709 20955 4767 20961
rect 4614 20924 4620 20936
rect 2700 20896 4620 20924
rect 1596 20865 1624 20896
rect 4614 20884 4620 20896
rect 4672 20924 4678 20936
rect 4724 20924 4752 20955
rect 4672 20896 4752 20924
rect 4672 20884 4678 20896
rect 1581 20859 1639 20865
rect 1581 20825 1593 20859
rect 1627 20825 1639 20859
rect 1581 20819 1639 20825
rect 2222 20816 2228 20868
rect 2280 20856 2286 20868
rect 2501 20859 2559 20865
rect 2501 20856 2513 20859
rect 2280 20828 2513 20856
rect 2280 20816 2286 20828
rect 2501 20825 2513 20828
rect 2547 20825 2559 20859
rect 4522 20856 4528 20868
rect 4483 20828 4528 20856
rect 2501 20819 2559 20825
rect 4522 20816 4528 20828
rect 4580 20816 4586 20868
rect 4341 20791 4399 20797
rect 4341 20757 4353 20791
rect 4387 20788 4399 20791
rect 4430 20788 4436 20800
rect 4387 20760 4436 20788
rect 4387 20757 4399 20760
rect 4341 20751 4399 20757
rect 4430 20748 4436 20760
rect 4488 20748 4494 20800
rect 5552 20797 5580 20964
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6733 20995 6791 21001
rect 6733 20961 6745 20995
rect 6779 20992 6791 20995
rect 7190 20992 7196 21004
rect 6779 20964 7196 20992
rect 6779 20961 6791 20964
rect 6733 20955 6791 20961
rect 7190 20952 7196 20964
rect 7248 20992 7254 21004
rect 9582 20992 9588 21004
rect 7248 20964 9588 20992
rect 7248 20952 7254 20964
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20893 7803 20927
rect 7745 20887 7803 20893
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 5994 20788 6000 20800
rect 5583 20760 6000 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 5994 20748 6000 20760
rect 6052 20748 6058 20800
rect 7558 20788 7564 20800
rect 7519 20760 7564 20788
rect 7558 20748 7564 20760
rect 7616 20788 7622 20800
rect 7760 20788 7788 20887
rect 10318 20856 10324 20868
rect 10279 20828 10324 20856
rect 10318 20816 10324 20828
rect 10376 20816 10382 20868
rect 7616 20760 7788 20788
rect 7616 20748 7622 20760
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 9033 20791 9091 20797
rect 9033 20788 9045 20791
rect 8260 20760 9045 20788
rect 8260 20748 8266 20760
rect 9033 20757 9045 20760
rect 9079 20788 9091 20791
rect 9766 20788 9772 20800
rect 9079 20760 9772 20788
rect 9079 20757 9091 20760
rect 9033 20751 9091 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 3142 20544 3148 20596
rect 3200 20584 3206 20596
rect 4062 20584 4068 20596
rect 3200 20556 4068 20584
rect 3200 20544 3206 20556
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 4522 20544 4528 20596
rect 4580 20584 4586 20596
rect 5261 20587 5319 20593
rect 5261 20584 5273 20587
rect 4580 20556 5273 20584
rect 4580 20544 4586 20556
rect 5261 20553 5273 20556
rect 5307 20553 5319 20587
rect 5261 20547 5319 20553
rect 5626 20544 5632 20596
rect 5684 20584 5690 20596
rect 5905 20587 5963 20593
rect 5905 20584 5917 20587
rect 5684 20556 5917 20584
rect 5684 20544 5690 20556
rect 5905 20553 5917 20556
rect 5951 20584 5963 20587
rect 7190 20584 7196 20596
rect 5951 20556 7196 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 8110 20584 8116 20596
rect 8071 20556 8116 20584
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 9677 20587 9735 20593
rect 9677 20584 9689 20587
rect 9548 20556 9689 20584
rect 9548 20544 9554 20556
rect 9677 20553 9689 20556
rect 9723 20553 9735 20587
rect 9677 20547 9735 20553
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 15470 20584 15476 20596
rect 10183 20556 15476 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 15470 20544 15476 20556
rect 15528 20544 15534 20596
rect 1857 20519 1915 20525
rect 1857 20485 1869 20519
rect 1903 20516 1915 20519
rect 4246 20516 4252 20528
rect 1903 20488 4252 20516
rect 1903 20485 1915 20488
rect 1857 20479 1915 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 4614 20476 4620 20528
rect 4672 20516 4678 20528
rect 5074 20516 5080 20528
rect 4672 20488 5080 20516
rect 4672 20476 4678 20488
rect 5074 20476 5080 20488
rect 5132 20476 5138 20528
rect 9125 20519 9183 20525
rect 9125 20485 9137 20519
rect 9171 20516 9183 20519
rect 9858 20516 9864 20528
rect 9171 20488 9864 20516
rect 9171 20485 9183 20488
rect 9125 20479 9183 20485
rect 9858 20476 9864 20488
rect 9916 20516 9922 20528
rect 10873 20519 10931 20525
rect 10873 20516 10885 20519
rect 9916 20488 10885 20516
rect 9916 20476 9922 20488
rect 10873 20485 10885 20488
rect 10919 20485 10931 20519
rect 10873 20479 10931 20485
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 4709 20451 4767 20457
rect 4709 20448 4721 20451
rect 1636 20420 4721 20448
rect 1636 20408 1642 20420
rect 4709 20417 4721 20420
rect 4755 20417 4767 20451
rect 8202 20448 8208 20460
rect 8163 20420 8208 20448
rect 4709 20411 4767 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 1670 20380 1676 20392
rect 1631 20352 1676 20380
rect 1670 20340 1676 20352
rect 1728 20340 1734 20392
rect 2593 20383 2651 20389
rect 2593 20349 2605 20383
rect 2639 20380 2651 20383
rect 2958 20380 2964 20392
rect 2639 20352 2964 20380
rect 2639 20349 2651 20352
rect 2593 20343 2651 20349
rect 2958 20340 2964 20352
rect 3016 20380 3022 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 3016 20352 3341 20380
rect 3016 20340 3022 20352
rect 3329 20349 3341 20352
rect 3375 20380 3387 20383
rect 4062 20380 4068 20392
rect 3375 20352 4068 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 4246 20380 4252 20392
rect 4207 20352 4252 20380
rect 4246 20340 4252 20352
rect 4304 20340 4310 20392
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20349 4399 20383
rect 4341 20343 4399 20349
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20349 4583 20383
rect 4525 20343 4583 20349
rect 2130 20272 2136 20324
rect 2188 20312 2194 20324
rect 2682 20312 2688 20324
rect 2188 20284 2688 20312
rect 2188 20272 2194 20284
rect 2682 20272 2688 20284
rect 2740 20272 2746 20324
rect 3418 20312 3424 20324
rect 3331 20284 3424 20312
rect 3418 20272 3424 20284
rect 3476 20312 3482 20324
rect 3697 20315 3755 20321
rect 3697 20312 3709 20315
rect 3476 20284 3709 20312
rect 3476 20272 3482 20284
rect 3697 20281 3709 20284
rect 3743 20312 3755 20315
rect 4356 20312 4384 20343
rect 3743 20284 4384 20312
rect 3743 20281 3755 20284
rect 3697 20275 3755 20281
rect 2222 20244 2228 20256
rect 2183 20216 2228 20244
rect 2222 20204 2228 20216
rect 2280 20204 2286 20256
rect 3142 20204 3148 20256
rect 3200 20244 3206 20256
rect 4154 20244 4160 20256
rect 3200 20216 4160 20244
rect 3200 20204 3206 20216
rect 4154 20204 4160 20216
rect 4212 20244 4218 20256
rect 4540 20244 4568 20343
rect 5166 20340 5172 20392
rect 5224 20380 5230 20392
rect 6178 20380 6184 20392
rect 5224 20352 6184 20380
rect 5224 20340 5230 20352
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 7006 20380 7012 20392
rect 6967 20352 7012 20380
rect 7006 20340 7012 20352
rect 7064 20380 7070 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 7064 20352 7665 20380
rect 7064 20340 7070 20352
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 7653 20343 7711 20349
rect 8110 20340 8116 20392
rect 8168 20380 8174 20392
rect 9953 20383 10011 20389
rect 9953 20380 9965 20383
rect 8168 20352 9965 20380
rect 8168 20340 8174 20352
rect 9953 20349 9965 20352
rect 9999 20380 10011 20383
rect 10505 20383 10563 20389
rect 10505 20380 10517 20383
rect 9999 20352 10517 20380
rect 9999 20349 10011 20352
rect 9953 20343 10011 20349
rect 10505 20349 10517 20352
rect 10551 20380 10563 20383
rect 10778 20380 10784 20392
rect 10551 20352 10784 20380
rect 10551 20349 10563 20352
rect 10505 20343 10563 20349
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 4706 20272 4712 20324
rect 4764 20312 4770 20324
rect 6549 20315 6607 20321
rect 6549 20312 6561 20315
rect 4764 20284 6561 20312
rect 4764 20272 4770 20284
rect 6549 20281 6561 20284
rect 6595 20312 6607 20315
rect 6825 20315 6883 20321
rect 6825 20312 6837 20315
rect 6595 20284 6837 20312
rect 6595 20281 6607 20284
rect 6549 20275 6607 20281
rect 6825 20281 6837 20284
rect 6871 20281 6883 20315
rect 6825 20275 6883 20281
rect 8018 20272 8024 20324
rect 8076 20312 8082 20324
rect 8526 20315 8584 20321
rect 8526 20312 8538 20315
rect 8076 20284 8538 20312
rect 8076 20272 8082 20284
rect 8526 20281 8538 20284
rect 8572 20281 8584 20315
rect 8526 20275 8584 20281
rect 4212 20216 4568 20244
rect 4212 20204 4218 20216
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6696 20216 7113 20244
rect 6696 20204 6702 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 1946 20040 1952 20052
rect 1412 20012 1952 20040
rect 1412 19913 1440 20012
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 3418 20040 3424 20052
rect 3379 20012 3424 20040
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 4798 20040 4804 20052
rect 4759 20012 4804 20040
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 7190 20040 7196 20052
rect 7151 20012 7196 20040
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 9766 20040 9772 20052
rect 9727 20012 9772 20040
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 1670 19932 1676 19984
rect 1728 19972 1734 19984
rect 2317 19975 2375 19981
rect 2317 19972 2329 19975
rect 1728 19944 2329 19972
rect 1728 19932 1734 19944
rect 2317 19941 2329 19944
rect 2363 19972 2375 19975
rect 3326 19972 3332 19984
rect 2363 19944 3332 19972
rect 2363 19941 2375 19944
rect 2317 19935 2375 19941
rect 3326 19932 3332 19944
rect 3384 19932 3390 19984
rect 3510 19932 3516 19984
rect 3568 19972 3574 19984
rect 4614 19972 4620 19984
rect 3568 19944 4620 19972
rect 3568 19932 3574 19944
rect 4614 19932 4620 19944
rect 4672 19932 4678 19984
rect 4890 19932 4896 19984
rect 4948 19972 4954 19984
rect 6411 19975 6469 19981
rect 6411 19972 6423 19975
rect 4948 19944 6423 19972
rect 4948 19932 4954 19944
rect 6411 19941 6423 19944
rect 6457 19941 6469 19975
rect 6411 19935 6469 19941
rect 7831 19975 7889 19981
rect 7831 19941 7843 19975
rect 7877 19972 7889 19975
rect 8018 19972 8024 19984
rect 7877 19944 8024 19972
rect 7877 19941 7889 19944
rect 7831 19935 7889 19941
rect 8018 19932 8024 19944
rect 8076 19972 8082 19984
rect 8665 19975 8723 19981
rect 8665 19972 8677 19975
rect 8076 19944 8677 19972
rect 8076 19932 8082 19944
rect 8665 19941 8677 19944
rect 8711 19941 8723 19975
rect 8665 19935 8723 19941
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19873 1455 19907
rect 1397 19867 1455 19873
rect 2590 19864 2596 19916
rect 2648 19904 2654 19916
rect 3053 19907 3111 19913
rect 3053 19904 3065 19907
rect 2648 19876 3065 19904
rect 2648 19864 2654 19876
rect 3053 19873 3065 19876
rect 3099 19904 3111 19907
rect 4522 19904 4528 19916
rect 3099 19876 4528 19904
rect 3099 19873 3111 19876
rect 3053 19867 3111 19873
rect 4522 19864 4528 19876
rect 4580 19864 4586 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4902 19876 5181 19904
rect 2222 19796 2228 19848
rect 2280 19836 2286 19848
rect 3145 19839 3203 19845
rect 3145 19836 3157 19839
rect 2280 19808 3157 19836
rect 2280 19796 2286 19808
rect 3145 19805 3157 19808
rect 3191 19805 3203 19839
rect 3145 19799 3203 19805
rect 3160 19768 3188 19799
rect 3970 19796 3976 19848
rect 4028 19836 4034 19848
rect 4902 19836 4930 19876
rect 5169 19873 5181 19876
rect 5215 19873 5227 19907
rect 5169 19867 5227 19873
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 6324 19907 6382 19913
rect 6324 19904 6336 19907
rect 5868 19876 6336 19904
rect 5868 19864 5874 19876
rect 6324 19873 6336 19876
rect 6370 19904 6382 19907
rect 6730 19904 6736 19916
rect 6370 19876 6736 19904
rect 6370 19873 6382 19876
rect 6324 19867 6382 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9674 19904 9680 19916
rect 9456 19876 9680 19904
rect 9456 19864 9462 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 7466 19836 7472 19848
rect 4028 19808 4930 19836
rect 7427 19808 7472 19836
rect 4028 19796 4034 19808
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 10152 19836 10180 19867
rect 9548 19808 10180 19836
rect 9548 19796 9554 19808
rect 4706 19768 4712 19780
rect 3160 19740 4712 19768
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 4798 19728 4804 19780
rect 4856 19768 4862 19780
rect 6089 19771 6147 19777
rect 6089 19768 6101 19771
rect 4856 19740 6101 19768
rect 4856 19728 4862 19740
rect 6089 19737 6101 19740
rect 6135 19737 6147 19771
rect 6089 19731 6147 19737
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 1762 19700 1768 19712
rect 1627 19672 1768 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 3234 19660 3240 19712
rect 3292 19700 3298 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3292 19672 3801 19700
rect 3292 19660 3298 19672
rect 3789 19669 3801 19672
rect 3835 19700 3847 19703
rect 4246 19700 4252 19712
rect 3835 19672 4252 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4430 19700 4436 19712
rect 4391 19672 4436 19700
rect 4430 19660 4436 19672
rect 4488 19660 4494 19712
rect 4617 19703 4675 19709
rect 4617 19669 4629 19703
rect 4663 19700 4675 19703
rect 5534 19700 5540 19712
rect 4663 19672 5540 19700
rect 4663 19669 4675 19672
rect 4617 19663 4675 19669
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 5813 19703 5871 19709
rect 5813 19669 5825 19703
rect 5859 19700 5871 19703
rect 5994 19700 6000 19712
rect 5859 19672 6000 19700
rect 5859 19669 5871 19672
rect 5813 19663 5871 19669
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7098 19700 7104 19712
rect 6963 19672 7104 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 4522 19456 4528 19508
rect 4580 19496 4586 19508
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 4580 19468 4629 19496
rect 4580 19456 4586 19468
rect 4617 19465 4629 19468
rect 4663 19496 4675 19499
rect 4663 19468 4936 19496
rect 4663 19465 4675 19468
rect 4617 19459 4675 19465
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2590 19428 2596 19440
rect 2547 19400 2596 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2590 19388 2596 19400
rect 2648 19388 2654 19440
rect 3050 19388 3056 19440
rect 3108 19428 3114 19440
rect 4908 19437 4936 19468
rect 5810 19456 5816 19508
rect 5868 19496 5874 19508
rect 10594 19496 10600 19508
rect 5868 19468 10600 19496
rect 5868 19456 5874 19468
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 3375 19431 3433 19437
rect 3375 19428 3387 19431
rect 3108 19400 3387 19428
rect 3108 19388 3114 19400
rect 3375 19397 3387 19400
rect 3421 19397 3433 19431
rect 3375 19391 3433 19397
rect 3513 19431 3571 19437
rect 3513 19397 3525 19431
rect 3559 19397 3571 19431
rect 3513 19391 3571 19397
rect 4893 19431 4951 19437
rect 4893 19397 4905 19431
rect 4939 19397 4951 19431
rect 4893 19391 4951 19397
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 3068 19360 3096 19388
rect 2179 19332 3096 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 3142 19320 3148 19372
rect 3200 19360 3206 19372
rect 3200 19332 3372 19360
rect 3200 19320 3206 19332
rect 1486 19292 1492 19304
rect 1447 19264 1492 19292
rect 1486 19252 1492 19264
rect 1544 19252 1550 19304
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3344 19292 3372 19332
rect 2924 19264 3372 19292
rect 2924 19252 2930 19264
rect 1762 19184 1768 19236
rect 1820 19224 1826 19236
rect 2314 19224 2320 19236
rect 1820 19196 2320 19224
rect 1820 19184 1826 19196
rect 2314 19184 2320 19196
rect 2372 19224 2378 19236
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 2372 19196 3249 19224
rect 2372 19184 2378 19196
rect 3237 19193 3249 19196
rect 3283 19193 3295 19227
rect 3344 19224 3372 19264
rect 3418 19252 3424 19304
rect 3476 19292 3482 19304
rect 3528 19292 3556 19391
rect 5258 19388 5264 19440
rect 5316 19428 5322 19440
rect 6914 19428 6920 19440
rect 5316 19400 6920 19428
rect 5316 19388 5322 19400
rect 6914 19388 6920 19400
rect 6972 19428 6978 19440
rect 7929 19431 7987 19437
rect 7929 19428 7941 19431
rect 6972 19400 7941 19428
rect 6972 19388 6978 19400
rect 7929 19397 7941 19400
rect 7975 19428 7987 19431
rect 8018 19428 8024 19440
rect 7975 19400 8024 19428
rect 7975 19397 7987 19400
rect 7929 19391 7987 19397
rect 8018 19388 8024 19400
rect 8076 19388 8082 19440
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 9217 19431 9275 19437
rect 9217 19428 9229 19431
rect 8812 19400 9229 19428
rect 8812 19388 8818 19400
rect 9217 19397 9229 19400
rect 9263 19397 9275 19431
rect 9217 19391 9275 19397
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3476 19264 3556 19292
rect 3476 19252 3482 19264
rect 3620 19224 3648 19323
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 4430 19360 4436 19372
rect 3752 19332 4436 19360
rect 3752 19320 3758 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 7558 19360 7564 19372
rect 7519 19332 7564 19360
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19360 8539 19363
rect 8665 19363 8723 19369
rect 8665 19360 8677 19363
rect 8527 19332 8677 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8665 19329 8677 19332
rect 8711 19360 8723 19363
rect 10137 19363 10195 19369
rect 10137 19360 10149 19363
rect 8711 19332 10149 19360
rect 8711 19329 8723 19332
rect 8665 19323 8723 19329
rect 10137 19329 10149 19332
rect 10183 19329 10195 19363
rect 10137 19323 10195 19329
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 4798 19292 4804 19304
rect 3936 19264 4804 19292
rect 3936 19252 3942 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5994 19292 6000 19304
rect 5123 19264 6000 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5994 19252 6000 19264
rect 6052 19252 6058 19304
rect 7098 19292 7104 19304
rect 7059 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7190 19252 7196 19304
rect 7248 19292 7254 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7248 19264 7297 19292
rect 7248 19252 7254 19264
rect 7285 19261 7297 19264
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 3344 19196 3648 19224
rect 3237 19187 3295 19193
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 4982 19224 4988 19236
rect 4212 19196 4988 19224
rect 4212 19184 4218 19196
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 8386 19184 8392 19236
rect 8444 19224 8450 19236
rect 8757 19227 8815 19233
rect 8757 19224 8769 19227
rect 8444 19196 8769 19224
rect 8444 19184 8450 19196
rect 8757 19193 8769 19196
rect 8803 19193 8815 19227
rect 8757 19187 8815 19193
rect 9490 19184 9496 19236
rect 9548 19224 9554 19236
rect 10597 19227 10655 19233
rect 10597 19224 10609 19227
rect 9548 19196 10609 19224
rect 9548 19184 9554 19196
rect 10597 19193 10609 19196
rect 10643 19193 10655 19227
rect 10597 19187 10655 19193
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3881 19159 3939 19165
rect 3881 19156 3893 19159
rect 3384 19128 3893 19156
rect 3384 19116 3390 19128
rect 3881 19125 3893 19128
rect 3927 19125 3939 19159
rect 3881 19119 3939 19125
rect 3970 19116 3976 19168
rect 4028 19156 4034 19168
rect 4246 19156 4252 19168
rect 4028 19128 4252 19156
rect 4028 19116 4034 19128
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 5261 19159 5319 19165
rect 5261 19156 5273 19159
rect 4764 19128 5273 19156
rect 4764 19116 4770 19128
rect 5261 19125 5273 19128
rect 5307 19125 5319 19159
rect 5261 19119 5319 19125
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 5813 19159 5871 19165
rect 5813 19156 5825 19159
rect 5592 19128 5825 19156
rect 5592 19116 5598 19128
rect 5813 19125 5825 19128
rect 5859 19125 5871 19159
rect 5813 19119 5871 19125
rect 6365 19159 6423 19165
rect 6365 19125 6377 19159
rect 6411 19156 6423 19159
rect 6730 19156 6736 19168
rect 6411 19128 6736 19156
rect 6411 19125 6423 19128
rect 6365 19119 6423 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 9674 19156 9680 19168
rect 8260 19128 9680 19156
rect 8260 19116 8266 19128
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 1394 18912 1400 18964
rect 1452 18952 1458 18964
rect 2869 18955 2927 18961
rect 2869 18952 2881 18955
rect 1452 18924 2881 18952
rect 1452 18912 1458 18924
rect 2869 18921 2881 18924
rect 2915 18921 2927 18955
rect 2869 18915 2927 18921
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3108 18924 3801 18952
rect 3108 18912 3114 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 5994 18952 6000 18964
rect 5955 18924 6000 18952
rect 3789 18915 3847 18921
rect 5994 18912 6000 18924
rect 6052 18912 6058 18964
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8444 18924 8585 18952
rect 8444 18912 8450 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 9766 18952 9772 18964
rect 9727 18924 9772 18952
rect 8573 18915 8631 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 2317 18887 2375 18893
rect 2317 18853 2329 18887
rect 2363 18884 2375 18887
rect 3068 18884 3096 18912
rect 2363 18856 3096 18884
rect 5163 18887 5221 18893
rect 2363 18853 2375 18856
rect 2317 18847 2375 18853
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1578 18816 1584 18828
rect 1443 18788 1584 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 2424 18825 2452 18856
rect 5163 18853 5175 18887
rect 5209 18884 5221 18887
rect 5258 18884 5264 18896
rect 5209 18856 5264 18884
rect 5209 18853 5221 18856
rect 5163 18847 5221 18853
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 5534 18844 5540 18896
rect 5592 18884 5598 18896
rect 7285 18887 7343 18893
rect 5592 18856 6592 18884
rect 5592 18844 5598 18856
rect 2409 18819 2467 18825
rect 2409 18816 2421 18819
rect 2387 18788 2421 18816
rect 2409 18785 2421 18788
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 2685 18819 2743 18825
rect 2685 18785 2697 18819
rect 2731 18816 2743 18819
rect 2866 18816 2872 18828
rect 2731 18788 2872 18816
rect 2731 18785 2743 18788
rect 2685 18779 2743 18785
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 2958 18776 2964 18828
rect 3016 18816 3022 18828
rect 6365 18819 6423 18825
rect 6365 18816 6377 18819
rect 3016 18788 6377 18816
rect 3016 18776 3022 18788
rect 6365 18785 6377 18788
rect 6411 18816 6423 18819
rect 6454 18816 6460 18828
rect 6411 18788 6460 18816
rect 6411 18785 6423 18788
rect 6365 18779 6423 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 6564 18825 6592 18856
rect 7285 18853 7297 18887
rect 7331 18884 7343 18887
rect 7466 18884 7472 18896
rect 7331 18856 7472 18884
rect 7331 18853 7343 18856
rect 7285 18847 7343 18853
rect 7466 18844 7472 18856
rect 7524 18884 7530 18896
rect 7561 18887 7619 18893
rect 7561 18884 7573 18887
rect 7524 18856 7573 18884
rect 7524 18844 7530 18856
rect 7561 18853 7573 18856
rect 7607 18853 7619 18887
rect 7561 18847 7619 18853
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7190 18816 7196 18828
rect 7147 18788 7196 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 8110 18816 8116 18828
rect 8071 18788 8116 18816
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9548 18788 9689 18816
rect 9548 18776 9554 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 10134 18816 10140 18828
rect 10095 18788 10140 18816
rect 9677 18779 9735 18785
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 3418 18748 3424 18760
rect 2372 18720 3424 18748
rect 2372 18708 2378 18720
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 4338 18748 4344 18760
rect 3568 18720 4344 18748
rect 3568 18708 3574 18720
rect 4338 18708 4344 18720
rect 4396 18708 4402 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 5258 18748 5264 18760
rect 4847 18720 5264 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 1581 18683 1639 18689
rect 1581 18649 1593 18683
rect 1627 18680 1639 18683
rect 2501 18683 2559 18689
rect 1627 18652 2452 18680
rect 1627 18649 1639 18652
rect 1581 18643 1639 18649
rect 658 18572 664 18624
rect 716 18612 722 18624
rect 1486 18612 1492 18624
rect 716 18584 1492 18612
rect 716 18572 722 18584
rect 1486 18572 1492 18584
rect 1544 18612 1550 18624
rect 1857 18615 1915 18621
rect 1857 18612 1869 18615
rect 1544 18584 1869 18612
rect 1544 18572 1550 18584
rect 1857 18581 1869 18584
rect 1903 18581 1915 18615
rect 2424 18612 2452 18652
rect 2501 18649 2513 18683
rect 2547 18680 2559 18683
rect 4062 18680 4068 18692
rect 2547 18652 4068 18680
rect 2547 18649 2559 18652
rect 2501 18643 2559 18649
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 4706 18680 4712 18692
rect 4663 18652 4712 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 4706 18640 4712 18652
rect 4764 18680 4770 18692
rect 10134 18680 10140 18692
rect 4764 18652 10140 18680
rect 4764 18640 4770 18652
rect 10134 18640 10140 18652
rect 10192 18640 10198 18692
rect 4246 18612 4252 18624
rect 2424 18584 4252 18612
rect 1857 18575 1915 18581
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 5721 18615 5779 18621
rect 5721 18612 5733 18615
rect 5040 18584 5733 18612
rect 5040 18572 5046 18584
rect 5721 18581 5733 18584
rect 5767 18581 5779 18615
rect 5721 18575 5779 18581
rect 8251 18615 8309 18621
rect 8251 18581 8263 18615
rect 8297 18612 8309 18615
rect 10410 18612 10416 18624
rect 8297 18584 10416 18612
rect 8297 18581 8309 18584
rect 8251 18575 8309 18581
rect 10410 18572 10416 18584
rect 10468 18612 10474 18624
rect 10689 18615 10747 18621
rect 10689 18612 10701 18615
rect 10468 18584 10701 18612
rect 10468 18572 10474 18584
rect 10689 18581 10701 18584
rect 10735 18581 10747 18615
rect 10689 18575 10747 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2409 18411 2467 18417
rect 2409 18408 2421 18411
rect 2004 18380 2421 18408
rect 2004 18368 2010 18380
rect 2409 18377 2421 18380
rect 2455 18408 2467 18411
rect 2593 18411 2651 18417
rect 2593 18408 2605 18411
rect 2455 18380 2605 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 2593 18377 2605 18380
rect 2639 18377 2651 18411
rect 2593 18371 2651 18377
rect 2682 18368 2688 18420
rect 2740 18408 2746 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2740 18380 2789 18408
rect 2740 18368 2746 18380
rect 2777 18377 2789 18380
rect 2823 18408 2835 18411
rect 4062 18408 4068 18420
rect 2823 18380 3366 18408
rect 4023 18380 4068 18408
rect 2823 18377 2835 18380
rect 2777 18371 2835 18377
rect 1857 18343 1915 18349
rect 1857 18309 1869 18343
rect 1903 18340 1915 18343
rect 2866 18340 2872 18352
rect 1903 18312 2872 18340
rect 1903 18309 1915 18312
rect 1857 18303 1915 18309
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 3068 18349 3096 18380
rect 3053 18343 3111 18349
rect 3053 18309 3065 18343
rect 3099 18309 3111 18343
rect 3053 18303 3111 18309
rect 3234 18300 3240 18352
rect 3292 18300 3298 18352
rect 3338 18340 3366 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 4341 18411 4399 18417
rect 4341 18408 4353 18411
rect 4304 18380 4353 18408
rect 4304 18368 4310 18380
rect 4341 18377 4353 18380
rect 4387 18408 4399 18411
rect 4387 18380 5028 18408
rect 4387 18377 4399 18380
rect 4341 18371 4399 18377
rect 4798 18340 4804 18352
rect 3338 18312 4804 18340
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3252 18272 3280 18300
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 2639 18244 3188 18272
rect 3252 18244 3433 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 1946 18204 1952 18216
rect 1910 18176 1952 18204
rect 1946 18164 1952 18176
rect 2004 18213 2010 18216
rect 2004 18207 2058 18213
rect 2004 18173 2012 18207
rect 2046 18204 2058 18207
rect 2774 18204 2780 18216
rect 2046 18176 2780 18204
rect 2046 18173 2058 18176
rect 2004 18167 2058 18173
rect 2004 18164 2010 18167
rect 2774 18164 2780 18176
rect 2832 18164 2838 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 3050 18204 3056 18216
rect 3007 18176 3056 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3160 18204 3188 18244
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3237 18207 3295 18213
rect 3237 18204 3249 18207
rect 3160 18176 3249 18204
rect 3237 18173 3249 18176
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4706 18204 4712 18216
rect 4028 18176 4712 18204
rect 4028 18164 4034 18176
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5000 18213 5028 18380
rect 5350 18368 5356 18420
rect 5408 18408 5414 18420
rect 8110 18408 8116 18420
rect 5408 18380 7328 18408
rect 8071 18380 8116 18408
rect 5408 18368 5414 18380
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 5537 18343 5595 18349
rect 5537 18340 5549 18343
rect 5500 18312 5549 18340
rect 5500 18300 5506 18312
rect 5537 18309 5549 18312
rect 5583 18309 5595 18343
rect 5537 18303 5595 18309
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 7300 18340 7328 18380
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 10134 18408 10140 18420
rect 10095 18380 10140 18408
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 6696 18312 7236 18340
rect 7300 18312 10548 18340
rect 6696 18300 6702 18312
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 7208 18281 7236 18312
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6512 18244 6929 18272
rect 6512 18232 6518 18244
rect 6917 18241 6929 18244
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 9490 18232 9496 18284
rect 9548 18272 9554 18284
rect 9769 18275 9827 18281
rect 9769 18272 9781 18275
rect 9548 18244 9781 18272
rect 9548 18232 9554 18244
rect 9769 18241 9781 18244
rect 9815 18241 9827 18275
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 9769 18235 9827 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10520 18272 10548 18312
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10520 18244 10701 18272
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10689 18235 10747 18241
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 6181 18207 6239 18213
rect 6181 18204 6193 18207
rect 5592 18176 6193 18204
rect 5592 18164 5598 18176
rect 6181 18173 6193 18176
rect 6227 18173 6239 18207
rect 6181 18167 6239 18173
rect 2087 18139 2145 18145
rect 2087 18105 2099 18139
rect 2133 18136 2145 18139
rect 5074 18136 5080 18148
rect 2133 18108 5080 18136
rect 2133 18105 2145 18108
rect 2087 18099 2145 18105
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 5258 18136 5264 18148
rect 5219 18108 5264 18136
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 7006 18136 7012 18148
rect 6967 18108 7012 18136
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 8846 18136 8852 18148
rect 8807 18108 8852 18136
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 8941 18139 8999 18145
rect 8941 18105 8953 18139
rect 8987 18105 8999 18139
rect 8941 18099 8999 18105
rect 9493 18139 9551 18145
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 10505 18139 10563 18145
rect 9539 18108 9996 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 6641 18071 6699 18077
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 7190 18068 7196 18080
rect 6687 18040 7196 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8573 18071 8631 18077
rect 8573 18068 8585 18071
rect 8352 18040 8585 18068
rect 8352 18028 8358 18040
rect 8573 18037 8585 18040
rect 8619 18068 8631 18071
rect 8956 18068 8984 18099
rect 8619 18040 8984 18068
rect 9968 18068 9996 18108
rect 10505 18105 10517 18139
rect 10551 18136 10563 18139
rect 10686 18136 10692 18148
rect 10551 18108 10692 18136
rect 10551 18105 10563 18108
rect 10505 18099 10563 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 10594 18068 10600 18080
rect 9968 18040 10600 18068
rect 8619 18037 8631 18040
rect 8573 18031 8631 18037
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3108 17836 3341 17864
rect 3108 17824 3114 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 3329 17827 3387 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 7193 17867 7251 17873
rect 7193 17833 7205 17867
rect 7239 17864 7251 17867
rect 7374 17864 7380 17876
rect 7239 17836 7380 17864
rect 7239 17833 7251 17836
rect 7193 17827 7251 17833
rect 7374 17824 7380 17836
rect 7432 17864 7438 17876
rect 9766 17864 9772 17876
rect 7432 17836 9772 17864
rect 7432 17824 7438 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2222 17796 2228 17808
rect 1820 17768 2228 17796
rect 1820 17756 1826 17768
rect 2222 17756 2228 17768
rect 2280 17756 2286 17808
rect 4341 17799 4399 17805
rect 4341 17765 4353 17799
rect 4387 17796 4399 17799
rect 4982 17796 4988 17808
rect 4387 17768 4988 17796
rect 4387 17765 4399 17768
rect 4341 17759 4399 17765
rect 4982 17756 4988 17768
rect 5040 17756 5046 17808
rect 5074 17756 5080 17808
rect 5132 17796 5138 17808
rect 5537 17799 5595 17805
rect 5537 17796 5549 17799
rect 5132 17768 5549 17796
rect 5132 17756 5138 17768
rect 5537 17765 5549 17768
rect 5583 17796 5595 17799
rect 5813 17799 5871 17805
rect 5813 17796 5825 17799
rect 5583 17768 5825 17796
rect 5583 17765 5595 17768
rect 5537 17759 5595 17765
rect 5813 17765 5825 17768
rect 5859 17765 5871 17799
rect 5813 17759 5871 17765
rect 5905 17799 5963 17805
rect 5905 17765 5917 17799
rect 5951 17796 5963 17799
rect 5994 17796 6000 17808
rect 5951 17768 6000 17796
rect 5951 17765 5963 17768
rect 5905 17759 5963 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 6086 17756 6092 17808
rect 6144 17796 6150 17808
rect 9490 17796 9496 17808
rect 6144 17768 9496 17796
rect 6144 17756 6150 17768
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3142 17728 3148 17740
rect 3007 17700 3148 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 7300 17737 7328 17768
rect 9490 17756 9496 17768
rect 9548 17756 9554 17808
rect 9861 17799 9919 17805
rect 9861 17765 9873 17799
rect 9907 17796 9919 17799
rect 10134 17796 10140 17808
rect 9907 17768 10140 17796
rect 9907 17765 9919 17768
rect 9861 17759 9919 17765
rect 10134 17756 10140 17768
rect 10192 17756 10198 17808
rect 7285 17731 7343 17737
rect 7285 17697 7297 17731
rect 7331 17697 7343 17731
rect 7834 17728 7840 17740
rect 7795 17700 7840 17728
rect 7285 17691 7343 17697
rect 7834 17688 7840 17700
rect 7892 17688 7898 17740
rect 10502 17688 10508 17740
rect 10560 17728 10566 17740
rect 11276 17731 11334 17737
rect 11276 17728 11288 17731
rect 10560 17700 11288 17728
rect 10560 17688 10566 17700
rect 11276 17697 11288 17700
rect 11322 17728 11334 17731
rect 11698 17728 11704 17740
rect 11322 17700 11704 17728
rect 11322 17697 11334 17700
rect 11276 17691 11334 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 2314 17660 2320 17672
rect 2275 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 4120 17632 4261 17660
rect 4120 17620 4126 17632
rect 4249 17629 4261 17632
rect 4295 17660 4307 17663
rect 4890 17660 4896 17672
rect 4295 17632 4896 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4890 17620 4896 17632
rect 4948 17620 4954 17672
rect 4982 17620 4988 17672
rect 5040 17660 5046 17672
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 5040 17632 6745 17660
rect 5040 17620 5046 17632
rect 6733 17629 6745 17632
rect 6779 17660 6791 17663
rect 7006 17660 7012 17672
rect 6779 17632 7012 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 8018 17660 8024 17672
rect 7979 17632 8024 17660
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9539 17632 9781 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 9769 17629 9781 17632
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10410 17660 10416 17672
rect 10371 17632 10416 17660
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 4801 17595 4859 17601
rect 4801 17561 4813 17595
rect 4847 17592 4859 17595
rect 5350 17592 5356 17604
rect 4847 17564 5356 17592
rect 4847 17561 4859 17564
rect 4801 17555 4859 17561
rect 5350 17552 5356 17564
rect 5408 17552 5414 17604
rect 6365 17595 6423 17601
rect 6365 17561 6377 17595
rect 6411 17592 6423 17595
rect 6638 17592 6644 17604
rect 6411 17564 6644 17592
rect 6411 17561 6423 17564
rect 6365 17555 6423 17561
rect 6638 17552 6644 17564
rect 6696 17552 6702 17604
rect 10686 17592 10692 17604
rect 8541 17564 10692 17592
rect 2222 17484 2228 17536
rect 2280 17524 2286 17536
rect 5810 17524 5816 17536
rect 2280 17496 5816 17524
rect 2280 17484 2286 17496
rect 5810 17484 5816 17496
rect 5868 17484 5874 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 8541 17524 8569 17564
rect 10686 17552 10692 17564
rect 10744 17552 10750 17604
rect 8846 17524 8852 17536
rect 6052 17496 8569 17524
rect 8807 17496 8852 17524
rect 6052 17484 6058 17496
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11379 17527 11437 17533
rect 11379 17524 11391 17527
rect 10836 17496 11391 17524
rect 10836 17484 10842 17496
rect 11379 17493 11391 17496
rect 11425 17493 11437 17527
rect 11379 17487 11437 17493
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2314 17320 2320 17332
rect 2271 17292 2320 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4982 17320 4988 17332
rect 4943 17292 4988 17320
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 12575 17323 12633 17329
rect 12575 17320 12587 17323
rect 8904 17292 12587 17320
rect 8904 17280 8910 17292
rect 12575 17289 12587 17292
rect 12621 17289 12633 17323
rect 12575 17283 12633 17289
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 13078 17320 13084 17332
rect 13035 17292 13084 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 2130 17212 2136 17264
rect 2188 17252 2194 17264
rect 4295 17255 4353 17261
rect 2188 17224 4154 17252
rect 2188 17212 2194 17224
rect 2590 17144 2596 17196
rect 2648 17184 2654 17196
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 2648 17156 2697 17184
rect 2648 17144 2654 17156
rect 2685 17153 2697 17156
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 4126 17128 4154 17224
rect 4295 17221 4307 17255
rect 4341 17252 4353 17255
rect 10318 17252 10324 17264
rect 4341 17224 10324 17252
rect 4341 17221 4353 17224
rect 4295 17215 4353 17221
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 11698 17252 11704 17264
rect 11659 17224 11704 17252
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 6638 17184 6644 17196
rect 5307 17156 6644 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6972 17156 7205 17184
rect 6972 17144 6978 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7374 17184 7380 17196
rect 7335 17156 7380 17184
rect 7193 17147 7251 17153
rect 4062 17076 4068 17128
rect 4120 17116 4154 17128
rect 4224 17119 4282 17125
rect 4224 17116 4236 17119
rect 4120 17088 4236 17116
rect 4120 17076 4126 17088
rect 4224 17085 4236 17088
rect 4270 17116 4282 17119
rect 4617 17119 4675 17125
rect 4617 17116 4629 17119
rect 4270 17088 4629 17116
rect 4270 17085 4282 17088
rect 4224 17079 4282 17085
rect 4617 17085 4629 17088
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6178 17116 6184 17128
rect 5960 17088 6184 17116
rect 5960 17076 5966 17088
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 1394 17008 1400 17060
rect 1452 17048 1458 17060
rect 1857 17051 1915 17057
rect 1857 17048 1869 17051
rect 1452 17020 1869 17048
rect 1452 17008 1458 17020
rect 1857 17017 1869 17020
rect 1903 17048 1915 17051
rect 2409 17051 2467 17057
rect 2409 17048 2421 17051
rect 1903 17020 2421 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 2409 17017 2421 17020
rect 2455 17017 2467 17051
rect 2409 17011 2467 17017
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17017 2559 17051
rect 2501 17011 2559 17017
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 2516 16980 2544 17011
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 5408 17020 5453 17048
rect 5408 17008 5414 17020
rect 6086 17008 6092 17060
rect 6144 17048 6150 17060
rect 6549 17051 6607 17057
rect 6549 17048 6561 17051
rect 6144 17020 6561 17048
rect 6144 17008 6150 17020
rect 6549 17017 6561 17020
rect 6595 17048 6607 17051
rect 6822 17048 6828 17060
rect 6595 17020 6828 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 7208 17048 7236 17147
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 9306 17184 9312 17196
rect 9263 17156 9312 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10468 17156 11069 17184
rect 10468 17144 10474 17156
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12504 17119 12562 17125
rect 12504 17116 12516 17119
rect 12032 17088 12516 17116
rect 12032 17076 12038 17088
rect 12504 17085 12516 17088
rect 12550 17116 12562 17119
rect 13004 17116 13032 17283
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 13630 17320 13636 17332
rect 13591 17292 13636 17320
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 12550 17088 13032 17116
rect 13449 17119 13507 17125
rect 12550 17085 12562 17088
rect 12504 17079 12562 17085
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 7466 17048 7472 17060
rect 7208 17020 7472 17048
rect 7466 17008 7472 17020
rect 7524 17048 7530 17060
rect 7698 17051 7756 17057
rect 7698 17048 7710 17051
rect 7524 17020 7710 17048
rect 7524 17008 7530 17020
rect 7698 17017 7710 17020
rect 7744 17017 7756 17051
rect 7698 17011 7756 17017
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8573 17051 8631 17057
rect 8573 17048 8585 17051
rect 7892 17020 8585 17048
rect 7892 17008 7898 17020
rect 8573 17017 8585 17020
rect 8619 17017 8631 17051
rect 8573 17011 8631 17017
rect 9309 17051 9367 17057
rect 9309 17017 9321 17051
rect 9355 17017 9367 17051
rect 9858 17048 9864 17060
rect 9771 17020 9864 17048
rect 9309 17011 9367 17017
rect 2372 16952 2544 16980
rect 2372 16940 2378 16952
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 3329 16983 3387 16989
rect 3329 16980 3341 16983
rect 3200 16952 3341 16980
rect 3200 16940 3206 16952
rect 3329 16949 3341 16952
rect 3375 16949 3387 16983
rect 3329 16943 3387 16949
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4982 16980 4988 16992
rect 4304 16952 4988 16980
rect 4304 16940 4310 16952
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6181 16983 6239 16989
rect 6181 16980 6193 16983
rect 6052 16952 6193 16980
rect 6052 16940 6058 16952
rect 6181 16949 6193 16952
rect 6227 16949 6239 16983
rect 8294 16980 8300 16992
rect 8255 16952 8300 16980
rect 6181 16943 6239 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8478 16940 8484 16992
rect 8536 16980 8542 16992
rect 9033 16983 9091 16989
rect 9033 16980 9045 16983
rect 8536 16952 9045 16980
rect 8536 16940 8542 16952
rect 9033 16949 9045 16952
rect 9079 16980 9091 16983
rect 9324 16980 9352 17011
rect 9858 17008 9864 17020
rect 9916 17048 9922 17060
rect 10410 17048 10416 17060
rect 9916 17020 10416 17048
rect 9916 17008 9922 17020
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 10594 17008 10600 17060
rect 10652 17048 10658 17060
rect 10781 17051 10839 17057
rect 10781 17048 10793 17051
rect 10652 17020 10793 17048
rect 10652 17008 10658 17020
rect 10781 17017 10793 17020
rect 10827 17017 10839 17051
rect 10781 17011 10839 17017
rect 10873 17051 10931 17057
rect 10873 17017 10885 17051
rect 10919 17017 10931 17051
rect 10873 17011 10931 17017
rect 9950 16980 9956 16992
rect 9079 16952 9956 16980
rect 9079 16949 9091 16952
rect 9033 16943 9091 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 10134 16980 10140 16992
rect 10095 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10502 16980 10508 16992
rect 10463 16952 10508 16980
rect 10502 16940 10508 16952
rect 10560 16980 10566 16992
rect 10888 16980 10916 17011
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 13464 17048 13492 17079
rect 14001 17051 14059 17057
rect 14001 17048 14013 17051
rect 11020 17020 14013 17048
rect 11020 17008 11026 17020
rect 14001 17017 14013 17020
rect 14047 17017 14059 17051
rect 14001 17011 14059 17017
rect 10560 16952 10916 16980
rect 10560 16940 10566 16952
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 1394 16776 1400 16788
rect 1355 16748 1400 16776
rect 1394 16736 1400 16748
rect 1452 16736 1458 16788
rect 7466 16776 7472 16788
rect 7427 16748 7472 16776
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8573 16779 8631 16785
rect 8573 16745 8585 16779
rect 8619 16776 8631 16779
rect 10134 16776 10140 16788
rect 8619 16748 10140 16776
rect 8619 16745 8631 16748
rect 8573 16739 8631 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10594 16736 10600 16788
rect 10652 16776 10658 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 10652 16748 10701 16776
rect 10652 16736 10658 16748
rect 10689 16745 10701 16748
rect 10735 16776 10747 16779
rect 10735 16748 12020 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 2593 16711 2651 16717
rect 2593 16708 2605 16711
rect 2363 16680 2605 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 2593 16677 2605 16680
rect 2639 16708 2651 16711
rect 3142 16708 3148 16720
rect 2639 16680 3148 16708
rect 2639 16677 2651 16680
rect 2593 16671 2651 16677
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 4246 16708 4252 16720
rect 4207 16680 4252 16708
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 5902 16708 5908 16720
rect 5500 16680 5908 16708
rect 5500 16668 5506 16680
rect 5902 16668 5908 16680
rect 5960 16668 5966 16720
rect 5997 16711 6055 16717
rect 5997 16677 6009 16711
rect 6043 16708 6055 16711
rect 6086 16708 6092 16720
rect 6043 16680 6092 16708
rect 6043 16677 6055 16680
rect 5997 16671 6055 16677
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 7484 16708 7512 16736
rect 7974 16711 8032 16717
rect 7974 16708 7986 16711
rect 7484 16680 7986 16708
rect 7974 16677 7986 16680
rect 8020 16677 8032 16711
rect 7974 16671 8032 16677
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 9858 16708 9864 16720
rect 8352 16680 9864 16708
rect 8352 16668 8358 16680
rect 9858 16668 9864 16680
rect 9916 16668 9922 16720
rect 9950 16668 9956 16720
rect 10008 16708 10014 16720
rect 11425 16711 11483 16717
rect 11425 16708 11437 16711
rect 10008 16680 11437 16708
rect 10008 16668 10014 16680
rect 11425 16677 11437 16680
rect 11471 16708 11483 16711
rect 11698 16708 11704 16720
rect 11471 16680 11704 16708
rect 11471 16677 11483 16680
rect 11425 16671 11483 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 11992 16717 12020 16748
rect 11977 16711 12035 16717
rect 11977 16677 11989 16711
rect 12023 16677 12035 16711
rect 11977 16671 12035 16677
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 6696 16612 6929 16640
rect 6696 16600 6702 16612
rect 6917 16609 6929 16612
rect 6963 16640 6975 16643
rect 9398 16640 9404 16652
rect 6963 16612 9404 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2501 16575 2559 16581
rect 2501 16572 2513 16575
rect 2188 16544 2513 16572
rect 2188 16532 2194 16544
rect 2501 16541 2513 16544
rect 2547 16572 2559 16575
rect 2547 16544 3188 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 3053 16507 3111 16513
rect 3053 16504 3065 16507
rect 2648 16476 3065 16504
rect 2648 16464 2654 16476
rect 3053 16473 3065 16476
rect 3099 16473 3111 16507
rect 3160 16504 3188 16544
rect 4154 16532 4160 16584
rect 4212 16572 4218 16584
rect 4798 16572 4804 16584
rect 4212 16544 4257 16572
rect 4759 16544 4804 16572
rect 4212 16532 4218 16544
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 6178 16572 6184 16584
rect 6139 16544 6184 16572
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 7653 16575 7711 16581
rect 7653 16541 7665 16575
rect 7699 16572 7711 16575
rect 8570 16572 8576 16584
rect 7699 16544 8576 16572
rect 7699 16541 7711 16544
rect 7653 16535 7711 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 9769 16575 9827 16581
rect 8680 16544 9444 16572
rect 4816 16504 4844 16532
rect 3160 16476 4844 16504
rect 3053 16467 3111 16473
rect 4890 16464 4896 16516
rect 4948 16504 4954 16516
rect 8680 16504 8708 16544
rect 4948 16476 5672 16504
rect 4948 16464 4954 16476
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 1857 16439 1915 16445
rect 1857 16436 1869 16439
rect 1636 16408 1869 16436
rect 1636 16396 1642 16408
rect 1857 16405 1869 16408
rect 1903 16405 1915 16439
rect 3418 16436 3424 16448
rect 3379 16408 3424 16436
rect 1857 16399 1915 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 5258 16436 5264 16448
rect 5219 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5644 16445 5672 16476
rect 6748 16476 8708 16504
rect 5629 16439 5687 16445
rect 5629 16405 5641 16439
rect 5675 16436 5687 16439
rect 6748 16436 6776 16476
rect 5675 16408 6776 16436
rect 9217 16439 9275 16445
rect 5675 16405 5687 16408
rect 5629 16399 5687 16405
rect 9217 16405 9229 16439
rect 9263 16436 9275 16439
rect 9306 16436 9312 16448
rect 9263 16408 9312 16436
rect 9263 16405 9275 16408
rect 9217 16399 9275 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9416 16436 9444 16544
rect 9769 16541 9781 16575
rect 9815 16541 9827 16575
rect 10410 16572 10416 16584
rect 10371 16544 10416 16572
rect 9769 16535 9827 16541
rect 9784 16504 9812 16535
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11379 16544 12296 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 10778 16504 10784 16516
rect 9784 16476 10784 16504
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 12268 16448 12296 16544
rect 12066 16436 12072 16448
rect 9416 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12250 16396 12256 16448
rect 12308 16436 12314 16448
rect 12943 16439 13001 16445
rect 12943 16436 12955 16439
rect 12308 16408 12955 16436
rect 12308 16396 12314 16408
rect 12943 16405 12955 16408
rect 12989 16405 13001 16439
rect 12943 16399 13001 16405
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 4246 16232 4252 16244
rect 3896 16204 4154 16232
rect 4207 16204 4252 16232
rect 2041 16167 2099 16173
rect 2041 16133 2053 16167
rect 2087 16164 2099 16167
rect 3896 16164 3924 16204
rect 2087 16136 3924 16164
rect 4126 16164 4154 16204
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 5902 16192 5908 16244
rect 5960 16232 5966 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5960 16204 6193 16232
rect 5960 16192 5966 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 6181 16195 6239 16201
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7466 16232 7472 16244
rect 7331 16204 7472 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8478 16232 8484 16244
rect 8343 16204 8484 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10502 16232 10508 16244
rect 10091 16204 10508 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11330 16232 11336 16244
rect 11291 16204 11336 16232
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 11698 16232 11704 16244
rect 11659 16204 11704 16232
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12161 16235 12219 16241
rect 12161 16201 12173 16235
rect 12207 16232 12219 16235
rect 12250 16232 12256 16244
rect 12207 16204 12256 16232
rect 12207 16201 12219 16204
rect 12161 16195 12219 16201
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 5920 16164 5948 16192
rect 4126 16136 5948 16164
rect 7484 16164 7512 16192
rect 8941 16167 8999 16173
rect 8941 16164 8953 16167
rect 7484 16136 8953 16164
rect 2087 16133 2099 16136
rect 2041 16127 2099 16133
rect 8941 16133 8953 16136
rect 8987 16164 8999 16167
rect 8987 16136 9260 16164
rect 8987 16133 8999 16136
rect 8941 16127 8999 16133
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 3418 16096 3424 16108
rect 1535 16068 3424 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 4798 16056 4804 16108
rect 4856 16096 4862 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 4856 16068 5089 16096
rect 4856 16056 4862 16068
rect 5077 16065 5089 16068
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 8018 16056 8024 16108
rect 8076 16096 8082 16108
rect 9122 16096 9128 16108
rect 8076 16068 9128 16096
rect 8076 16056 8082 16068
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9232 16096 9260 16136
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 11011 16167 11069 16173
rect 11011 16164 11023 16167
rect 9364 16136 11023 16164
rect 9364 16124 9370 16136
rect 11011 16133 11023 16136
rect 11057 16133 11069 16167
rect 11011 16127 11069 16133
rect 9490 16096 9496 16108
rect 9232 16068 9496 16096
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9916 16068 10333 16096
rect 9916 16056 9922 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2866 16028 2872 16040
rect 2547 16000 2872 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2866 15988 2872 16000
rect 2924 16028 2930 16040
rect 2961 16031 3019 16037
rect 2961 16028 2973 16031
rect 2924 16000 2973 16028
rect 2924 15988 2930 16000
rect 2961 15997 2973 16000
rect 3007 15997 3019 16031
rect 2961 15991 3019 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 6687 16000 7389 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7377 15997 7389 16000
rect 7423 16028 7435 16031
rect 9950 16028 9956 16040
rect 7423 16000 9956 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10940 16031 10998 16037
rect 10940 15997 10952 16031
rect 10986 16028 10998 16031
rect 11330 16028 11336 16040
rect 10986 16000 11336 16028
rect 10986 15997 10998 16000
rect 10940 15991 10998 15997
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 1578 15960 1584 15972
rect 1539 15932 1584 15960
rect 1578 15920 1584 15932
rect 1636 15920 1642 15972
rect 3282 15963 3340 15969
rect 3282 15960 3294 15963
rect 2792 15932 3294 15960
rect 2314 15852 2320 15904
rect 2372 15892 2378 15904
rect 2792 15901 2820 15932
rect 3282 15929 3294 15932
rect 3328 15929 3340 15963
rect 4798 15960 4804 15972
rect 4759 15932 4804 15960
rect 3282 15923 3340 15929
rect 4798 15920 4804 15932
rect 4856 15920 4862 15972
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15929 4951 15963
rect 4893 15923 4951 15929
rect 2777 15895 2835 15901
rect 2777 15892 2789 15895
rect 2372 15864 2789 15892
rect 2372 15852 2378 15864
rect 2777 15861 2789 15864
rect 2823 15861 2835 15895
rect 2777 15855 2835 15861
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 3108 15864 3893 15892
rect 3108 15852 3114 15864
rect 3881 15861 3893 15864
rect 3927 15892 3939 15895
rect 4246 15892 4252 15904
rect 3927 15864 4252 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4430 15852 4436 15904
rect 4488 15892 4494 15904
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4488 15864 4537 15892
rect 4488 15852 4494 15864
rect 4525 15861 4537 15864
rect 4571 15892 4583 15895
rect 4908 15892 4936 15923
rect 7466 15920 7472 15972
rect 7524 15960 7530 15972
rect 7698 15963 7756 15969
rect 7698 15960 7710 15963
rect 7524 15932 7710 15960
rect 7524 15920 7530 15932
rect 7698 15929 7710 15932
rect 7744 15929 7756 15963
rect 7698 15923 7756 15929
rect 8110 15920 8116 15972
rect 8168 15960 8174 15972
rect 9490 15969 9496 15972
rect 9487 15960 9496 15969
rect 8168 15932 9352 15960
rect 9451 15932 9496 15960
rect 8168 15920 8174 15932
rect 4571 15864 4936 15892
rect 5905 15895 5963 15901
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 5905 15861 5917 15895
rect 5951 15892 5963 15895
rect 6086 15892 6092 15904
rect 5951 15864 6092 15892
rect 5951 15861 5963 15864
rect 5905 15855 5963 15861
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 8570 15892 8576 15904
rect 8531 15864 8576 15892
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 9324 15892 9352 15932
rect 9487 15923 9496 15932
rect 9490 15920 9496 15923
rect 9548 15920 9554 15972
rect 12802 15892 12808 15904
rect 9324 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3142 15688 3148 15700
rect 3103 15660 3148 15688
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 6411 15691 6469 15697
rect 6411 15688 6423 15691
rect 3476 15660 6423 15688
rect 3476 15648 3482 15660
rect 6411 15657 6423 15660
rect 6457 15657 6469 15691
rect 8846 15688 8852 15700
rect 8759 15660 8852 15688
rect 6411 15651 6469 15657
rect 8846 15648 8852 15660
rect 8904 15688 8910 15700
rect 11379 15691 11437 15697
rect 11379 15688 11391 15691
rect 8904 15660 11391 15688
rect 8904 15648 8910 15660
rect 11379 15657 11391 15660
rect 11425 15657 11437 15691
rect 11379 15651 11437 15657
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12391 15691 12449 15697
rect 12391 15688 12403 15691
rect 12124 15660 12403 15688
rect 12124 15648 12130 15660
rect 12391 15657 12403 15660
rect 12437 15657 12449 15691
rect 12391 15651 12449 15657
rect 2314 15580 2320 15632
rect 2372 15620 2378 15632
rect 2546 15623 2604 15629
rect 2546 15620 2558 15623
rect 2372 15592 2558 15620
rect 2372 15580 2378 15592
rect 2546 15589 2558 15592
rect 2592 15620 2604 15623
rect 4246 15620 4252 15632
rect 2592 15592 4252 15620
rect 2592 15589 2604 15592
rect 2546 15583 2604 15589
rect 4246 15580 4252 15592
rect 4304 15620 4310 15632
rect 4846 15623 4904 15629
rect 4846 15620 4858 15623
rect 4304 15592 4858 15620
rect 4304 15580 4310 15592
rect 4846 15589 4858 15592
rect 4892 15589 4904 15623
rect 4846 15583 4904 15589
rect 4982 15580 4988 15632
rect 5040 15620 5046 15632
rect 6825 15623 6883 15629
rect 6825 15620 6837 15623
rect 5040 15592 6837 15620
rect 5040 15580 5046 15592
rect 6825 15589 6837 15592
rect 6871 15589 6883 15623
rect 6825 15583 6883 15589
rect 7466 15580 7472 15632
rect 7524 15620 7530 15632
rect 7790 15623 7848 15629
rect 7790 15620 7802 15623
rect 7524 15592 7802 15620
rect 7524 15580 7530 15592
rect 7790 15589 7802 15592
rect 7836 15589 7848 15623
rect 9122 15620 9128 15632
rect 9083 15592 9128 15620
rect 7790 15583 7848 15589
rect 9122 15580 9128 15592
rect 9180 15580 9186 15632
rect 9858 15620 9864 15632
rect 9819 15592 9864 15620
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 10410 15620 10416 15632
rect 10371 15592 10416 15620
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 11146 15580 11152 15632
rect 11204 15620 11210 15632
rect 11204 15592 12363 15620
rect 11204 15580 11210 15592
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 1636 15524 5457 15552
rect 1636 15512 1642 15524
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2774 15484 2780 15496
rect 2464 15456 2780 15484
rect 2464 15444 2470 15456
rect 2774 15444 2780 15456
rect 2832 15484 2838 15496
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 2832 15456 3433 15484
rect 2832 15444 2838 15456
rect 3421 15453 3433 15456
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15453 4583 15487
rect 5460 15484 5488 15515
rect 5718 15512 5724 15564
rect 5776 15552 5782 15564
rect 6270 15552 6276 15564
rect 6328 15561 6334 15564
rect 6328 15555 6366 15561
rect 5776 15524 6276 15552
rect 5776 15512 5782 15524
rect 6270 15512 6276 15524
rect 6354 15521 6366 15555
rect 11238 15552 11244 15564
rect 11199 15524 11244 15552
rect 6328 15515 6366 15521
rect 6328 15512 6334 15515
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 12335 15561 12363 15592
rect 12320 15555 12378 15561
rect 12320 15521 12332 15555
rect 12366 15552 12378 15555
rect 12618 15552 12624 15564
rect 12366 15524 12624 15552
rect 12366 15521 12378 15524
rect 12320 15515 12378 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 7469 15487 7527 15493
rect 5460 15456 7420 15484
rect 4525 15447 4583 15453
rect 4540 15360 4568 15447
rect 4890 15376 4896 15428
rect 4948 15416 4954 15428
rect 5813 15419 5871 15425
rect 5813 15416 5825 15419
rect 4948 15388 5825 15416
rect 4948 15376 4954 15388
rect 5813 15385 5825 15388
rect 5859 15416 5871 15419
rect 6914 15416 6920 15428
rect 5859 15388 6920 15416
rect 5859 15385 5871 15388
rect 5813 15379 5871 15385
rect 6914 15376 6920 15388
rect 6972 15376 6978 15428
rect 7392 15416 7420 15456
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8202 15484 8208 15496
rect 7515 15456 8208 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10226 15416 10232 15428
rect 7392 15388 10232 15416
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 3510 15308 3516 15360
rect 3568 15348 3574 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 3568 15320 3801 15348
rect 3568 15308 3574 15320
rect 3789 15317 3801 15320
rect 3835 15348 3847 15351
rect 4154 15348 4160 15360
rect 3835 15320 4160 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4433 15351 4491 15357
rect 4433 15317 4445 15351
rect 4479 15348 4491 15351
rect 4522 15348 4528 15360
rect 4479 15320 4528 15348
rect 4479 15317 4491 15320
rect 4433 15311 4491 15317
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 8389 15351 8447 15357
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 8662 15348 8668 15360
rect 8435 15320 8668 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10778 15348 10784 15360
rect 9456 15320 10784 15348
rect 9456 15308 9462 15320
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 2314 15144 2320 15156
rect 2275 15116 2320 15144
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5316 15116 5825 15144
rect 5316 15104 5322 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 5813 15107 5871 15113
rect 6270 15104 6276 15116
rect 6328 15144 6334 15156
rect 8110 15144 8116 15156
rect 6328 15116 8116 15144
rect 6328 15104 6334 15116
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 8662 15144 8668 15156
rect 8623 15116 8668 15144
rect 8662 15104 8668 15116
rect 8720 15144 8726 15156
rect 9858 15144 9864 15156
rect 8720 15116 9864 15144
rect 8720 15104 8726 15116
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 10226 15144 10232 15156
rect 10187 15116 10232 15144
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 12618 15144 12624 15156
rect 12579 15116 12624 15144
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 4246 15036 4252 15088
rect 4304 15076 4310 15088
rect 4433 15079 4491 15085
rect 4433 15076 4445 15079
rect 4304 15048 4445 15076
rect 4304 15036 4310 15048
rect 4433 15045 4445 15048
rect 4479 15076 4491 15079
rect 4801 15079 4859 15085
rect 4801 15076 4813 15079
rect 4479 15048 4813 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4801 15045 4813 15048
rect 4847 15076 4859 15079
rect 5166 15076 5172 15088
rect 4847 15048 5172 15076
rect 4847 15045 4859 15048
rect 4801 15039 4859 15045
rect 5166 15036 5172 15048
rect 5224 15076 5230 15088
rect 7466 15076 7472 15088
rect 5224 15048 7472 15076
rect 5224 15036 5230 15048
rect 7466 15036 7472 15048
rect 7524 15076 7530 15088
rect 7837 15079 7895 15085
rect 7837 15076 7849 15079
rect 7524 15048 7849 15076
rect 7524 15036 7530 15048
rect 7837 15045 7849 15048
rect 7883 15045 7895 15079
rect 7837 15039 7895 15045
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 8904 15048 8984 15076
rect 8904 15036 8910 15048
rect 4890 15008 4896 15020
rect 4851 14980 4896 15008
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 8956 15017 8984 15048
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 11238 15076 11244 15088
rect 9732 15048 11244 15076
rect 9732 15036 9738 15048
rect 11238 15036 11244 15048
rect 11296 15076 11302 15088
rect 11425 15079 11483 15085
rect 11425 15076 11437 15079
rect 11296 15048 11437 15076
rect 11296 15036 11302 15048
rect 11425 15045 11437 15048
rect 11471 15045 11483 15079
rect 11425 15039 11483 15045
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 10594 15008 10600 15020
rect 9631 14980 10600 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 10778 15008 10784 15020
rect 10739 14980 10784 15008
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14940 1639 14943
rect 1670 14940 1676 14952
rect 1627 14912 1676 14940
rect 1627 14909 1639 14912
rect 1581 14903 1639 14909
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 3418 14940 3424 14952
rect 3379 14912 3424 14940
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 1397 14875 1455 14881
rect 1397 14841 1409 14875
rect 1443 14872 1455 14875
rect 1854 14872 1860 14884
rect 1443 14844 1860 14872
rect 1443 14841 1455 14844
rect 1397 14835 1455 14841
rect 1854 14832 1860 14844
rect 1912 14832 1918 14884
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 2498 14872 2504 14884
rect 1995 14844 2504 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2498 14832 2504 14844
rect 2556 14832 2562 14884
rect 2685 14875 2743 14881
rect 2685 14841 2697 14875
rect 2731 14872 2743 14875
rect 2958 14872 2964 14884
rect 2731 14844 2964 14872
rect 2731 14841 2743 14844
rect 2685 14835 2743 14841
rect 2958 14832 2964 14844
rect 3016 14872 3022 14884
rect 3620 14872 3648 14903
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 4212 14912 6837 14940
rect 4212 14900 4218 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7190 14940 7196 14952
rect 6871 14912 7196 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 7466 14940 7472 14952
rect 7423 14912 7472 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 5810 14872 5816 14884
rect 3016 14844 3648 14872
rect 3712 14844 5816 14872
rect 3016 14832 3022 14844
rect 2866 14804 2872 14816
rect 2827 14776 2872 14804
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3712 14804 3740 14844
rect 5810 14832 5816 14844
rect 5868 14872 5874 14884
rect 7650 14872 7656 14884
rect 5868 14844 7656 14872
rect 5868 14832 5874 14844
rect 7650 14832 7656 14844
rect 7708 14832 7714 14884
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 9033 14875 9091 14881
rect 9033 14872 9045 14875
rect 8720 14844 9045 14872
rect 8720 14832 8726 14844
rect 9033 14841 9045 14844
rect 9079 14841 9091 14875
rect 9033 14835 9091 14841
rect 10318 14832 10324 14884
rect 10376 14872 10382 14884
rect 10505 14875 10563 14881
rect 10505 14872 10517 14875
rect 10376 14844 10517 14872
rect 10376 14832 10382 14844
rect 10505 14841 10517 14844
rect 10551 14841 10563 14875
rect 10505 14835 10563 14841
rect 10597 14875 10655 14881
rect 10597 14841 10609 14875
rect 10643 14841 10655 14875
rect 10597 14835 10655 14841
rect 3200 14776 3740 14804
rect 3200 14764 3206 14776
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4246 14804 4252 14816
rect 4028 14776 4252 14804
rect 4028 14764 4034 14776
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5261 14807 5319 14813
rect 5261 14804 5273 14807
rect 5224 14776 5273 14804
rect 5224 14764 5230 14776
rect 5261 14773 5273 14776
rect 5307 14773 5319 14807
rect 6914 14804 6920 14816
rect 6875 14776 6920 14804
rect 5261 14767 5319 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10612 14804 10640 14835
rect 10284 14776 10640 14804
rect 10284 14764 10290 14776
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 1535 14603 1593 14609
rect 1535 14569 1547 14603
rect 1581 14600 1593 14603
rect 3510 14600 3516 14612
rect 1581 14572 3516 14600
rect 1581 14569 1593 14572
rect 1535 14563 1593 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4338 14600 4344 14612
rect 4299 14572 4344 14600
rect 4338 14560 4344 14572
rect 4396 14600 4402 14612
rect 5258 14600 5264 14612
rect 4396 14572 5264 14600
rect 4396 14560 4402 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 6086 14600 6092 14612
rect 6047 14572 6092 14600
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 8754 14600 8760 14612
rect 8628 14572 8760 14600
rect 8628 14560 8634 14572
rect 8754 14560 8760 14572
rect 8812 14560 8818 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9766 14600 9772 14612
rect 9539 14572 9772 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10318 14560 10324 14612
rect 10376 14600 10382 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10376 14572 10701 14600
rect 10376 14560 10382 14572
rect 10689 14569 10701 14572
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 3145 14535 3203 14541
rect 3145 14501 3157 14535
rect 3191 14532 3203 14535
rect 4430 14532 4436 14544
rect 3191 14504 4436 14532
rect 3191 14501 3203 14504
rect 3145 14495 3203 14501
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 5166 14492 5172 14544
rect 5224 14532 5230 14544
rect 5490 14535 5548 14541
rect 5490 14532 5502 14535
rect 5224 14504 5502 14532
rect 5224 14492 5230 14504
rect 5490 14501 5502 14504
rect 5536 14532 5548 14535
rect 5718 14532 5724 14544
rect 5536 14504 5724 14532
rect 5536 14501 5548 14504
rect 5490 14495 5548 14501
rect 5718 14492 5724 14504
rect 5776 14492 5782 14544
rect 7653 14535 7711 14541
rect 7653 14501 7665 14535
rect 7699 14532 7711 14535
rect 8202 14532 8208 14544
rect 7699 14504 8208 14532
rect 7699 14501 7711 14504
rect 7653 14495 7711 14501
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 1464 14467 1522 14473
rect 1464 14433 1476 14467
rect 1510 14464 1522 14467
rect 2038 14464 2044 14476
rect 1510 14436 2044 14464
rect 1510 14433 1522 14436
rect 1464 14427 1522 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2406 14424 2412 14476
rect 2464 14464 2470 14476
rect 2501 14467 2559 14473
rect 2501 14464 2513 14467
rect 2464 14436 2513 14464
rect 2464 14424 2470 14436
rect 2501 14433 2513 14436
rect 2547 14464 2559 14467
rect 3050 14464 3056 14476
rect 2547 14436 3056 14464
rect 2547 14433 2559 14436
rect 2501 14427 2559 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3418 14464 3424 14476
rect 3379 14436 3424 14464
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4157 14467 4215 14473
rect 4157 14464 4169 14467
rect 4028 14436 4169 14464
rect 4028 14424 4034 14436
rect 4157 14433 4169 14436
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6880 14436 6929 14464
rect 6880 14424 6886 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 1854 14356 1860 14408
rect 1912 14396 1918 14408
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1912 14368 1961 14396
rect 1912 14356 1918 14368
rect 1949 14365 1961 14368
rect 1995 14396 2007 14399
rect 2682 14396 2688 14408
rect 1995 14368 2688 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 3436 14396 3464 14424
rect 5166 14396 5172 14408
rect 2740 14368 3464 14396
rect 5127 14368 5172 14396
rect 2740 14356 2746 14368
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 6932 14328 6960 14427
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7064 14436 7389 14464
rect 7064 14424 7070 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8516 14467 8574 14473
rect 8516 14464 8528 14467
rect 8168 14436 8528 14464
rect 8168 14424 8174 14436
rect 8516 14433 8528 14436
rect 8562 14433 8574 14467
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 8516 14427 8574 14433
rect 9600 14436 9689 14464
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 8846 14396 8852 14408
rect 7248 14368 8852 14396
rect 7248 14356 7254 14368
rect 8846 14356 8852 14368
rect 8904 14396 8910 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8904 14368 8953 14396
rect 8904 14356 8910 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 7926 14328 7932 14340
rect 6932 14300 7932 14328
rect 7208 14272 7236 14300
rect 7926 14288 7932 14300
rect 7984 14328 7990 14340
rect 9600 14328 9628 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 10134 14464 10140 14476
rect 10095 14436 10140 14464
rect 9677 14427 9735 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 9674 14328 9680 14340
rect 7984 14300 9680 14328
rect 7984 14288 7990 14300
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 2317 14263 2375 14269
rect 2317 14260 2329 14263
rect 2280 14232 2329 14260
rect 2280 14220 2286 14232
rect 2317 14229 2329 14232
rect 2363 14260 2375 14263
rect 2866 14260 2872 14272
rect 2363 14232 2872 14260
rect 2363 14229 2375 14232
rect 2317 14223 2375 14229
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 4798 14260 4804 14272
rect 4759 14232 4804 14260
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 7190 14220 7196 14272
rect 7248 14220 7254 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8619 14263 8677 14269
rect 8619 14260 8631 14263
rect 8536 14232 8631 14260
rect 8536 14220 8542 14232
rect 8619 14229 8631 14232
rect 8665 14229 8677 14263
rect 8619 14223 8677 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 2682 14056 2688 14068
rect 2643 14028 2688 14056
rect 2682 14016 2688 14028
rect 2740 14016 2746 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 4488 14028 4629 14056
rect 4488 14016 4494 14028
rect 4617 14025 4629 14028
rect 4663 14056 4675 14059
rect 4982 14056 4988 14068
rect 4663 14028 4988 14056
rect 4663 14025 4675 14028
rect 4617 14019 4675 14025
rect 4982 14016 4988 14028
rect 5040 14056 5046 14068
rect 5350 14056 5356 14068
rect 5040 14028 5356 14056
rect 5040 14016 5046 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5718 14056 5724 14068
rect 5500 14028 5724 14056
rect 5500 14016 5506 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14056 6515 14059
rect 7466 14056 7472 14068
rect 6503 14028 7472 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 2038 13988 2044 14000
rect 1951 13960 2044 13988
rect 2038 13948 2044 13960
rect 2096 13988 2102 14000
rect 3142 13988 3148 14000
rect 2096 13960 3148 13988
rect 2096 13948 2102 13960
rect 3142 13948 3148 13960
rect 3200 13948 3206 14000
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 5626 13988 5632 14000
rect 4856 13960 5632 13988
rect 4856 13948 4862 13960
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3476 13892 3525 13920
rect 3476 13880 3482 13892
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1670 13852 1676 13864
rect 1443 13824 1676 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1670 13812 1676 13824
rect 1728 13852 1734 13864
rect 2130 13852 2136 13864
rect 1728 13824 2136 13852
rect 1728 13812 1734 13824
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 3602 13852 3608 13864
rect 3563 13824 3608 13852
rect 2869 13815 2927 13821
rect 2774 13744 2780 13796
rect 2832 13784 2838 13796
rect 2884 13784 2912 13815
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 5000 13861 5028 13960
rect 5626 13948 5632 13960
rect 5684 13988 5690 14000
rect 7282 13988 7288 14000
rect 5684 13960 7288 13988
rect 5684 13948 5690 13960
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 7006 13920 7012 13932
rect 6196 13892 7012 13920
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13821 5043 13855
rect 4985 13815 5043 13821
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5350 13852 5356 13864
rect 5307 13824 5356 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 6196 13796 6224 13892
rect 6932 13861 6960 13892
rect 7006 13880 7012 13892
rect 7064 13880 7070 13932
rect 7386 13861 7414 14028
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7926 14056 7932 14068
rect 7887 14028 7932 14056
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 8168 14028 8309 14056
rect 8168 14016 8174 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 8297 14019 8355 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10091 14059 10149 14065
rect 10091 14056 10103 14059
rect 9824 14028 10103 14056
rect 9824 14016 9830 14028
rect 10091 14025 10103 14028
rect 10137 14025 10149 14059
rect 10091 14019 10149 14025
rect 7944 13920 7972 14016
rect 7944 13892 8432 13920
rect 8404 13861 8432 13892
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 9548 13892 10425 13920
rect 9548 13880 9554 13892
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13821 8447 13855
rect 8846 13852 8852 13864
rect 8807 13824 8852 13852
rect 8389 13815 8447 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 10035 13861 10063 13892
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 10413 13883 10471 13889
rect 10004 13855 10063 13861
rect 10004 13821 10016 13855
rect 10050 13824 10063 13855
rect 10050 13821 10062 13824
rect 10004 13815 10062 13821
rect 3418 13784 3424 13796
rect 2832 13756 3424 13784
rect 2832 13744 2838 13756
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 6178 13784 6184 13796
rect 4172 13756 6184 13784
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 3970 13716 3976 13728
rect 3568 13688 3976 13716
rect 3568 13676 3574 13688
rect 3970 13676 3976 13688
rect 4028 13716 4034 13728
rect 4172 13725 4200 13756
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 4028 13688 4169 13716
rect 4028 13676 4034 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4798 13716 4804 13728
rect 4759 13688 4804 13716
rect 4157 13679 4215 13685
rect 4798 13676 4804 13688
rect 4856 13676 4862 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 5408 13688 6469 13716
rect 5408 13676 5414 13688
rect 6457 13685 6469 13688
rect 6503 13716 6515 13719
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6503 13688 6561 13716
rect 6503 13685 6515 13688
rect 6457 13679 6515 13685
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6549 13679 6607 13685
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 2406 13512 2412 13524
rect 2367 13484 2412 13512
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 3108 13484 3157 13512
rect 3108 13472 3114 13484
rect 3145 13481 3157 13484
rect 3191 13512 3203 13515
rect 3234 13512 3240 13524
rect 3191 13484 3240 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3418 13512 3424 13524
rect 3379 13484 3424 13512
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4304 13484 4537 13512
rect 4304 13472 4310 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 5166 13512 5172 13524
rect 5127 13484 5172 13512
rect 4525 13475 4583 13481
rect 2222 13444 2228 13456
rect 1964 13416 2228 13444
rect 1964 13385 1992 13416
rect 2222 13404 2228 13416
rect 2280 13444 2286 13456
rect 3326 13444 3332 13456
rect 2280 13416 3332 13444
rect 2280 13404 2286 13416
rect 3326 13404 3332 13416
rect 3384 13404 3390 13456
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13345 2007 13379
rect 1949 13339 2007 13345
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 2648 13348 2973 13376
rect 2648 13336 2654 13348
rect 2961 13345 2973 13348
rect 3007 13376 3019 13379
rect 4264 13376 4292 13472
rect 4540 13444 4568 13475
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6052 13484 6285 13512
rect 6052 13472 6058 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 7009 13515 7067 13521
rect 7009 13481 7021 13515
rect 7055 13512 7067 13515
rect 7190 13512 7196 13524
rect 7055 13484 7196 13512
rect 7055 13481 7067 13484
rect 7009 13475 7067 13481
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 10134 13512 10140 13524
rect 7340 13484 10140 13512
rect 7340 13472 7346 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 5074 13444 5080 13456
rect 4540 13416 5080 13444
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 5442 13404 5448 13456
rect 5500 13444 5506 13456
rect 5715 13447 5773 13453
rect 5715 13444 5727 13447
rect 5500 13416 5727 13444
rect 5500 13404 5506 13416
rect 5715 13413 5727 13416
rect 5761 13444 5773 13447
rect 5902 13444 5908 13456
rect 5761 13416 5908 13444
rect 5761 13413 5773 13416
rect 5715 13407 5773 13413
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 7926 13404 7932 13456
rect 7984 13444 7990 13456
rect 8205 13447 8263 13453
rect 8205 13444 8217 13447
rect 7984 13416 8217 13444
rect 7984 13404 7990 13416
rect 8205 13413 8217 13416
rect 8251 13413 8263 13447
rect 8205 13407 8263 13413
rect 3007 13348 4292 13376
rect 4341 13379 4399 13385
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4798 13376 4804 13388
rect 4387 13348 4804 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 9712 13379 9770 13385
rect 9712 13376 9724 13379
rect 9640 13348 9724 13376
rect 9640 13336 9646 13348
rect 9712 13345 9724 13348
rect 9758 13376 9770 13379
rect 11974 13376 11980 13388
rect 9758 13348 11980 13376
rect 9758 13345 9770 13348
rect 9712 13339 9770 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3418 13308 3424 13320
rect 2915 13280 3424 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3418 13268 3424 13280
rect 3476 13308 3482 13320
rect 3602 13308 3608 13320
rect 3476 13280 3608 13308
rect 3476 13268 3482 13280
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5350 13308 5356 13320
rect 4764 13280 5212 13308
rect 5311 13280 5356 13308
rect 4764 13268 4770 13280
rect 2133 13243 2191 13249
rect 2133 13209 2145 13243
rect 2179 13240 2191 13243
rect 4982 13240 4988 13252
rect 2179 13212 4988 13240
rect 2179 13209 2191 13212
rect 2133 13203 2191 13209
rect 4982 13200 4988 13212
rect 5040 13200 5046 13252
rect 4798 13172 4804 13184
rect 4759 13144 4804 13172
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 5184 13172 5212 13280
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8846 13308 8852 13320
rect 8159 13280 8852 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8846 13268 8852 13280
rect 8904 13308 8910 13320
rect 9815 13311 9873 13317
rect 9815 13308 9827 13311
rect 8904 13280 9827 13308
rect 8904 13268 8910 13280
rect 9815 13277 9827 13280
rect 9861 13277 9873 13311
rect 9815 13271 9873 13277
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 6880 13212 7297 13240
rect 6880 13200 6886 13212
rect 7285 13209 7297 13212
rect 7331 13209 7343 13243
rect 7285 13203 7343 13209
rect 8665 13243 8723 13249
rect 8665 13209 8677 13243
rect 8711 13240 8723 13243
rect 8754 13240 8760 13252
rect 8711 13212 8760 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 9398 13172 9404 13184
rect 5184 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 2222 12968 2228 12980
rect 2183 12940 2228 12968
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 2590 12968 2596 12980
rect 2551 12940 2596 12968
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 4341 12971 4399 12977
rect 4341 12968 4353 12971
rect 2915 12940 4353 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 4341 12937 4353 12940
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 4525 12971 4583 12977
rect 4525 12968 4537 12971
rect 4488 12940 4537 12968
rect 4488 12928 4494 12940
rect 4525 12937 4537 12940
rect 4571 12937 4583 12971
rect 4525 12931 4583 12937
rect 2406 12860 2412 12912
rect 2464 12900 2470 12912
rect 3881 12903 3939 12909
rect 3881 12900 3893 12903
rect 2464 12872 3893 12900
rect 2464 12860 2470 12872
rect 3881 12869 3893 12872
rect 3927 12900 3939 12903
rect 4154 12900 4160 12912
rect 3927 12872 4160 12900
rect 3927 12869 3939 12872
rect 3881 12863 3939 12869
rect 4154 12860 4160 12872
rect 4212 12900 4218 12912
rect 4212 12872 4476 12900
rect 4212 12860 4218 12872
rect 4448 12844 4476 12872
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 2700 12804 3249 12832
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 2700 12773 2728 12804
rect 3237 12801 3249 12804
rect 3283 12832 3295 12835
rect 3283 12804 4154 12832
rect 3283 12801 3295 12804
rect 3237 12795 3295 12801
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12733 2743 12767
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 2685 12727 2743 12733
rect 3528 12736 3709 12764
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3528 12637 3556 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 4126 12696 4154 12804
rect 4430 12792 4436 12844
rect 4488 12792 4494 12844
rect 4540 12832 4568 12931
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 5408 12940 6193 12968
rect 5408 12928 5414 12940
rect 6181 12937 6193 12940
rect 6227 12968 6239 12971
rect 6914 12968 6920 12980
rect 6227 12940 6920 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 11514 12968 11520 12980
rect 10551 12940 11520 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 5166 12860 5172 12912
rect 5224 12900 5230 12912
rect 5224 12872 5304 12900
rect 5224 12860 5230 12872
rect 5276 12841 5304 12872
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 9582 12900 9588 12912
rect 6788 12872 9588 12900
rect 6788 12860 6794 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 9769 12903 9827 12909
rect 9769 12900 9781 12903
rect 9640 12872 9781 12900
rect 9640 12860 9646 12872
rect 9769 12869 9781 12872
rect 9815 12869 9827 12903
rect 9769 12863 9827 12869
rect 5261 12835 5319 12841
rect 4540 12804 5212 12832
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4890 12764 4896 12776
rect 4387 12736 4896 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 5184 12773 5212 12804
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5718 12832 5724 12844
rect 5261 12795 5319 12801
rect 5362 12804 5724 12832
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12733 5043 12767
rect 4985 12727 5043 12733
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 4249 12699 4307 12705
rect 4249 12696 4261 12699
rect 4126 12668 4261 12696
rect 4249 12665 4261 12668
rect 4295 12696 4307 12699
rect 4522 12696 4528 12708
rect 4295 12668 4528 12696
rect 4295 12665 4307 12668
rect 4249 12659 4307 12665
rect 4522 12656 4528 12668
rect 4580 12696 4586 12708
rect 5000 12696 5028 12727
rect 5362 12696 5390 12804
rect 5718 12792 5724 12804
rect 5776 12832 5782 12844
rect 7834 12832 7840 12844
rect 5776 12804 7840 12832
rect 5776 12792 5782 12804
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 8478 12832 8484 12844
rect 8439 12804 8484 12832
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12832 8818 12844
rect 9674 12832 9680 12844
rect 8812 12804 9680 12832
rect 8812 12792 8818 12804
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 6822 12764 6828 12776
rect 6236 12736 6828 12764
rect 6236 12724 6242 12736
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 10020 12767 10078 12773
rect 10020 12733 10032 12767
rect 10066 12764 10078 12767
rect 10318 12764 10324 12776
rect 10066 12736 10324 12764
rect 10066 12733 10078 12736
rect 10020 12727 10078 12733
rect 7300 12696 7328 12727
rect 10318 12724 10324 12736
rect 10376 12764 10382 12776
rect 10520 12764 10548 12931
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 10376 12736 10548 12764
rect 10376 12724 10382 12736
rect 4580 12668 5390 12696
rect 6564 12668 7328 12696
rect 8573 12699 8631 12705
rect 4580 12656 4586 12668
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 3200 12600 3525 12628
rect 3200 12588 3206 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 5902 12628 5908 12640
rect 5859 12600 5908 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 6564 12637 6592 12668
rect 8573 12665 8585 12699
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6052 12600 6561 12628
rect 6052 12588 6058 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7282 12628 7288 12640
rect 7147 12600 7288 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8076 12600 8217 12628
rect 8076 12588 8082 12600
rect 8205 12597 8217 12600
rect 8251 12628 8263 12631
rect 8588 12628 8616 12659
rect 8251 12600 8616 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10091 12631 10149 12637
rect 10091 12628 10103 12631
rect 9824 12600 10103 12628
rect 9824 12588 9830 12600
rect 10091 12597 10103 12600
rect 10137 12597 10149 12631
rect 10091 12591 10149 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 4580 12396 4629 12424
rect 4580 12384 4586 12396
rect 4617 12393 4629 12396
rect 4663 12393 4675 12427
rect 6822 12424 6828 12436
rect 6783 12396 6828 12424
rect 4617 12387 4675 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 8478 12424 8484 12436
rect 8439 12396 8484 12424
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8846 12424 8852 12436
rect 8807 12396 8852 12424
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 7006 12356 7012 12368
rect 5960 12328 7012 12356
rect 5960 12316 5966 12328
rect 7006 12316 7012 12328
rect 7064 12356 7070 12368
rect 7330 12359 7388 12365
rect 7330 12356 7342 12359
rect 7064 12328 7342 12356
rect 7064 12316 7070 12328
rect 7330 12325 7342 12328
rect 7376 12325 7388 12359
rect 9766 12356 9772 12368
rect 9727 12328 9772 12356
rect 7330 12319 7388 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 9916 12328 9961 12356
rect 9916 12316 9922 12328
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2406 12288 2412 12300
rect 1995 12260 2412 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 2961 12291 3019 12297
rect 2961 12288 2973 12291
rect 2924 12260 2973 12288
rect 2924 12248 2930 12260
rect 2961 12257 2973 12260
rect 3007 12288 3019 12291
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3007 12260 3433 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4706 12288 4712 12300
rect 4479 12260 4712 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5626 12288 5632 12300
rect 5587 12260 5632 12288
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 5994 12288 6000 12300
rect 5955 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 11308 12291 11366 12297
rect 11308 12257 11320 12291
rect 11354 12288 11366 12291
rect 11422 12288 11428 12300
rect 11354 12260 11428 12288
rect 11354 12257 11366 12260
rect 11308 12251 11366 12257
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6472 12192 7021 12220
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 1765 12155 1823 12161
rect 1765 12152 1777 12155
rect 1728 12124 1777 12152
rect 1728 12112 1734 12124
rect 1765 12121 1777 12124
rect 1811 12152 1823 12155
rect 3145 12155 3203 12161
rect 3145 12152 3157 12155
rect 1811 12124 3157 12152
rect 1811 12121 1823 12124
rect 1765 12115 1823 12121
rect 3145 12121 3157 12124
rect 3191 12152 3203 12155
rect 5626 12152 5632 12164
rect 3191 12124 5632 12152
rect 3191 12121 3203 12124
rect 3145 12115 3203 12121
rect 5626 12112 5632 12124
rect 5684 12112 5690 12164
rect 6472 12096 6500 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 7009 12183 7067 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 7926 12152 7932 12164
rect 7839 12124 7932 12152
rect 7926 12112 7932 12124
rect 7984 12152 7990 12164
rect 9858 12152 9864 12164
rect 7984 12124 9864 12152
rect 7984 12112 7990 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 2133 12087 2191 12093
rect 2133 12053 2145 12087
rect 2179 12084 2191 12087
rect 3050 12084 3056 12096
rect 2179 12056 3056 12084
rect 2179 12053 2191 12056
rect 2133 12047 2191 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4764 12056 4905 12084
rect 4764 12044 4770 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 6454 12084 6460 12096
rect 6415 12056 6460 12084
rect 4893 12047 4951 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 11379 12087 11437 12093
rect 11379 12084 11391 12087
rect 10652 12056 11391 12084
rect 10652 12044 10658 12056
rect 11379 12053 11391 12056
rect 11425 12053 11437 12087
rect 11379 12047 11437 12053
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2406 11880 2412 11892
rect 2367 11852 2412 11880
rect 2406 11840 2412 11852
rect 2464 11840 2470 11892
rect 3418 11880 3424 11892
rect 3379 11852 3424 11880
rect 3418 11840 3424 11852
rect 3476 11880 3482 11892
rect 4062 11880 4068 11892
rect 3476 11852 4068 11880
rect 3476 11840 3482 11852
rect 4062 11840 4068 11852
rect 4120 11880 4126 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4120 11852 4537 11880
rect 4120 11840 4126 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 4982 11880 4988 11892
rect 4943 11852 4988 11880
rect 4525 11843 4583 11849
rect 4982 11840 4988 11852
rect 5040 11880 5046 11892
rect 5994 11880 6000 11892
rect 5040 11852 6000 11880
rect 5040 11840 5046 11852
rect 2041 11815 2099 11821
rect 2041 11781 2053 11815
rect 2087 11812 2099 11815
rect 2087 11784 4154 11812
rect 2087 11781 2099 11784
rect 2041 11775 2099 11781
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2056 11676 2084 11775
rect 1443 11648 2084 11676
rect 3421 11679 3479 11685
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3436 11552 3464 11639
rect 4126 11608 4154 11784
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5132 11716 5304 11744
rect 5132 11704 5138 11716
rect 5276 11685 5304 11716
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11645 5319 11679
rect 5552 11676 5580 11852
rect 5994 11840 6000 11852
rect 6052 11880 6058 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 6052 11852 6193 11880
rect 6052 11840 6058 11852
rect 6181 11849 6193 11852
rect 6227 11849 6239 11883
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 6181 11843 6239 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6454 11744 6460 11756
rect 5951 11716 6460 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 8938 11744 8944 11756
rect 8711 11716 8944 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5552 11648 5641 11676
rect 5261 11639 5319 11645
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6236 11648 7021 11676
rect 6236 11636 6242 11648
rect 7009 11645 7021 11648
rect 7055 11676 7067 11679
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7055 11648 8217 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 6914 11608 6920 11620
rect 4126 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7330 11611 7388 11617
rect 7330 11608 7342 11611
rect 7024 11580 7342 11608
rect 7024 11552 7052 11580
rect 7330 11577 7342 11580
rect 7376 11577 7388 11611
rect 7330 11571 7388 11577
rect 8849 11611 8907 11617
rect 8849 11577 8861 11611
rect 8895 11577 8907 11611
rect 8849 11571 8907 11577
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 3016 11512 3065 11540
rect 3016 11500 3022 11512
rect 3053 11509 3065 11512
rect 3099 11540 3111 11543
rect 3418 11540 3424 11552
rect 3099 11512 3424 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 6641 11543 6699 11549
rect 4212 11512 4257 11540
rect 4212 11500 4218 11512
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 7006 11540 7012 11552
rect 6687 11512 7012 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7926 11540 7932 11552
rect 7887 11512 7932 11540
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 8864 11540 8892 11571
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9493 11611 9551 11617
rect 8996 11580 9041 11608
rect 8996 11568 9002 11580
rect 9493 11577 9505 11611
rect 9539 11608 9551 11611
rect 10226 11608 10232 11620
rect 9539 11580 10232 11608
rect 9539 11577 9551 11580
rect 9493 11571 9551 11577
rect 10226 11568 10232 11580
rect 10284 11608 10290 11620
rect 10413 11611 10471 11617
rect 10413 11608 10425 11611
rect 10284 11580 10425 11608
rect 10284 11568 10290 11580
rect 10413 11577 10425 11580
rect 10459 11577 10471 11611
rect 10413 11571 10471 11577
rect 10505 11611 10563 11617
rect 10505 11577 10517 11611
rect 10551 11577 10563 11611
rect 10505 11571 10563 11577
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 11514 11608 11520 11620
rect 11103 11580 11520 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 10134 11540 10140 11552
rect 8812 11512 8892 11540
rect 10095 11512 10140 11540
rect 8812 11500 8818 11512
rect 10134 11500 10140 11512
rect 10192 11540 10198 11552
rect 10520 11540 10548 11571
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 11422 11540 11428 11552
rect 10192 11512 10548 11540
rect 11335 11512 11428 11540
rect 10192 11500 10198 11512
rect 11422 11500 11428 11512
rect 11480 11540 11486 11552
rect 12618 11540 12624 11552
rect 11480 11512 12624 11540
rect 11480 11500 11486 11512
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 3510 11336 3516 11348
rect 1627 11308 3516 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5626 11336 5632 11348
rect 5587 11308 5632 11336
rect 5169 11299 5227 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 8205 11339 8263 11345
rect 8205 11305 8217 11339
rect 8251 11336 8263 11339
rect 8938 11336 8944 11348
rect 8251 11308 8944 11336
rect 8251 11305 8263 11308
rect 8205 11299 8263 11305
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9493 11339 9551 11345
rect 9493 11305 9505 11339
rect 9539 11336 9551 11339
rect 9766 11336 9772 11348
rect 9539 11308 9772 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 3142 11268 3148 11280
rect 2424 11240 2912 11268
rect 3103 11240 3148 11268
rect 2424 11212 2452 11240
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2406 11200 2412 11212
rect 2319 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2774 11200 2780 11212
rect 2731 11172 2780 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2700 11132 2728 11163
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 2884 11200 2912 11240
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 7606 11271 7664 11277
rect 7606 11268 7618 11271
rect 7064 11240 7618 11268
rect 7064 11228 7070 11240
rect 7606 11237 7618 11240
rect 7652 11237 7664 11271
rect 7606 11231 7664 11237
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 9858 11268 9864 11280
rect 7984 11240 9864 11268
rect 7984 11228 7990 11240
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 11422 11268 11428 11280
rect 11383 11240 11428 11268
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 4062 11200 4068 11212
rect 2884 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4338 11200 4344 11212
rect 4212 11172 4257 11200
rect 4299 11172 4344 11200
rect 4212 11160 4218 11172
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 5718 11200 5724 11212
rect 5679 11172 5724 11200
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 6052 11172 6193 11200
rect 6052 11160 6058 11172
rect 6181 11169 6193 11172
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 2363 11104 2728 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 3016 11104 4537 11132
rect 3016 11092 3022 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 7190 11132 7196 11144
rect 6503 11104 7196 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 9769 11135 9827 11141
rect 7340 11104 7385 11132
rect 7340 11092 7346 11104
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 9769 11095 9827 11101
rect 2498 11064 2504 11076
rect 2459 11036 2504 11064
rect 2498 11024 2504 11036
rect 2556 11024 2562 11076
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 7098 11064 7104 11076
rect 3108 11036 7104 11064
rect 3108 11024 3114 11036
rect 7098 11024 7104 11036
rect 7156 11064 7162 11076
rect 7650 11064 7656 11076
rect 7156 11036 7656 11064
rect 7156 11024 7162 11036
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 9784 11064 9812 11095
rect 10226 11092 10232 11104
rect 10284 11132 10290 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 10284 11104 10701 11132
rect 10284 11092 10290 11104
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 10594 11064 10600 11076
rect 9784 11036 10600 11064
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 3697 10999 3755 11005
rect 3697 10965 3709 10999
rect 3743 10996 3755 10999
rect 4246 10996 4252 11008
rect 3743 10968 4252 10996
rect 3743 10965 3755 10968
rect 3697 10959 3755 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 7006 10996 7012 11008
rect 6967 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 11348 10996 11376 11095
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11572 11104 11621 11132
rect 11572 11092 11578 11104
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 11606 10996 11612 11008
rect 9732 10968 11612 10996
rect 9732 10956 9738 10968
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 4982 10792 4988 10804
rect 4943 10764 4988 10792
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 6052 10764 6193 10792
rect 6052 10752 6058 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6181 10755 6239 10761
rect 7282 10752 7288 10804
rect 7340 10792 7346 10804
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 7340 10764 8585 10792
rect 7340 10752 7346 10764
rect 8573 10761 8585 10764
rect 8619 10761 8631 10795
rect 8573 10755 8631 10761
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8904 10764 8953 10792
rect 8904 10752 8910 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 9916 10764 10241 10792
rect 9916 10752 9922 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10594 10792 10600 10804
rect 10555 10764 10600 10792
rect 10229 10755 10287 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11606 10792 11612 10804
rect 11567 10764 11612 10792
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 3050 10684 3056 10736
rect 3108 10724 3114 10736
rect 3970 10724 3976 10736
rect 3108 10696 3976 10724
rect 3108 10684 3114 10696
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 8297 10727 8355 10733
rect 8297 10693 8309 10727
rect 8343 10724 8355 10727
rect 10134 10724 10140 10736
rect 8343 10696 10140 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 2498 10616 2504 10668
rect 2556 10656 2562 10668
rect 3145 10659 3203 10665
rect 3145 10656 3157 10659
rect 2556 10628 3157 10656
rect 2556 10616 2562 10628
rect 3145 10625 3157 10628
rect 3191 10656 3203 10659
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3191 10628 3709 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3697 10625 3709 10628
rect 3743 10656 3755 10659
rect 4246 10656 4252 10668
rect 3743 10628 4252 10656
rect 3743 10625 3755 10628
rect 3697 10619 3755 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 8260 10628 11253 10656
rect 8260 10616 8266 10628
rect 11241 10625 11253 10628
rect 11287 10656 11299 10659
rect 11422 10656 11428 10668
rect 11287 10628 11428 10656
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2682 10588 2688 10600
rect 1995 10560 2688 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 3528 10560 3617 10588
rect 2774 10520 2780 10532
rect 2735 10492 2780 10520
rect 2774 10480 2780 10492
rect 2832 10480 2838 10532
rect 3528 10464 3556 10560
rect 3605 10557 3617 10560
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 3881 10591 3939 10597
rect 3881 10557 3893 10591
rect 3927 10588 3939 10591
rect 3970 10588 3976 10600
rect 3927 10560 3976 10588
rect 3927 10557 3939 10560
rect 3881 10551 3939 10557
rect 3970 10548 3976 10560
rect 4028 10588 4034 10600
rect 4338 10588 4344 10600
rect 4028 10560 4344 10588
rect 4028 10548 4034 10560
rect 4338 10548 4344 10560
rect 4396 10588 4402 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4396 10560 4629 10588
rect 4396 10548 4402 10560
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 5534 10588 5540 10600
rect 5491 10560 5540 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 5994 10588 6000 10600
rect 5767 10560 6000 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 5994 10548 6000 10560
rect 6052 10548 6058 10600
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7156 10560 7389 10588
rect 7156 10548 7162 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 5902 10520 5908 10532
rect 5863 10492 5908 10520
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 7006 10520 7012 10532
rect 6687 10492 7012 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7006 10480 7012 10492
rect 7064 10520 7070 10532
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 7064 10492 7297 10520
rect 7064 10480 7070 10492
rect 7285 10489 7297 10492
rect 7331 10520 7343 10523
rect 7739 10523 7797 10529
rect 7739 10520 7751 10523
rect 7331 10492 7751 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7739 10489 7751 10492
rect 7785 10520 7797 10523
rect 8110 10520 8116 10532
rect 7785 10492 8116 10520
rect 7785 10489 7797 10492
rect 7739 10483 7797 10489
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 9214 10520 9220 10532
rect 9175 10492 9220 10520
rect 9214 10480 9220 10492
rect 9272 10480 9278 10532
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9324 10452 9352 10483
rect 9674 10480 9680 10532
rect 9732 10520 9738 10532
rect 9861 10523 9919 10529
rect 9861 10520 9873 10523
rect 9732 10492 9873 10520
rect 9732 10480 9738 10492
rect 9861 10489 9873 10492
rect 9907 10489 9919 10523
rect 9861 10483 9919 10489
rect 8904 10424 9352 10452
rect 8904 10412 8910 10424
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2406 10248 2412 10260
rect 2363 10220 2412 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2866 10248 2872 10260
rect 2827 10220 2872 10248
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5534 10248 5540 10260
rect 5307 10220 5540 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5718 10248 5724 10260
rect 5675 10220 5724 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 9214 10248 9220 10260
rect 9175 10220 9220 10248
rect 9214 10208 9220 10220
rect 9272 10248 9278 10260
rect 9815 10251 9873 10257
rect 9815 10248 9827 10251
rect 9272 10220 9827 10248
rect 9272 10208 9278 10220
rect 9815 10217 9827 10220
rect 9861 10217 9873 10251
rect 9815 10211 9873 10217
rect 1394 10140 1400 10192
rect 1452 10180 1458 10192
rect 1673 10183 1731 10189
rect 1673 10180 1685 10183
rect 1452 10152 1685 10180
rect 1452 10140 1458 10152
rect 1673 10149 1685 10152
rect 1719 10180 1731 10183
rect 4062 10180 4068 10192
rect 1719 10152 4068 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 6457 10183 6515 10189
rect 6457 10149 6469 10183
rect 6503 10180 6515 10183
rect 7098 10180 7104 10192
rect 6503 10152 7104 10180
rect 6503 10149 6515 10152
rect 6457 10143 6515 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7647 10183 7705 10189
rect 7647 10149 7659 10183
rect 7693 10180 7705 10183
rect 8110 10180 8116 10192
rect 7693 10152 8116 10180
rect 7693 10149 7705 10152
rect 7647 10143 7705 10149
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2556 10084 2601 10112
rect 2556 10072 2562 10084
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 4246 10112 4252 10124
rect 2740 10084 2833 10112
rect 4207 10084 4252 10112
rect 2740 10072 2746 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 5166 10112 5172 10124
rect 4488 10084 5172 10112
rect 4488 10072 4494 10084
rect 5166 10072 5172 10084
rect 5224 10112 5230 10124
rect 5721 10115 5779 10121
rect 5721 10112 5733 10115
rect 5224 10084 5733 10112
rect 5224 10072 5230 10084
rect 5721 10081 5733 10084
rect 5767 10081 5779 10115
rect 5721 10075 5779 10081
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6052 10084 6193 10112
rect 6052 10072 6058 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7248 10084 7297 10112
rect 7248 10072 7254 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 9744 10115 9802 10121
rect 9744 10081 9756 10115
rect 9790 10081 9802 10115
rect 9744 10075 9802 10081
rect 2700 10044 2728 10072
rect 3697 10047 3755 10053
rect 3697 10044 3709 10047
rect 2700 10016 3709 10044
rect 3697 10013 3709 10016
rect 3743 10044 3755 10047
rect 3970 10044 3976 10056
rect 3743 10016 3976 10044
rect 3743 10013 3755 10016
rect 3697 10007 3755 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4801 10047 4859 10053
rect 4801 10044 4813 10047
rect 4212 10016 4813 10044
rect 4212 10004 4218 10016
rect 4801 10013 4813 10016
rect 4847 10044 4859 10047
rect 5350 10044 5356 10056
rect 4847 10016 5356 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 9582 10044 9588 10056
rect 6972 10016 9588 10044
rect 6972 10004 6978 10016
rect 9582 10004 9588 10016
rect 9640 10044 9646 10056
rect 9759 10044 9787 10075
rect 9640 10016 9787 10044
rect 9640 10004 9646 10016
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 5442 9976 5448 9988
rect 3200 9948 5448 9976
rect 3200 9936 3206 9948
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 2133 9707 2191 9713
rect 2133 9673 2145 9707
rect 2179 9704 2191 9707
rect 2406 9704 2412 9716
rect 2179 9676 2412 9704
rect 2179 9673 2191 9676
rect 2133 9667 2191 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2777 9707 2835 9713
rect 2777 9704 2789 9707
rect 2556 9676 2789 9704
rect 2556 9664 2562 9676
rect 2777 9673 2789 9676
rect 2823 9673 2835 9707
rect 3142 9704 3148 9716
rect 3103 9676 3148 9704
rect 2777 9667 2835 9673
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3513 9707 3571 9713
rect 3513 9673 3525 9707
rect 3559 9704 3571 9707
rect 3970 9704 3976 9716
rect 3559 9676 3976 9704
rect 3559 9673 3571 9676
rect 3513 9667 3571 9673
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4985 9707 5043 9713
rect 4985 9704 4997 9707
rect 4304 9676 4997 9704
rect 4304 9664 4310 9676
rect 4985 9673 4997 9676
rect 5031 9673 5043 9707
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 4985 9667 5043 9673
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5994 9704 6000 9716
rect 5955 9676 6000 9704
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 8389 9707 8447 9713
rect 8389 9704 8401 9707
rect 7248 9676 8401 9704
rect 7248 9664 7254 9676
rect 8389 9673 8401 9676
rect 8435 9673 8447 9707
rect 8389 9667 8447 9673
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 8895 9707 8953 9713
rect 8895 9704 8907 9707
rect 8812 9676 8907 9704
rect 8812 9664 8818 9676
rect 8895 9673 8907 9676
rect 8941 9673 8953 9707
rect 9582 9704 9588 9716
rect 9543 9676 9588 9704
rect 8895 9667 8953 9673
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10318 9704 10324 9716
rect 10279 9676 10324 9704
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 11020 9676 11253 9704
rect 11020 9664 11026 9676
rect 11241 9673 11253 9676
rect 11287 9673 11299 9707
rect 11241 9667 11299 9673
rect 4062 9636 4068 9648
rect 4023 9608 4068 9636
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5721 9639 5779 9645
rect 5721 9605 5733 9639
rect 5767 9636 5779 9639
rect 8294 9636 8300 9648
rect 5767 9608 8300 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 7208 9580 7236 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2682 9568 2688 9580
rect 2547 9540 2688 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 4430 9568 4436 9580
rect 3292 9540 4436 9568
rect 3292 9528 3298 9540
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5316 9540 6561 9568
rect 5316 9528 5322 9540
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 6595 9540 7052 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 2958 9500 2964 9512
rect 2919 9472 2964 9500
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3804 9472 3985 9500
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3804 9373 3832 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4338 9500 4344 9512
rect 4295 9472 4344 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4338 9460 4344 9472
rect 4396 9460 4402 9512
rect 5534 9500 5540 9512
rect 5495 9472 5540 9500
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 7024 9509 7052 9540
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7009 9463 7067 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8824 9503 8882 9509
rect 8824 9469 8836 9503
rect 8870 9500 8882 9503
rect 9836 9503 9894 9509
rect 8870 9472 9352 9500
rect 8870 9469 8882 9472
rect 8824 9463 8882 9469
rect 7742 9432 7748 9444
rect 7703 9404 7748 9432
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 9324 9441 9352 9472
rect 9836 9469 9848 9503
rect 9882 9500 9894 9503
rect 10318 9500 10324 9512
rect 9882 9472 10324 9500
rect 9882 9469 9894 9472
rect 9836 9463 9894 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10848 9503 10906 9509
rect 10848 9469 10860 9503
rect 10894 9500 10906 9503
rect 10962 9500 10968 9512
rect 10894 9472 10968 9500
rect 10894 9469 10906 9472
rect 10848 9463 10906 9469
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9490 9432 9496 9444
rect 9355 9404 9496 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9490 9392 9496 9404
rect 9548 9432 9554 9444
rect 10686 9432 10692 9444
rect 9548 9404 10692 9432
rect 9548 9392 9554 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3568 9336 3801 9364
rect 3568 9324 3574 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 3789 9327 3847 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 9907 9367 9965 9373
rect 9907 9364 9919 9367
rect 9732 9336 9919 9364
rect 9732 9324 9738 9336
rect 9907 9333 9919 9336
rect 9953 9333 9965 9367
rect 9907 9327 9965 9333
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10919 9367 10977 9373
rect 10919 9364 10931 9367
rect 10560 9336 10931 9364
rect 10560 9324 10566 9336
rect 10919 9333 10931 9336
rect 10965 9333 10977 9367
rect 10919 9327 10977 9333
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2958 9160 2964 9172
rect 2919 9132 2964 9160
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 5166 9160 5172 9172
rect 5127 9132 5172 9160
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9640 9132 10456 9160
rect 9640 9120 9646 9132
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 4798 9092 4804 9104
rect 2832 9064 4384 9092
rect 4759 9064 4804 9092
rect 2832 9052 2838 9064
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3568 8996 4077 9024
rect 3568 8984 3574 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4246 9024 4252 9036
rect 4203 8996 4252 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4172 8888 4200 8987
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4356 9033 4384 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 6638 9092 6644 9104
rect 6135 9064 6644 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 9861 9095 9919 9101
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 10226 9092 10232 9104
rect 9907 9064 10232 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 10226 9052 10232 9064
rect 10284 9052 10290 9104
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 4982 9024 4988 9036
rect 4387 8996 4988 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 10428 9024 10456 9132
rect 11238 9024 11244 9036
rect 11296 9033 11302 9036
rect 11296 9027 11334 9033
rect 10428 8996 11244 9024
rect 7929 8987 7987 8993
rect 5994 8956 6000 8968
rect 5955 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 6730 8956 6736 8968
rect 6687 8928 6736 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7484 8888 7512 8987
rect 7834 8888 7840 8900
rect 4028 8860 4200 8888
rect 5092 8860 7840 8888
rect 4028 8848 4034 8860
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 5092 8820 5120 8860
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 7098 8820 7104 8832
rect 3384 8792 5120 8820
rect 7059 8792 7104 8820
rect 3384 8780 3390 8792
rect 7098 8780 7104 8792
rect 7156 8820 7162 8832
rect 7558 8820 7564 8832
rect 7156 8792 7564 8820
rect 7156 8780 7162 8792
rect 7558 8780 7564 8792
rect 7616 8820 7622 8832
rect 7944 8820 7972 8987
rect 11238 8984 11244 8996
rect 11322 9024 11334 9027
rect 11422 9024 11428 9036
rect 11322 8996 11428 9024
rect 11322 8993 11334 8996
rect 11296 8987 11334 8993
rect 11296 8984 11302 8987
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 9815 8928 10640 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 10410 8888 10416 8900
rect 10367 8860 10416 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 10612 8832 10640 8928
rect 7616 8792 7972 8820
rect 7616 8780 7622 8792
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 11379 8823 11437 8829
rect 11379 8820 11391 8823
rect 10652 8792 11391 8820
rect 10652 8780 10658 8792
rect 11379 8789 11391 8792
rect 11425 8789 11437 8823
rect 11379 8783 11437 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3510 8616 3516 8628
rect 2924 8588 3516 8616
rect 2924 8576 2930 8588
rect 3510 8576 3516 8588
rect 3568 8616 3574 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 3568 8588 4629 8616
rect 3568 8576 3574 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4982 8616 4988 8628
rect 4943 8588 4988 8616
rect 4617 8579 4675 8585
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 7834 8616 7840 8628
rect 7795 8588 7840 8616
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11480 8588 11529 8616
rect 11480 8576 11486 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 2041 8551 2099 8557
rect 2041 8548 2053 8551
rect 1811 8520 2053 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 2041 8517 2053 8520
rect 2087 8548 2099 8551
rect 3050 8548 3056 8560
rect 2087 8520 3056 8548
rect 2087 8517 2099 8520
rect 2041 8511 2099 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 4341 8551 4399 8557
rect 4341 8548 4353 8551
rect 4120 8520 4353 8548
rect 4120 8508 4126 8520
rect 4341 8517 4353 8520
rect 4387 8517 4399 8551
rect 5810 8548 5816 8560
rect 5723 8520 5816 8548
rect 4341 8511 4399 8517
rect 5810 8508 5816 8520
rect 5868 8548 5874 8560
rect 7469 8551 7527 8557
rect 7469 8548 7481 8551
rect 5868 8520 7481 8548
rect 5868 8508 5874 8520
rect 7469 8517 7481 8520
rect 7515 8517 7527 8551
rect 7469 8511 7527 8517
rect 106 8440 112 8492
rect 164 8480 170 8492
rect 164 8452 2452 8480
rect 164 8440 170 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 1443 8384 1777 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1765 8381 1777 8384
rect 1811 8381 1823 8415
rect 2424 8412 2452 8452
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 3384 8452 6929 8480
rect 3384 8440 3390 8452
rect 6917 8449 6929 8452
rect 6963 8480 6975 8483
rect 7282 8480 7288 8492
rect 6963 8452 7288 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 9214 8480 9220 8492
rect 9127 8452 9220 8480
rect 9214 8440 9220 8452
rect 9272 8480 9278 8492
rect 9674 8480 9680 8492
rect 9272 8452 9680 8480
rect 9272 8440 9278 8452
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 3180 8415 3238 8421
rect 3180 8412 3192 8415
rect 2424 8384 3192 8412
rect 1765 8375 1823 8381
rect 3180 8381 3192 8384
rect 3226 8412 3238 8415
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3226 8384 3617 8412
rect 3226 8381 3238 8384
rect 3180 8375 3238 8381
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4614 8412 4620 8424
rect 4203 8384 4620 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 10778 8421 10784 8424
rect 10756 8415 10784 8421
rect 10756 8412 10768 8415
rect 10691 8384 10768 8412
rect 10756 8381 10768 8384
rect 10836 8412 10842 8424
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 10836 8384 11161 8412
rect 10756 8375 10784 8381
rect 10778 8372 10784 8375
rect 10836 8372 10842 8384
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 3283 8347 3341 8353
rect 3283 8313 3295 8347
rect 3329 8344 3341 8347
rect 3786 8344 3792 8356
rect 3329 8316 3792 8344
rect 3329 8313 3341 8316
rect 3283 8307 3341 8313
rect 3786 8304 3792 8316
rect 3844 8344 3850 8356
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 3844 8316 5273 8344
rect 3844 8304 3850 8316
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8313 5411 8347
rect 5353 8307 5411 8313
rect 7009 8347 7067 8353
rect 7009 8313 7021 8347
rect 7055 8313 7067 8347
rect 9030 8344 9036 8356
rect 8943 8316 9036 8344
rect 7009 8307 7067 8313
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 5368 8276 5396 8307
rect 6178 8276 6184 8288
rect 5368 8248 6184 8276
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 6638 8236 6644 8248
rect 6696 8276 6702 8288
rect 7024 8276 7052 8307
rect 9030 8304 9036 8316
rect 9088 8344 9094 8356
rect 9286 8347 9344 8353
rect 9286 8344 9298 8347
rect 9088 8316 9298 8344
rect 9088 8304 9094 8316
rect 9286 8313 9298 8316
rect 9332 8313 9344 8347
rect 9858 8344 9864 8356
rect 9819 8316 9864 8344
rect 9286 8307 9344 8313
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 6696 8248 7052 8276
rect 6696 8236 6702 8248
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7466 8276 7472 8288
rect 7156 8248 7472 8276
rect 7156 8236 7162 8248
rect 7466 8236 7472 8248
rect 7524 8276 7530 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7524 8248 8217 8276
rect 7524 8236 7530 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 10226 8276 10232 8288
rect 10187 8248 10232 8276
rect 8205 8239 8263 8245
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 10827 8279 10885 8285
rect 10827 8276 10839 8279
rect 10652 8248 10839 8276
rect 10652 8236 10658 8248
rect 10827 8245 10839 8248
rect 10873 8245 10885 8279
rect 10827 8239 10885 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 3099 8075 3157 8081
rect 3099 8041 3111 8075
rect 3145 8072 3157 8075
rect 3326 8072 3332 8084
rect 3145 8044 3332 8072
rect 3145 8041 3157 8044
rect 3099 8035 3157 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4203 8075 4261 8081
rect 4203 8041 4215 8075
rect 4249 8072 4261 8075
rect 5994 8072 6000 8084
rect 4249 8044 6000 8072
rect 4249 8041 4261 8044
rect 4203 8035 4261 8041
rect 5994 8032 6000 8044
rect 6052 8072 6058 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6052 8044 6653 8072
rect 6052 8032 6058 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 7282 8072 7288 8084
rect 7243 8044 7288 8072
rect 6641 8035 6699 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 8110 8032 8116 8084
rect 8168 8072 8174 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 8168 8044 8217 8072
rect 8168 8032 8174 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 8205 8035 8263 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 4614 8004 4620 8016
rect 4575 7976 4620 8004
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 5330 8007 5388 8013
rect 5330 7973 5342 8007
rect 5376 8004 5388 8007
rect 5442 8004 5448 8016
rect 5376 7976 5448 8004
rect 5376 7973 5388 7976
rect 5330 7967 5388 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 9582 8004 9588 8016
rect 9088 7976 9588 8004
rect 9088 7964 9094 7976
rect 9582 7964 9588 7976
rect 9640 8004 9646 8016
rect 9861 8007 9919 8013
rect 9861 8004 9873 8007
rect 9640 7976 9873 8004
rect 9640 7964 9646 7976
rect 9861 7973 9873 7976
rect 9907 7973 9919 8007
rect 10410 8004 10416 8016
rect 10371 7976 10416 8004
rect 9861 7967 9919 7973
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2958 7936 2964 7948
rect 3016 7945 3022 7948
rect 3016 7939 3054 7945
rect 2188 7908 2964 7936
rect 2188 7896 2194 7908
rect 2958 7896 2964 7908
rect 3042 7905 3054 7939
rect 3016 7899 3054 7905
rect 4132 7939 4190 7945
rect 4132 7905 4144 7939
rect 4178 7936 4190 7939
rect 4430 7936 4436 7948
rect 4178 7908 4436 7936
rect 4178 7905 4190 7908
rect 4132 7899 4190 7905
rect 3016 7896 3022 7899
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 6822 7936 6828 7948
rect 6783 7908 6828 7936
rect 6822 7896 6828 7908
rect 6880 7896 6886 7948
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7800 7908 7849 7936
rect 7800 7896 7806 7908
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 11308 7939 11366 7945
rect 11308 7905 11320 7939
rect 11354 7936 11366 7939
rect 11514 7936 11520 7948
rect 11354 7908 11520 7936
rect 11354 7905 11366 7908
rect 11308 7899 11366 7905
rect 11514 7896 11520 7908
rect 11572 7936 11578 7948
rect 12066 7936 12072 7948
rect 11572 7908 12072 7936
rect 11572 7896 11578 7908
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5166 7868 5172 7880
rect 5123 7840 5172 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9548 7840 9781 7868
rect 9548 7828 9554 7840
rect 9769 7837 9781 7840
rect 9815 7868 9827 7871
rect 10502 7868 10508 7880
rect 9815 7840 10508 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7800 8815 7803
rect 10226 7800 10232 7812
rect 8803 7772 10232 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7732 3571 7735
rect 4062 7732 4068 7744
rect 3559 7704 4068 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4982 7732 4988 7744
rect 4943 7704 4988 7732
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6178 7732 6184 7744
rect 6043 7704 6184 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6546 7732 6552 7744
rect 6328 7704 6552 7732
rect 6328 7692 6334 7704
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7009 7735 7067 7741
rect 7009 7701 7021 7735
rect 7055 7732 7067 7735
rect 7466 7732 7472 7744
rect 7055 7704 7472 7732
rect 7055 7701 7067 7704
rect 7009 7695 7067 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 11379 7735 11437 7741
rect 11379 7732 11391 7735
rect 10744 7704 11391 7732
rect 10744 7692 10750 7704
rect 11379 7701 11391 7704
rect 11425 7701 11437 7735
rect 11379 7695 11437 7701
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 2958 7528 2964 7540
rect 2919 7500 2964 7528
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4430 7528 4436 7540
rect 4391 7500 4436 7528
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6270 7528 6276 7540
rect 5951 7500 6276 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 9640 7500 9689 7528
rect 9640 7488 9646 7500
rect 9677 7497 9689 7500
rect 9723 7528 9735 7531
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9723 7500 9965 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 11514 7528 11520 7540
rect 11475 7500 11520 7528
rect 9953 7491 10011 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 2590 7420 2596 7472
rect 2648 7460 2654 7472
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 2648 7432 6193 7460
rect 2648 7420 2654 7432
rect 6181 7429 6193 7432
rect 6227 7460 6239 7463
rect 6822 7460 6828 7472
rect 6227 7432 6828 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 9916 7432 10916 7460
rect 9916 7420 9922 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4982 7392 4988 7404
rect 4203 7364 4988 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5902 7352 5908 7404
rect 5960 7392 5966 7404
rect 7006 7392 7012 7404
rect 5960 7364 7012 7392
rect 5960 7352 5966 7364
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8260 7364 8769 7392
rect 8260 7352 8266 7364
rect 8757 7361 8769 7364
rect 8803 7392 8815 7395
rect 9030 7392 9036 7404
rect 8803 7364 9036 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 10888 7401 10916 7432
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4062 7324 4068 7336
rect 4019 7296 4068 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 4890 7324 4896 7336
rect 4120 7296 4896 7324
rect 4120 7284 4126 7296
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 8662 7324 8668 7336
rect 5000 7296 8668 7324
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 5000 7256 5028 7296
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 3016 7228 5028 7256
rect 5306 7259 5364 7265
rect 3016 7216 3022 7228
rect 5306 7225 5318 7259
rect 5352 7225 5364 7259
rect 5306 7219 5364 7225
rect 7371 7259 7429 7265
rect 7371 7225 7383 7259
rect 7417 7256 7429 7259
rect 9078 7259 9136 7265
rect 7417 7228 8156 7256
rect 7417 7225 7429 7228
rect 7371 7219 7429 7225
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 5321 7188 5349 7219
rect 8128 7200 8156 7228
rect 9078 7225 9090 7259
rect 9124 7225 9136 7259
rect 9078 7219 9136 7225
rect 5442 7188 5448 7200
rect 4939 7160 5448 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 5442 7148 5448 7160
rect 5500 7188 5506 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 5500 7160 6561 7188
rect 5500 7148 5506 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 7926 7188 7932 7200
rect 7887 7160 7932 7188
rect 6549 7151 6607 7157
rect 7926 7148 7932 7160
rect 7984 7148 7990 7200
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 8168 7160 8217 7188
rect 8168 7148 8174 7160
rect 8205 7157 8217 7160
rect 8251 7188 8263 7191
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8251 7160 8585 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 8573 7157 8585 7160
rect 8619 7188 8631 7191
rect 9093 7188 9121 7219
rect 10226 7216 10232 7268
rect 10284 7256 10290 7268
rect 10413 7259 10471 7265
rect 10413 7256 10425 7259
rect 10284 7228 10425 7256
rect 10284 7216 10290 7228
rect 10413 7225 10425 7228
rect 10459 7256 10471 7259
rect 10689 7259 10747 7265
rect 10689 7256 10701 7259
rect 10459 7228 10701 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 10689 7225 10701 7228
rect 10735 7225 10747 7259
rect 10689 7219 10747 7225
rect 8619 7160 9121 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 3418 6984 3424 6996
rect 3379 6956 3424 6984
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 5258 6984 5264 6996
rect 4724 6956 5264 6984
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4724 6857 4752 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7006 6984 7012 6996
rect 6967 6956 7012 6984
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 8168 6956 8217 6984
rect 8168 6944 8174 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 8205 6947 8263 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 10652 6956 10701 6984
rect 10652 6944 10658 6956
rect 10689 6953 10701 6956
rect 10735 6953 10747 6987
rect 10689 6947 10747 6953
rect 5166 6916 5172 6928
rect 5127 6888 5172 6916
rect 5166 6876 5172 6888
rect 5224 6916 5230 6928
rect 5813 6919 5871 6925
rect 5813 6916 5825 6919
rect 5224 6888 5825 6916
rect 5224 6876 5230 6888
rect 5813 6885 5825 6888
rect 5859 6885 5871 6919
rect 6178 6916 6184 6928
rect 6139 6888 6184 6916
rect 5813 6879 5871 6885
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 6730 6916 6736 6928
rect 6691 6888 6736 6916
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 9306 6876 9312 6928
rect 9364 6916 9370 6928
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 9364 6888 9873 6916
rect 9364 6876 9370 6888
rect 9861 6885 9873 6888
rect 9907 6885 9919 6919
rect 10410 6916 10416 6928
rect 10371 6888 10416 6916
rect 9861 6879 9919 6885
rect 10410 6876 10416 6888
rect 10468 6876 10474 6928
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4120 6820 4721 6848
rect 4120 6808 4126 6820
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 4890 6848 4896 6860
rect 4851 6820 4896 6848
rect 4709 6811 4767 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 12320 6851 12378 6857
rect 12320 6817 12332 6851
rect 12366 6848 12378 6851
rect 12618 6848 12624 6860
rect 12366 6820 12624 6848
rect 12366 6817 12378 6820
rect 12320 6811 12378 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 6086 6780 6092 6792
rect 6047 6752 6092 6780
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 10686 6780 10692 6792
rect 9815 6752 10692 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 11238 6780 11244 6792
rect 11199 6752 11244 6780
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 7742 6712 7748 6724
rect 3108 6684 7748 6712
rect 3108 6672 3114 6684
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 5442 6644 5448 6656
rect 5403 6616 5448 6644
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 12391 6647 12449 6653
rect 12391 6644 12403 6647
rect 9548 6616 12403 6644
rect 9548 6604 9554 6616
rect 12391 6613 12403 6616
rect 12437 6613 12449 6647
rect 12391 6607 12449 6613
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 1854 6400 1860 6452
rect 1912 6440 1918 6452
rect 5721 6443 5779 6449
rect 1912 6412 4476 6440
rect 1912 6400 1918 6412
rect 4062 6372 4068 6384
rect 4023 6344 4068 6372
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 4448 6245 4476 6412
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 6086 6440 6092 6452
rect 5767 6412 6092 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8294 6440 8300 6452
rect 7708 6412 8300 6440
rect 7708 6400 7714 6412
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8812 6412 8953 6440
rect 8812 6400 8818 6412
rect 8941 6409 8953 6412
rect 8987 6440 8999 6443
rect 9306 6440 9312 6452
rect 8987 6412 9312 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9306 6400 9312 6412
rect 9364 6440 9370 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 9364 6412 10149 6440
rect 9364 6400 9370 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6440 11023 6443
rect 11241 6443 11299 6449
rect 11241 6440 11253 6443
rect 11011 6412 11253 6440
rect 11011 6409 11023 6412
rect 10965 6403 11023 6409
rect 11241 6409 11253 6412
rect 11287 6440 11299 6443
rect 11422 6440 11428 6452
rect 11287 6412 11428 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6178 6372 6184 6384
rect 6043 6344 6184 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6178 6332 6184 6344
rect 6236 6332 6242 6384
rect 10827 6375 10885 6381
rect 10827 6341 10839 6375
rect 10873 6372 10885 6375
rect 15102 6372 15108 6384
rect 10873 6344 15108 6372
rect 10873 6341 10885 6344
rect 10827 6335 10885 6341
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 7653 6307 7711 6313
rect 4816 6276 6684 6304
rect 4816 6245 4844 6276
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4479 6208 4813 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4801 6205 4813 6208
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 4890 6196 4896 6248
rect 4948 6236 4954 6248
rect 6656 6245 6684 6276
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7834 6304 7840 6316
rect 7699 6276 7840 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 7834 6264 7840 6276
rect 7892 6304 7898 6316
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7892 6276 8309 6304
rect 7892 6264 7898 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 9217 6307 9275 6313
rect 9217 6273 9229 6307
rect 9263 6304 9275 6307
rect 9490 6304 9496 6316
rect 9263 6276 9496 6304
rect 9263 6273 9275 6276
rect 9217 6267 9275 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4948 6208 4997 6236
rect 4948 6196 4954 6208
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6687 6208 6929 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 7466 6236 7472 6248
rect 7427 6208 7472 6236
rect 6917 6199 6975 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10756 6239 10814 6245
rect 10756 6236 10768 6239
rect 10560 6208 10768 6236
rect 10560 6196 10566 6208
rect 10756 6205 10768 6208
rect 10802 6236 10814 6239
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10802 6208 10977 6236
rect 10802 6205 10814 6208
rect 10756 6199 10814 6205
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 106 6128 112 6180
rect 164 6168 170 6180
rect 2038 6168 2044 6180
rect 164 6140 2044 6168
rect 164 6128 170 6140
rect 2038 6128 2044 6140
rect 2096 6168 2102 6180
rect 7006 6168 7012 6180
rect 2096 6140 7012 6168
rect 2096 6128 2102 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 9858 6168 9864 6180
rect 9364 6140 9409 6168
rect 9819 6140 9864 6168
rect 9364 6128 9370 6140
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8110 6100 8116 6112
rect 8067 6072 8116 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 12618 6100 12624 6112
rect 12579 6072 12624 6100
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4890 5896 4896 5908
rect 4571 5868 4896 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 5767 5899 5825 5905
rect 5767 5865 5779 5899
rect 5813 5896 5825 5899
rect 6086 5896 6092 5908
rect 5813 5868 6092 5896
rect 5813 5865 5825 5868
rect 5767 5859 5825 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 9490 5896 9496 5908
rect 9263 5868 9496 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 7009 5831 7067 5837
rect 7009 5797 7021 5831
rect 7055 5828 7067 5831
rect 7055 5800 7512 5828
rect 7055 5797 7067 5800
rect 7009 5791 7067 5797
rect 7484 5772 7512 5800
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 7984 5800 9873 5828
rect 7984 5788 7990 5800
rect 9861 5797 9873 5800
rect 9907 5828 9919 5831
rect 10042 5828 10048 5840
rect 9907 5800 10048 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10413 5831 10471 5837
rect 10413 5797 10425 5831
rect 10459 5828 10471 5831
rect 10502 5828 10508 5840
rect 10459 5800 10508 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 10502 5788 10508 5800
rect 10560 5788 10566 5840
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 5626 5760 5632 5772
rect 5583 5732 5632 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7248 5732 7297 5760
rect 7248 5720 7254 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7524 5732 7849 5760
rect 7524 5720 7530 5732
rect 7837 5729 7849 5732
rect 7883 5760 7895 5763
rect 8478 5760 8484 5772
rect 7883 5732 8484 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 9766 5692 9772 5704
rect 9679 5664 9772 5692
rect 9766 5652 9772 5664
rect 9824 5692 9830 5704
rect 11238 5692 11244 5704
rect 9824 5664 11244 5692
rect 9824 5652 9830 5664
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5684 5324 6193 5352
rect 5684 5312 5690 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 6503 5324 8125 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 8113 5321 8125 5324
rect 8159 5352 8171 5355
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 8159 5324 8217 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 8205 5315 8263 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10042 5352 10048 5364
rect 10003 5324 10048 5352
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 4632 5216 4660 5312
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 5960 5256 7052 5284
rect 5960 5244 5966 5256
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4632 5188 4997 5216
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6788 5188 6929 5216
rect 6788 5176 6794 5188
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 7024 5216 7052 5256
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7024 5188 7205 5216
rect 6917 5179 6975 5185
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 7975 5188 8524 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8496 5160 8524 5188
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 4764 5120 6469 5148
rect 4764 5108 4770 5120
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8159 5120 8401 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 8536 5120 8953 5148
rect 8536 5108 8542 5120
rect 8941 5117 8953 5120
rect 8987 5148 8999 5151
rect 10226 5148 10232 5160
rect 8987 5120 10232 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 5306 5083 5364 5089
rect 5306 5080 5318 5083
rect 4816 5052 5318 5080
rect 4816 5024 4844 5052
rect 5306 5049 5318 5052
rect 5352 5080 5364 5083
rect 5442 5080 5448 5092
rect 5352 5052 5448 5080
rect 5352 5049 5364 5052
rect 5306 5043 5364 5049
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5049 7067 5083
rect 7009 5043 7067 5049
rect 4798 5012 4804 5024
rect 4759 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6086 5012 6092 5024
rect 5951 4984 6092 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6822 5012 6828 5024
rect 6687 4984 6828 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6822 4972 6828 4984
rect 6880 5012 6886 5024
rect 7024 5012 7052 5043
rect 8478 5012 8484 5024
rect 6880 4984 7052 5012
rect 8439 4984 8484 5012
rect 6880 4972 6886 4984
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 5408 4780 5457 4808
rect 5408 4768 5414 4780
rect 5445 4777 5457 4780
rect 5491 4808 5503 4811
rect 5810 4808 5816 4820
rect 5491 4780 5816 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 6730 4808 6736 4820
rect 6656 4780 6736 4808
rect 6086 4740 6092 4752
rect 6047 4712 6092 4740
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 6656 4749 6684 4780
rect 6730 4768 6736 4780
rect 6788 4808 6794 4820
rect 6917 4811 6975 4817
rect 6917 4808 6929 4811
rect 6788 4780 6929 4808
rect 6788 4768 6794 4780
rect 6917 4777 6929 4780
rect 6963 4777 6975 4811
rect 6917 4771 6975 4777
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7248 4780 7297 4808
rect 7248 4768 7254 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8260 4780 8585 4808
rect 8260 4768 8266 4780
rect 8573 4777 8585 4780
rect 8619 4808 8631 4811
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 8619 4780 9781 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10468 4780 10701 4808
rect 10468 4768 10474 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 6641 4743 6699 4749
rect 6641 4709 6653 4743
rect 6687 4709 6699 4743
rect 7650 4740 7656 4752
rect 7611 4712 7656 4740
rect 6641 4703 6699 4709
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4706 4672 4712 4684
rect 4663 4644 4712 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 9674 4672 9680 4684
rect 9635 4644 9680 4672
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 10226 4672 10232 4684
rect 10139 4644 10232 4672
rect 10226 4632 10232 4644
rect 10284 4672 10290 4684
rect 10962 4672 10968 4684
rect 10284 4644 10968 4672
rect 10284 4632 10290 4644
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 4724 4536 4752 4632
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5994 4604 6000 4616
rect 5955 4576 6000 4604
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7340 4576 7573 4604
rect 7340 4564 7346 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 4982 4536 4988 4548
rect 4724 4508 4988 4536
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 7852 4536 7880 4567
rect 5868 4508 7880 4536
rect 5868 4496 5874 4508
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 8386 4468 8392 4480
rect 4212 4440 8392 4468
rect 4212 4428 4218 4440
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 3418 4264 3424 4276
rect 3160 4236 3424 4264
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4128 3111 4131
rect 3160 4128 3188 4236
rect 3418 4224 3424 4236
rect 3476 4264 3482 4276
rect 3697 4267 3755 4273
rect 3697 4264 3709 4267
rect 3476 4236 3709 4264
rect 3476 4224 3482 4236
rect 3697 4233 3709 4236
rect 3743 4264 3755 4267
rect 4154 4264 4160 4276
rect 3743 4236 4160 4264
rect 3743 4233 3755 4236
rect 3697 4227 3755 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4295 4267 4353 4273
rect 4295 4233 4307 4267
rect 4341 4264 4353 4267
rect 5994 4264 6000 4276
rect 4341 4236 6000 4264
rect 4341 4233 4353 4236
rect 4295 4227 4353 4233
rect 5994 4224 6000 4236
rect 6052 4264 6058 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6052 4236 6561 4264
rect 6052 4224 6058 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 9674 4264 9680 4276
rect 8352 4236 9680 4264
rect 8352 4224 8358 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10410 4264 10416 4276
rect 10060 4236 10416 4264
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 4890 4196 4896 4208
rect 4111 4168 4896 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 4982 4156 4988 4208
rect 5040 4196 5046 4208
rect 5040 4168 5085 4196
rect 5040 4156 5046 4168
rect 6086 4156 6092 4208
rect 6144 4196 6150 4208
rect 6181 4199 6239 4205
rect 6181 4196 6193 4199
rect 6144 4168 6193 4196
rect 6144 4156 6150 4168
rect 6181 4165 6193 4168
rect 6227 4196 6239 4199
rect 7469 4199 7527 4205
rect 7469 4196 7481 4199
rect 6227 4168 7481 4196
rect 6227 4165 6239 4168
rect 6181 4159 6239 4165
rect 7469 4165 7481 4168
rect 7515 4196 7527 4199
rect 7650 4196 7656 4208
rect 7515 4168 7656 4196
rect 7515 4165 7527 4168
rect 7469 4159 7527 4165
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 3099 4100 3188 4128
rect 3283 4131 3341 4137
rect 3099 4097 3111 4100
rect 3053 4091 3111 4097
rect 3283 4097 3295 4131
rect 3329 4128 3341 4131
rect 7282 4128 7288 4140
rect 3329 4100 7288 4128
rect 3329 4097 3341 4100
rect 3283 4091 3341 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 10060 4137 10088 4236
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 10962 4264 10968 4276
rect 10923 4236 10968 4264
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10023 4100 10057 4128
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10318 4128 10324 4140
rect 10279 4100 10324 4128
rect 10045 4091 10103 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 4224 4063 4282 4069
rect 4224 4029 4236 4063
rect 4270 4060 4282 4063
rect 4270 4032 4752 4060
rect 4270 4029 4282 4032
rect 4224 4023 4282 4029
rect 4724 3933 4752 4032
rect 5258 3992 5264 4004
rect 5219 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 5353 3995 5411 4001
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5442 3992 5448 4004
rect 5399 3964 5448 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5902 3992 5908 4004
rect 5863 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7374 3992 7380 4004
rect 6288 3964 7380 3992
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 6288 3924 6316 3964
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 8526 3995 8584 4001
rect 8526 3961 8538 3995
rect 8572 3961 8584 3995
rect 10134 3992 10140 4004
rect 10095 3964 10140 3992
rect 8526 3955 8584 3961
rect 4755 3896 6316 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6696 3896 6837 3924
rect 6696 3884 6702 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 6825 3887 6883 3893
rect 8110 3884 8116 3896
rect 8168 3924 8174 3936
rect 8541 3924 8569 3955
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 9122 3924 9128 3936
rect 8168 3896 8569 3924
rect 9083 3896 9128 3924
rect 8168 3884 8174 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 5132 3692 5733 3720
rect 5132 3680 5138 3692
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 6273 3723 6331 3729
rect 6273 3720 6285 3723
rect 6236 3692 6285 3720
rect 6236 3680 6242 3692
rect 6273 3689 6285 3692
rect 6319 3689 6331 3723
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6273 3683 6331 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8478 3720 8484 3732
rect 7791 3692 8484 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3553 4675 3587
rect 4890 3584 4896 3596
rect 4851 3556 4896 3584
rect 4617 3547 4675 3553
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4632 3516 4660 3547
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 7852 3593 7880 3692
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8757 3723 8815 3729
rect 8757 3689 8769 3723
rect 8803 3720 8815 3723
rect 10134 3720 10140 3732
rect 8803 3692 10140 3720
rect 8803 3689 8815 3692
rect 8757 3683 8815 3689
rect 10134 3680 10140 3692
rect 10192 3720 10198 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10192 3692 10701 3720
rect 10192 3680 10198 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 8110 3652 8116 3664
rect 8071 3624 8116 3652
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 9122 3612 9128 3664
rect 9180 3652 9186 3664
rect 9490 3652 9496 3664
rect 9180 3624 9496 3652
rect 9180 3612 9186 3624
rect 9490 3612 9496 3624
rect 9548 3652 9554 3664
rect 9861 3655 9919 3661
rect 9861 3652 9873 3655
rect 9548 3624 9873 3652
rect 9548 3612 9554 3624
rect 9861 3621 9873 3624
rect 9907 3621 9919 3655
rect 9861 3615 9919 3621
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 5077 3519 5135 3525
rect 4580 3488 5028 3516
rect 4580 3476 4586 3488
rect 5000 3448 5028 3488
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5123 3488 5917 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5905 3485 5917 3488
rect 5951 3516 5963 3519
rect 6546 3516 6552 3528
rect 5951 3488 6552 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8076 3488 9045 3516
rect 8076 3476 8082 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9033 3479 9091 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 10100 3488 11253 3516
rect 10100 3476 10106 3488
rect 11241 3485 11253 3488
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 8294 3448 8300 3460
rect 5000 3420 8300 3448
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 10318 3448 10324 3460
rect 10279 3420 10324 3448
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 5442 3380 5448 3392
rect 5403 3352 5448 3380
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 12618 3380 12624 3392
rect 5592 3352 12624 3380
rect 5592 3340 5598 3352
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 106 3136 112 3188
rect 164 3176 170 3188
rect 3970 3176 3976 3188
rect 164 3148 3976 3176
rect 164 3136 170 3148
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4522 3176 4528 3188
rect 4483 3148 4528 3176
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5500 3148 5917 3176
rect 5500 3136 5506 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 5905 3139 5963 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 9490 3176 9496 3188
rect 9451 3148 9496 3176
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 9824 3148 11345 3176
rect 9824 3136 9830 3148
rect 11333 3145 11345 3148
rect 11379 3145 11391 3179
rect 11333 3139 11391 3145
rect 3804 3080 5304 3108
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3375 2944 3709 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3697 2941 3709 2944
rect 3743 2972 3755 2975
rect 3804 2972 3832 3080
rect 4890 3040 4896 3052
rect 3988 3012 4896 3040
rect 3988 2984 4016 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5074 3040 5080 3052
rect 5031 3012 5080 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5276 3040 5304 3080
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 7009 3111 7067 3117
rect 7009 3108 7021 3111
rect 5776 3080 7021 3108
rect 5776 3068 5782 3080
rect 7009 3077 7021 3080
rect 7055 3077 7067 3111
rect 7009 3071 7067 3077
rect 7190 3040 7196 3052
rect 5276 3012 7196 3040
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 8076 3012 8217 3040
rect 8076 3000 8082 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10042 3040 10048 3052
rect 9907 3012 10048 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 3970 2972 3976 2984
rect 3743 2944 3832 2972
rect 3931 2944 3976 2972
rect 3743 2941 3755 2944
rect 3697 2935 3755 2941
rect 3970 2932 3976 2944
rect 4028 2932 4034 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 6730 2972 6736 2984
rect 4203 2944 6736 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 6914 2972 6920 2984
rect 6871 2944 6920 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 6914 2932 6920 2944
rect 6972 2972 6978 2984
rect 7374 2972 7380 2984
rect 6972 2944 7380 2972
rect 6972 2932 6978 2944
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 10778 2932 10784 2984
rect 10836 2972 10842 2984
rect 12504 2975 12562 2981
rect 12504 2972 12516 2975
rect 10836 2944 12516 2972
rect 10836 2932 10842 2944
rect 12504 2941 12516 2944
rect 12550 2972 12562 2975
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12550 2944 12909 2972
rect 12550 2941 12562 2944
rect 12504 2935 12562 2941
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 5306 2907 5364 2913
rect 5306 2873 5318 2907
rect 5352 2904 5364 2907
rect 6178 2904 6184 2916
rect 5352 2876 6184 2904
rect 5352 2873 5364 2876
rect 5306 2867 5364 2873
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 4798 2836 4804 2848
rect 1820 2808 4804 2836
rect 1820 2796 1826 2808
rect 4798 2796 4804 2808
rect 4856 2836 4862 2848
rect 5321 2836 5349 2867
rect 6178 2864 6184 2876
rect 6236 2864 6242 2916
rect 8526 2907 8584 2913
rect 8526 2873 8538 2907
rect 8572 2873 8584 2907
rect 10137 2907 10195 2913
rect 8526 2867 8584 2873
rect 9140 2876 9996 2904
rect 8018 2836 8024 2848
rect 4856 2808 5349 2836
rect 7979 2808 8024 2836
rect 4856 2796 4862 2808
rect 8018 2796 8024 2808
rect 8076 2836 8082 2848
rect 8541 2836 8569 2867
rect 9140 2845 9168 2876
rect 8076 2808 8569 2836
rect 9125 2839 9183 2845
rect 8076 2796 8082 2808
rect 9125 2805 9137 2839
rect 9171 2805 9183 2839
rect 9968 2836 9996 2876
rect 10137 2873 10149 2907
rect 10183 2873 10195 2907
rect 10137 2867 10195 2873
rect 10152 2836 10180 2867
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10376 2876 10701 2904
rect 10376 2864 10382 2876
rect 10689 2873 10701 2876
rect 10735 2904 10747 2907
rect 11054 2904 11060 2916
rect 10735 2876 11060 2904
rect 10735 2873 10747 2876
rect 10689 2867 10747 2873
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 9968 2808 10977 2836
rect 9125 2799 9183 2805
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 10965 2799 11023 2805
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12575 2839 12633 2845
rect 12575 2836 12587 2839
rect 12400 2808 12587 2836
rect 12400 2796 12406 2808
rect 12575 2805 12587 2808
rect 12621 2805 12633 2839
rect 12575 2799 12633 2805
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3970 2632 3976 2644
rect 3559 2604 3976 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4948 2604 5089 2632
rect 4948 2592 4954 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 5077 2595 5135 2601
rect 5460 2604 7849 2632
rect 5460 2573 5488 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 10410 2632 10416 2644
rect 10371 2604 10416 2632
rect 7837 2595 7895 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2564 3939 2567
rect 5445 2567 5503 2573
rect 5445 2564 5457 2567
rect 3927 2536 5457 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 5445 2533 5457 2536
rect 5491 2533 5503 2567
rect 5445 2527 5503 2533
rect 6365 2567 6423 2573
rect 6365 2533 6377 2567
rect 6411 2564 6423 2567
rect 6638 2564 6644 2576
rect 6411 2536 6644 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4203 2468 4844 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 4816 2369 4844 2468
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 6380 2428 6408 2527
rect 6638 2524 6644 2536
rect 6696 2524 6702 2576
rect 7190 2564 7196 2576
rect 7151 2536 7196 2564
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6788 2468 6929 2496
rect 6788 2456 6794 2468
rect 6917 2465 6929 2468
rect 6963 2496 6975 2499
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 6963 2468 8493 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8732 2499 8790 2505
rect 8732 2465 8744 2499
rect 8778 2496 8790 2499
rect 8846 2496 8852 2508
rect 8778 2468 8852 2496
rect 8778 2465 8790 2468
rect 8732 2459 8790 2465
rect 8846 2456 8852 2468
rect 8904 2496 8910 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8904 2468 9137 2496
rect 8904 2456 8910 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10428 2496 10456 2592
rect 9815 2468 10456 2496
rect 10873 2499 10931 2505
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10873 2465 10885 2499
rect 10919 2465 10931 2499
rect 10873 2459 10931 2465
rect 5399 2400 6408 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 10888 2428 10916 2459
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 12688 2499 12746 2505
rect 12688 2496 12700 2499
rect 11112 2468 12700 2496
rect 11112 2456 11118 2468
rect 12688 2465 12700 2468
rect 12734 2496 12746 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12734 2468 13093 2496
rect 12734 2465 12746 2468
rect 12688 2459 12746 2465
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13081 2459 13139 2465
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 7064 2400 11437 2428
rect 7064 2388 7070 2400
rect 11425 2397 11437 2400
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 4801 2363 4859 2369
rect 4801 2329 4813 2363
rect 4847 2360 4859 2363
rect 5534 2360 5540 2372
rect 4847 2332 5540 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 5902 2360 5908 2372
rect 5815 2332 5908 2360
rect 5902 2320 5908 2332
rect 5960 2360 5966 2372
rect 10778 2360 10784 2372
rect 5960 2332 10784 2360
rect 5960 2320 5966 2332
rect 10778 2320 10784 2332
rect 10836 2320 10842 2372
rect 12759 2363 12817 2369
rect 12759 2329 12771 2363
rect 12805 2360 12817 2363
rect 13354 2360 13360 2372
rect 12805 2332 13360 2360
rect 12805 2329 12817 2332
rect 12759 2323 12817 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 4522 2292 4528 2304
rect 4387 2264 4528 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6236 2264 6653 2292
rect 6236 2252 6242 2264
rect 6641 2261 6653 2264
rect 6687 2292 6699 2295
rect 7190 2292 7196 2304
rect 6687 2264 7196 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 7190 2252 7196 2264
rect 7248 2292 7254 2304
rect 8018 2292 8024 2304
rect 7248 2264 8024 2292
rect 7248 2252 7254 2264
rect 8018 2252 8024 2264
rect 8076 2292 8082 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 8076 2264 8125 2292
rect 8076 2252 8082 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8803 2295 8861 2301
rect 8803 2261 8815 2295
rect 8849 2292 8861 2295
rect 9766 2292 9772 2304
rect 8849 2264 9772 2292
rect 8849 2261 8861 2264
rect 8803 2255 8861 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 11054 2292 11060 2304
rect 11015 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
<< via1 >>
rect 572 39584 624 39636
rect 1216 39584 1268 39636
rect 2780 39584 2832 39636
rect 3516 39584 3568 39636
rect 13820 39584 13872 39636
rect 15384 39584 15436 39636
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 10048 35819 10100 35828
rect 10048 35785 10057 35819
rect 10057 35785 10091 35819
rect 10091 35785 10100 35819
rect 10048 35776 10100 35785
rect 5540 35572 5592 35624
rect 9312 35572 9364 35624
rect 5356 35504 5408 35556
rect 6736 35504 6788 35556
rect 8300 35547 8352 35556
rect 8300 35513 8309 35547
rect 8309 35513 8343 35547
rect 8343 35513 8352 35547
rect 8300 35504 8352 35513
rect 8392 35547 8444 35556
rect 8392 35513 8401 35547
rect 8401 35513 8435 35547
rect 8435 35513 8444 35547
rect 8392 35504 8444 35513
rect 6828 35436 6880 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 6828 35275 6880 35284
rect 6828 35241 6837 35275
rect 6837 35241 6871 35275
rect 6871 35241 6880 35275
rect 6828 35232 6880 35241
rect 8300 35232 8352 35284
rect 10508 35232 10560 35284
rect 7012 35164 7064 35216
rect 6184 35096 6236 35148
rect 9680 35139 9732 35148
rect 9680 35105 9689 35139
rect 9689 35105 9723 35139
rect 9723 35105 9732 35139
rect 9680 35096 9732 35105
rect 9772 35028 9824 35080
rect 8300 34935 8352 34944
rect 8300 34901 8309 34935
rect 8309 34901 8343 34935
rect 8343 34901 8352 34935
rect 8300 34892 8352 34901
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 5540 34731 5592 34740
rect 5540 34697 5549 34731
rect 5549 34697 5583 34731
rect 5583 34697 5592 34731
rect 5540 34688 5592 34697
rect 5724 34688 5776 34740
rect 6184 34731 6236 34740
rect 6184 34697 6193 34731
rect 6193 34697 6227 34731
rect 6227 34697 6236 34731
rect 6184 34688 6236 34697
rect 6736 34688 6788 34740
rect 9680 34731 9732 34740
rect 9680 34697 9689 34731
rect 9689 34697 9723 34731
rect 9723 34697 9732 34731
rect 9680 34688 9732 34697
rect 9956 34688 10008 34740
rect 12808 34688 12860 34740
rect 7104 34620 7156 34672
rect 7564 34663 7616 34672
rect 7564 34629 7573 34663
rect 7573 34629 7607 34663
rect 7607 34629 7616 34663
rect 7564 34620 7616 34629
rect 6828 34552 6880 34604
rect 8576 34595 8628 34604
rect 8576 34561 8585 34595
rect 8585 34561 8619 34595
rect 8619 34561 8628 34595
rect 8576 34552 8628 34561
rect 9312 34552 9364 34604
rect 5540 34484 5592 34536
rect 6000 34484 6052 34536
rect 10048 34527 10100 34536
rect 10048 34493 10057 34527
rect 10057 34493 10091 34527
rect 10091 34493 10100 34527
rect 10048 34484 10100 34493
rect 11244 34484 11296 34536
rect 7012 34416 7064 34468
rect 8668 34459 8720 34468
rect 8668 34425 8677 34459
rect 8677 34425 8711 34459
rect 8711 34425 8720 34459
rect 8668 34416 8720 34425
rect 7932 34391 7984 34400
rect 7932 34357 7941 34391
rect 7941 34357 7975 34391
rect 7975 34357 7984 34391
rect 7932 34348 7984 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 8300 34187 8352 34196
rect 8300 34153 8309 34187
rect 8309 34153 8343 34187
rect 8343 34153 8352 34187
rect 8300 34144 8352 34153
rect 8576 34187 8628 34196
rect 8576 34153 8585 34187
rect 8585 34153 8619 34187
rect 8619 34153 8628 34187
rect 8576 34144 8628 34153
rect 7472 34076 7524 34128
rect 9588 34076 9640 34128
rect 6092 34051 6144 34060
rect 6092 34017 6101 34051
rect 6101 34017 6135 34051
rect 6135 34017 6144 34051
rect 6092 34008 6144 34017
rect 6276 34051 6328 34060
rect 6276 34017 6285 34051
rect 6285 34017 6319 34051
rect 6319 34017 6328 34051
rect 6276 34008 6328 34017
rect 7932 34008 7984 34060
rect 4804 33983 4856 33992
rect 4804 33949 4813 33983
rect 4813 33949 4847 33983
rect 4847 33949 4856 33983
rect 4804 33940 4856 33949
rect 9772 33983 9824 33992
rect 9772 33949 9781 33983
rect 9781 33949 9815 33983
rect 9815 33949 9824 33983
rect 9772 33940 9824 33949
rect 9312 33872 9364 33924
rect 7012 33847 7064 33856
rect 7012 33813 7021 33847
rect 7021 33813 7055 33847
rect 7055 33813 7064 33847
rect 7012 33804 7064 33813
rect 8392 33804 8444 33856
rect 10048 33804 10100 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6276 33600 6328 33652
rect 7012 33600 7064 33652
rect 8668 33600 8720 33652
rect 9772 33600 9824 33652
rect 4068 33532 4120 33584
rect 3976 33328 4028 33380
rect 9312 33532 9364 33584
rect 4620 33328 4672 33380
rect 4712 33303 4764 33312
rect 4712 33269 4721 33303
rect 4721 33269 4755 33303
rect 4755 33269 4764 33303
rect 4712 33260 4764 33269
rect 4988 33328 5040 33380
rect 6644 33396 6696 33448
rect 8576 33439 8628 33448
rect 6276 33328 6328 33380
rect 6920 33328 6972 33380
rect 8576 33405 8585 33439
rect 8585 33405 8619 33439
rect 8619 33405 8628 33439
rect 8576 33396 8628 33405
rect 7472 33328 7524 33380
rect 6092 33260 6144 33312
rect 8668 33260 8720 33312
rect 9588 33260 9640 33312
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 4620 33099 4672 33108
rect 4620 33065 4629 33099
rect 4629 33065 4663 33099
rect 4663 33065 4672 33099
rect 4620 33056 4672 33065
rect 7472 33099 7524 33108
rect 7472 33065 7481 33099
rect 7481 33065 7515 33099
rect 7515 33065 7524 33099
rect 7472 33056 7524 33065
rect 9588 33056 9640 33108
rect 4988 32988 5040 33040
rect 4804 32895 4856 32904
rect 4804 32861 4813 32895
rect 4813 32861 4847 32895
rect 4847 32861 4856 32895
rect 4804 32852 4856 32861
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 4344 32784 4396 32836
rect 8576 32827 8628 32836
rect 8576 32793 8585 32827
rect 8585 32793 8619 32827
rect 8619 32793 8628 32827
rect 8576 32784 8628 32793
rect 5356 32716 5408 32768
rect 6644 32716 6696 32768
rect 6920 32759 6972 32768
rect 6920 32725 6929 32759
rect 6929 32725 6963 32759
rect 6963 32725 6972 32759
rect 6920 32716 6972 32725
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 7472 32512 7524 32564
rect 4160 32444 4212 32496
rect 4344 32419 4396 32428
rect 4344 32385 4353 32419
rect 4353 32385 4387 32419
rect 4387 32385 4396 32419
rect 4344 32376 4396 32385
rect 4896 32376 4948 32428
rect 4068 32351 4120 32360
rect 4068 32317 4077 32351
rect 4077 32317 4111 32351
rect 4111 32317 4120 32351
rect 4068 32308 4120 32317
rect 6920 32376 6972 32428
rect 8668 32351 8720 32360
rect 8668 32317 8677 32351
rect 8677 32317 8711 32351
rect 8711 32317 8720 32351
rect 8668 32308 8720 32317
rect 4344 32240 4396 32292
rect 5356 32283 5408 32292
rect 5356 32249 5365 32283
rect 5365 32249 5399 32283
rect 5399 32249 5408 32283
rect 5356 32240 5408 32249
rect 7012 32240 7064 32292
rect 9680 32308 9732 32360
rect 10048 32308 10100 32360
rect 10232 32240 10284 32292
rect 4988 32172 5040 32224
rect 6644 32172 6696 32224
rect 8484 32215 8536 32224
rect 8484 32181 8493 32215
rect 8493 32181 8527 32215
rect 8527 32181 8536 32215
rect 8484 32172 8536 32181
rect 9680 32172 9732 32224
rect 10048 32215 10100 32224
rect 10048 32181 10057 32215
rect 10057 32181 10091 32215
rect 10091 32181 10100 32215
rect 10048 32172 10100 32181
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 3424 31968 3476 32020
rect 4068 31968 4120 32020
rect 4804 32011 4856 32020
rect 4804 31977 4813 32011
rect 4813 31977 4847 32011
rect 4847 31977 4856 32011
rect 4804 31968 4856 31977
rect 9772 32011 9824 32020
rect 9772 31977 9781 32011
rect 9781 31977 9815 32011
rect 9815 31977 9824 32011
rect 9772 31968 9824 31977
rect 14004 31968 14056 32020
rect 4988 31900 5040 31952
rect 6920 31943 6972 31952
rect 6920 31909 6929 31943
rect 6929 31909 6963 31943
rect 6963 31909 6972 31943
rect 6920 31900 6972 31909
rect 7104 31900 7156 31952
rect 10048 31900 10100 31952
rect 9680 31875 9732 31884
rect 9680 31841 9689 31875
rect 9689 31841 9723 31875
rect 9723 31841 9732 31875
rect 9680 31832 9732 31841
rect 10232 31875 10284 31884
rect 10232 31841 10241 31875
rect 10241 31841 10275 31875
rect 10275 31841 10284 31875
rect 10232 31832 10284 31841
rect 10968 31832 11020 31884
rect 11428 31832 11480 31884
rect 4620 31764 4672 31816
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 7012 31764 7064 31816
rect 5908 31671 5960 31680
rect 5908 31637 5917 31671
rect 5917 31637 5951 31671
rect 5951 31637 5960 31671
rect 5908 31628 5960 31637
rect 8668 31628 8720 31680
rect 9496 31628 9548 31680
rect 10140 31628 10192 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 5632 31424 5684 31476
rect 6828 31424 6880 31476
rect 11428 31467 11480 31476
rect 11428 31433 11437 31467
rect 11437 31433 11471 31467
rect 11471 31433 11480 31467
rect 11428 31424 11480 31433
rect 6920 31356 6972 31408
rect 10416 31356 10468 31408
rect 4988 31288 5040 31340
rect 9772 31288 9824 31340
rect 10140 31331 10192 31340
rect 10140 31297 10149 31331
rect 10149 31297 10183 31331
rect 10183 31297 10192 31331
rect 10140 31288 10192 31297
rect 3976 31220 4028 31272
rect 9680 31263 9732 31272
rect 4620 31084 4672 31136
rect 4988 31152 5040 31204
rect 9680 31229 9689 31263
rect 9689 31229 9723 31263
rect 9723 31229 9732 31263
rect 9680 31220 9732 31229
rect 5540 31084 5592 31136
rect 8116 31127 8168 31136
rect 8116 31093 8125 31127
rect 8125 31093 8159 31127
rect 8159 31093 8168 31127
rect 10232 31195 10284 31204
rect 10232 31161 10241 31195
rect 10241 31161 10275 31195
rect 10275 31161 10284 31195
rect 10232 31152 10284 31161
rect 8116 31084 8168 31093
rect 9588 31084 9640 31136
rect 10968 31084 11020 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 3976 30880 4028 30932
rect 4252 30812 4304 30864
rect 3976 30744 4028 30796
rect 5908 30812 5960 30864
rect 8116 30880 8168 30932
rect 10232 30880 10284 30932
rect 7012 30812 7064 30864
rect 9864 30855 9916 30864
rect 9864 30821 9873 30855
rect 9873 30821 9907 30855
rect 9907 30821 9916 30855
rect 9864 30812 9916 30821
rect 10416 30855 10468 30864
rect 10416 30821 10425 30855
rect 10425 30821 10459 30855
rect 10459 30821 10468 30855
rect 10416 30812 10468 30821
rect 5356 30676 5408 30728
rect 7840 30719 7892 30728
rect 7840 30685 7849 30719
rect 7849 30685 7883 30719
rect 7883 30685 7892 30719
rect 7840 30676 7892 30685
rect 9772 30719 9824 30728
rect 9772 30685 9781 30719
rect 9781 30685 9815 30719
rect 9815 30685 9824 30719
rect 9772 30676 9824 30685
rect 4988 30583 5040 30592
rect 4988 30549 4997 30583
rect 4997 30549 5031 30583
rect 5031 30549 5040 30583
rect 4988 30540 5040 30549
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 3976 30336 4028 30388
rect 4068 30336 4120 30388
rect 5908 30336 5960 30388
rect 9772 30379 9824 30388
rect 9772 30345 9781 30379
rect 9781 30345 9815 30379
rect 9815 30345 9824 30379
rect 9772 30336 9824 30345
rect 9864 30336 9916 30388
rect 4988 30268 5040 30320
rect 8116 30311 8168 30320
rect 8116 30277 8125 30311
rect 8125 30277 8159 30311
rect 8159 30277 8168 30311
rect 8116 30268 8168 30277
rect 4344 30132 4396 30184
rect 7012 30200 7064 30252
rect 8484 30200 8536 30252
rect 10416 30243 10468 30252
rect 10416 30209 10425 30243
rect 10425 30209 10459 30243
rect 10459 30209 10468 30243
rect 10416 30200 10468 30209
rect 4436 30064 4488 30116
rect 6736 30132 6788 30184
rect 8116 30064 8168 30116
rect 10140 30107 10192 30116
rect 10140 30073 10149 30107
rect 10149 30073 10183 30107
rect 10183 30073 10192 30107
rect 10140 30064 10192 30073
rect 4620 29996 4672 30048
rect 5356 29996 5408 30048
rect 6828 29996 6880 30048
rect 9588 29996 9640 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 4160 29835 4212 29844
rect 4160 29801 4169 29835
rect 4169 29801 4203 29835
rect 4203 29801 4212 29835
rect 4160 29792 4212 29801
rect 8484 29792 8536 29844
rect 6828 29767 6880 29776
rect 6828 29733 6837 29767
rect 6837 29733 6871 29767
rect 6871 29733 6880 29767
rect 6828 29724 6880 29733
rect 7104 29767 7156 29776
rect 7104 29733 7113 29767
rect 7113 29733 7147 29767
rect 7147 29733 7156 29767
rect 7104 29724 7156 29733
rect 7840 29724 7892 29776
rect 10140 29792 10192 29844
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 4436 29656 4488 29708
rect 4620 29656 4672 29708
rect 5908 29699 5960 29708
rect 5908 29665 5952 29699
rect 5952 29665 5960 29699
rect 5908 29656 5960 29665
rect 8668 29656 8720 29708
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9680 29656 9732 29665
rect 9864 29656 9916 29708
rect 10968 29656 11020 29708
rect 9312 29588 9364 29640
rect 6920 29452 6972 29504
rect 8484 29452 8536 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 5908 29291 5960 29300
rect 5908 29257 5917 29291
rect 5917 29257 5951 29291
rect 5951 29257 5960 29291
rect 5908 29248 5960 29257
rect 7012 29180 7064 29232
rect 9680 29223 9732 29232
rect 9680 29189 9689 29223
rect 9689 29189 9723 29223
rect 9723 29189 9732 29223
rect 9680 29180 9732 29189
rect 4160 29155 4212 29164
rect 4160 29121 4169 29155
rect 4169 29121 4203 29155
rect 4203 29121 4212 29155
rect 6920 29155 6972 29164
rect 4160 29112 4212 29121
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 6920 29112 6972 29121
rect 7564 29155 7616 29164
rect 7564 29121 7573 29155
rect 7573 29121 7607 29155
rect 7607 29121 7616 29155
rect 7564 29112 7616 29121
rect 8300 29112 8352 29164
rect 8484 29155 8536 29164
rect 8484 29121 8493 29155
rect 8493 29121 8527 29155
rect 8527 29121 8536 29155
rect 8484 29112 8536 29121
rect 9312 29112 9364 29164
rect 4988 28976 5040 29028
rect 3884 28908 3936 28960
rect 5080 28951 5132 28960
rect 5080 28917 5089 28951
rect 5089 28917 5123 28951
rect 5123 28917 5132 28951
rect 5080 28908 5132 28917
rect 8116 28976 8168 29028
rect 7104 28908 7156 28960
rect 8668 28908 8720 28960
rect 9588 28908 9640 28960
rect 9864 28908 9916 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 1584 28747 1636 28756
rect 1584 28713 1593 28747
rect 1593 28713 1627 28747
rect 1627 28713 1636 28747
rect 1584 28704 1636 28713
rect 4436 28704 4488 28756
rect 4988 28704 5040 28756
rect 6184 28704 6236 28756
rect 5080 28636 5132 28688
rect 6920 28704 6972 28756
rect 8116 28679 8168 28688
rect 8116 28645 8125 28679
rect 8125 28645 8159 28679
rect 8159 28645 8168 28679
rect 8116 28636 8168 28645
rect 1400 28611 1452 28620
rect 1400 28577 1409 28611
rect 1409 28577 1443 28611
rect 1443 28577 1452 28611
rect 1400 28568 1452 28577
rect 2688 28568 2740 28620
rect 7104 28611 7156 28620
rect 7104 28577 7113 28611
rect 7113 28577 7147 28611
rect 7147 28577 7156 28611
rect 7104 28568 7156 28577
rect 9772 28611 9824 28620
rect 9772 28577 9790 28611
rect 9790 28577 9824 28611
rect 9772 28568 9824 28577
rect 11060 28568 11112 28620
rect 4344 28500 4396 28552
rect 5356 28543 5408 28552
rect 5356 28509 5365 28543
rect 5365 28509 5399 28543
rect 5399 28509 5408 28543
rect 5356 28500 5408 28509
rect 6092 28500 6144 28552
rect 6736 28432 6788 28484
rect 8300 28543 8352 28552
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 3976 28364 4028 28416
rect 4436 28364 4488 28416
rect 4988 28364 5040 28416
rect 7748 28407 7800 28416
rect 7748 28373 7757 28407
rect 7757 28373 7791 28407
rect 7791 28373 7800 28407
rect 7748 28364 7800 28373
rect 9956 28364 10008 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 5080 28160 5132 28212
rect 6184 28203 6236 28212
rect 6184 28169 6193 28203
rect 6193 28169 6227 28203
rect 6227 28169 6236 28203
rect 6184 28160 6236 28169
rect 7748 28160 7800 28212
rect 9772 28203 9824 28212
rect 9772 28169 9781 28203
rect 9781 28169 9815 28203
rect 9815 28169 9824 28203
rect 9772 28160 9824 28169
rect 1400 27956 1452 28008
rect 4620 28092 4672 28144
rect 4988 28067 5040 28076
rect 4988 28033 4997 28067
rect 4997 28033 5031 28067
rect 5031 28033 5040 28067
rect 4988 28024 5040 28033
rect 5632 28067 5684 28076
rect 5632 28033 5641 28067
rect 5641 28033 5675 28067
rect 5675 28033 5684 28067
rect 5632 28024 5684 28033
rect 2596 27888 2648 27940
rect 3700 27863 3752 27872
rect 3700 27829 3709 27863
rect 3709 27829 3743 27863
rect 3743 27829 3752 27863
rect 3700 27820 3752 27829
rect 4252 27820 4304 27872
rect 5080 27931 5132 27940
rect 5080 27897 5089 27931
rect 5089 27897 5123 27931
rect 5123 27897 5132 27931
rect 5080 27888 5132 27897
rect 6092 27888 6144 27940
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 10140 28024 10192 28076
rect 8760 27956 8812 28008
rect 10048 27931 10100 27940
rect 10048 27897 10057 27931
rect 10057 27897 10091 27931
rect 10091 27897 10100 27931
rect 10048 27888 10100 27897
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3976 27616 4028 27668
rect 4344 27659 4396 27668
rect 4344 27625 4353 27659
rect 4353 27625 4387 27659
rect 4387 27625 4396 27659
rect 4344 27616 4396 27625
rect 5080 27616 5132 27668
rect 8116 27616 8168 27668
rect 11520 27616 11572 27668
rect 4068 27548 4120 27600
rect 4988 27548 5040 27600
rect 6092 27548 6144 27600
rect 6184 27548 6236 27600
rect 8392 27548 8444 27600
rect 10048 27548 10100 27600
rect 11060 27548 11112 27600
rect 4804 27523 4856 27532
rect 4804 27489 4813 27523
rect 4813 27489 4847 27523
rect 4847 27489 4856 27523
rect 4804 27480 4856 27489
rect 5264 27523 5316 27532
rect 5264 27489 5273 27523
rect 5273 27489 5307 27523
rect 5307 27489 5316 27523
rect 5264 27480 5316 27489
rect 11428 27523 11480 27532
rect 11428 27489 11437 27523
rect 11437 27489 11471 27523
rect 11471 27489 11480 27523
rect 11428 27480 11480 27489
rect 4712 27412 4764 27464
rect 7932 27412 7984 27464
rect 9404 27412 9456 27464
rect 10232 27455 10284 27464
rect 10232 27421 10241 27455
rect 10241 27421 10275 27455
rect 10275 27421 10284 27455
rect 10232 27412 10284 27421
rect 2688 27344 2740 27396
rect 3700 27344 3752 27396
rect 4436 27344 4488 27396
rect 6000 27344 6052 27396
rect 8760 27387 8812 27396
rect 8760 27353 8769 27387
rect 8769 27353 8803 27387
rect 8803 27353 8812 27387
rect 8760 27344 8812 27353
rect 9956 27344 10008 27396
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 8852 27276 8904 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 3148 27072 3200 27124
rect 4436 27072 4488 27124
rect 3424 27004 3476 27056
rect 5264 27072 5316 27124
rect 5448 27072 5500 27124
rect 6184 27072 6236 27124
rect 7932 27115 7984 27124
rect 7932 27081 7941 27115
rect 7941 27081 7975 27115
rect 7975 27081 7984 27115
rect 7932 27072 7984 27081
rect 8392 27115 8444 27124
rect 8392 27081 8401 27115
rect 8401 27081 8435 27115
rect 8435 27081 8444 27115
rect 8392 27072 8444 27081
rect 11060 27115 11112 27124
rect 11060 27081 11069 27115
rect 11069 27081 11103 27115
rect 11103 27081 11112 27115
rect 11060 27072 11112 27081
rect 4804 27004 4856 27056
rect 4252 26936 4304 26988
rect 5816 26936 5868 26988
rect 7748 27004 7800 27056
rect 8852 26936 8904 26988
rect 10232 26936 10284 26988
rect 3976 26911 4028 26920
rect 3976 26877 3985 26911
rect 3985 26877 4019 26911
rect 4019 26877 4028 26911
rect 3976 26868 4028 26877
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 4344 26800 4396 26852
rect 5172 26843 5224 26852
rect 5172 26809 5181 26843
rect 5181 26809 5215 26843
rect 5215 26809 5224 26843
rect 5172 26800 5224 26809
rect 5356 26800 5408 26852
rect 6644 26800 6696 26852
rect 4804 26732 4856 26784
rect 5264 26732 5316 26784
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 7656 26843 7708 26852
rect 7656 26809 7665 26843
rect 7665 26809 7699 26843
rect 7699 26809 7708 26843
rect 7656 26800 7708 26809
rect 8668 26843 8720 26852
rect 8668 26809 8677 26843
rect 8677 26809 8711 26843
rect 8711 26809 8720 26843
rect 8668 26800 8720 26809
rect 9864 26800 9916 26852
rect 6000 26732 6052 26741
rect 9956 26732 10008 26784
rect 11428 26775 11480 26784
rect 11428 26741 11437 26775
rect 11437 26741 11471 26775
rect 11471 26741 11480 26775
rect 11428 26732 11480 26741
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 3424 26571 3476 26580
rect 3424 26537 3433 26571
rect 3433 26537 3467 26571
rect 3467 26537 3476 26571
rect 3424 26528 3476 26537
rect 3976 26528 4028 26580
rect 4252 26528 4304 26580
rect 6920 26528 6972 26580
rect 8668 26528 8720 26580
rect 9404 26571 9456 26580
rect 9404 26537 9413 26571
rect 9413 26537 9447 26571
rect 9447 26537 9456 26571
rect 9404 26528 9456 26537
rect 4528 26460 4580 26512
rect 5448 26460 5500 26512
rect 6276 26503 6328 26512
rect 6276 26469 6285 26503
rect 6285 26469 6319 26503
rect 6319 26469 6328 26503
rect 6276 26460 6328 26469
rect 7932 26460 7984 26512
rect 9864 26503 9916 26512
rect 9864 26469 9873 26503
rect 9873 26469 9907 26503
rect 9907 26469 9916 26503
rect 9864 26460 9916 26469
rect 10232 26460 10284 26512
rect 2044 26392 2096 26444
rect 3056 26392 3108 26444
rect 11428 26460 11480 26512
rect 4344 26367 4396 26376
rect 4344 26333 4353 26367
rect 4353 26333 4387 26367
rect 4387 26333 4396 26367
rect 4344 26324 4396 26333
rect 6644 26367 6696 26376
rect 6644 26333 6653 26367
rect 6653 26333 6687 26367
rect 6687 26333 6696 26367
rect 6644 26324 6696 26333
rect 7840 26367 7892 26376
rect 7840 26333 7849 26367
rect 7849 26333 7883 26367
rect 7883 26333 7892 26367
rect 7840 26324 7892 26333
rect 10876 26324 10928 26376
rect 6460 26256 6512 26308
rect 3332 26188 3384 26240
rect 5172 26188 5224 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4528 26027 4580 26036
rect 2044 25959 2096 25968
rect 2044 25925 2053 25959
rect 2053 25925 2087 25959
rect 2087 25925 2096 25959
rect 2044 25916 2096 25925
rect 4528 25993 4537 26027
rect 4537 25993 4571 26027
rect 4571 25993 4580 26027
rect 4528 25984 4580 25993
rect 4620 25984 4672 26036
rect 5724 25984 5776 26036
rect 6276 25984 6328 26036
rect 6460 26027 6512 26036
rect 6460 25993 6469 26027
rect 6469 25993 6503 26027
rect 6503 25993 6512 26027
rect 6460 25984 6512 25993
rect 8668 25984 8720 26036
rect 10048 25984 10100 26036
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 5264 25916 5316 25968
rect 5632 25959 5684 25968
rect 5632 25925 5641 25959
rect 5641 25925 5675 25959
rect 5675 25925 5684 25959
rect 5632 25916 5684 25925
rect 1768 25848 1820 25900
rect 2964 25848 3016 25900
rect 3332 25848 3384 25900
rect 2412 25823 2464 25832
rect 2412 25789 2421 25823
rect 2421 25789 2455 25823
rect 2455 25789 2464 25823
rect 2412 25780 2464 25789
rect 3884 25823 3936 25832
rect 3884 25789 3893 25823
rect 3893 25789 3927 25823
rect 3927 25789 3936 25823
rect 3884 25780 3936 25789
rect 4712 25780 4764 25832
rect 3976 25712 4028 25764
rect 7656 25848 7708 25900
rect 8944 25848 8996 25900
rect 10140 25848 10192 25900
rect 5816 25780 5868 25832
rect 5080 25755 5132 25764
rect 3056 25687 3108 25696
rect 3056 25653 3065 25687
rect 3065 25653 3099 25687
rect 3099 25653 3108 25687
rect 3056 25644 3108 25653
rect 5080 25721 5089 25755
rect 5089 25721 5123 25755
rect 5123 25721 5132 25755
rect 5080 25712 5132 25721
rect 5172 25755 5224 25764
rect 5172 25721 5181 25755
rect 5181 25721 5215 25755
rect 5215 25721 5224 25755
rect 5172 25712 5224 25721
rect 9956 25755 10008 25764
rect 4252 25644 4304 25696
rect 4712 25644 4764 25696
rect 7196 25644 7248 25696
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 9956 25721 9965 25755
rect 9965 25721 9999 25755
rect 9999 25721 10008 25755
rect 9956 25712 10008 25721
rect 10048 25755 10100 25764
rect 10048 25721 10057 25755
rect 10057 25721 10091 25755
rect 10091 25721 10100 25755
rect 10048 25712 10100 25721
rect 7932 25644 7984 25653
rect 9404 25687 9456 25696
rect 9404 25653 9413 25687
rect 9413 25653 9447 25687
rect 9447 25653 9456 25687
rect 9404 25644 9456 25653
rect 11428 25644 11480 25696
rect 12164 25644 12216 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 3884 25440 3936 25492
rect 4344 25483 4396 25492
rect 4344 25449 4353 25483
rect 4353 25449 4387 25483
rect 4387 25449 4396 25483
rect 4344 25440 4396 25449
rect 5080 25440 5132 25492
rect 8852 25440 8904 25492
rect 8944 25483 8996 25492
rect 8944 25449 8953 25483
rect 8953 25449 8987 25483
rect 8987 25449 8996 25483
rect 8944 25440 8996 25449
rect 9956 25440 10008 25492
rect 4528 25372 4580 25424
rect 7840 25372 7892 25424
rect 9404 25372 9456 25424
rect 9864 25415 9916 25424
rect 9864 25381 9873 25415
rect 9873 25381 9907 25415
rect 9907 25381 9916 25415
rect 9864 25372 9916 25381
rect 10416 25372 10468 25424
rect 3240 25304 3292 25356
rect 5264 25304 5316 25356
rect 6184 25304 6236 25356
rect 6920 25347 6972 25356
rect 6920 25313 6929 25347
rect 6929 25313 6963 25347
rect 6963 25313 6972 25347
rect 6920 25304 6972 25313
rect 3976 25236 4028 25288
rect 4620 25279 4672 25288
rect 4620 25245 4629 25279
rect 4629 25245 4663 25279
rect 4663 25245 4672 25279
rect 4620 25236 4672 25245
rect 4712 25236 4764 25288
rect 2412 25168 2464 25220
rect 4896 25168 4948 25220
rect 6000 25236 6052 25288
rect 8392 25304 8444 25356
rect 11244 25347 11296 25356
rect 11244 25313 11253 25347
rect 11253 25313 11287 25347
rect 11287 25313 11296 25347
rect 11244 25304 11296 25313
rect 9772 25279 9824 25288
rect 9772 25245 9781 25279
rect 9781 25245 9815 25279
rect 9815 25245 9824 25279
rect 9772 25236 9824 25245
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 6736 25168 6788 25220
rect 10508 25168 10560 25220
rect 6828 25143 6880 25152
rect 6828 25109 6837 25143
rect 6837 25109 6871 25143
rect 6871 25109 6880 25143
rect 6828 25100 6880 25109
rect 7104 25100 7156 25152
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4160 24939 4212 24948
rect 4160 24905 4169 24939
rect 4169 24905 4203 24939
rect 4203 24905 4212 24939
rect 4160 24896 4212 24905
rect 4528 24896 4580 24948
rect 9772 24896 9824 24948
rect 10416 24939 10468 24948
rect 10416 24905 10425 24939
rect 10425 24905 10459 24939
rect 10459 24905 10468 24939
rect 10416 24896 10468 24905
rect 11244 24939 11296 24948
rect 11244 24905 11253 24939
rect 11253 24905 11287 24939
rect 11287 24905 11296 24939
rect 11244 24896 11296 24905
rect 4068 24828 4120 24880
rect 4436 24828 4488 24880
rect 3884 24692 3936 24744
rect 4068 24692 4120 24744
rect 5816 24828 5868 24880
rect 6000 24828 6052 24880
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 6828 24760 6880 24812
rect 8484 24692 8536 24744
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 2228 24624 2280 24676
rect 5172 24667 5224 24676
rect 5172 24633 5181 24667
rect 5181 24633 5215 24667
rect 5215 24633 5224 24667
rect 5172 24624 5224 24633
rect 5264 24667 5316 24676
rect 5264 24633 5273 24667
rect 5273 24633 5307 24667
rect 5307 24633 5316 24667
rect 5264 24624 5316 24633
rect 5540 24624 5592 24676
rect 6000 24624 6052 24676
rect 7748 24667 7800 24676
rect 3240 24556 3292 24608
rect 3884 24599 3936 24608
rect 3884 24565 3893 24599
rect 3893 24565 3927 24599
rect 3927 24565 3936 24599
rect 3884 24556 3936 24565
rect 4988 24556 5040 24608
rect 5356 24556 5408 24608
rect 6920 24556 6972 24608
rect 7748 24633 7757 24667
rect 7757 24633 7791 24667
rect 7791 24633 7800 24667
rect 7748 24624 7800 24633
rect 7932 24624 7984 24676
rect 8392 24667 8444 24676
rect 8392 24633 8401 24667
rect 8401 24633 8435 24667
rect 8435 24633 8444 24667
rect 8392 24624 8444 24633
rect 9312 24624 9364 24676
rect 8024 24599 8076 24608
rect 8024 24565 8033 24599
rect 8033 24565 8067 24599
rect 8067 24565 8076 24599
rect 8024 24556 8076 24565
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 2504 24352 2556 24404
rect 4620 24352 4672 24404
rect 5264 24352 5316 24404
rect 6828 24352 6880 24404
rect 5172 24284 5224 24336
rect 8024 24284 8076 24336
rect 2228 24216 2280 24268
rect 2872 24216 2924 24268
rect 3976 24216 4028 24268
rect 4712 24216 4764 24268
rect 2044 24148 2096 24200
rect 4436 24148 4488 24200
rect 5908 24216 5960 24268
rect 6276 24259 6328 24268
rect 6276 24225 6320 24259
rect 6320 24225 6328 24259
rect 6276 24216 6328 24225
rect 7840 24148 7892 24200
rect 8852 24148 8904 24200
rect 4528 24080 4580 24132
rect 7104 24080 7156 24132
rect 1768 24012 1820 24064
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 5632 24012 5684 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 1676 23808 1728 23860
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 4804 23808 4856 23860
rect 3516 23783 3568 23792
rect 3516 23749 3525 23783
rect 3525 23749 3559 23783
rect 3559 23749 3568 23783
rect 3516 23740 3568 23749
rect 1768 23604 1820 23656
rect 2504 23604 2556 23656
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 3056 23468 3108 23520
rect 3424 23647 3476 23656
rect 3424 23613 3433 23647
rect 3433 23613 3467 23647
rect 3467 23613 3476 23647
rect 3424 23604 3476 23613
rect 4528 23672 4580 23724
rect 4804 23672 4856 23724
rect 5540 23808 5592 23860
rect 6276 23851 6328 23860
rect 6276 23817 6285 23851
rect 6285 23817 6319 23851
rect 6319 23817 6328 23851
rect 6276 23808 6328 23817
rect 15476 23808 15528 23860
rect 7840 23740 7892 23792
rect 8668 23715 8720 23724
rect 8668 23681 8677 23715
rect 8677 23681 8711 23715
rect 8711 23681 8720 23715
rect 8668 23672 8720 23681
rect 8852 23672 8904 23724
rect 5080 23604 5132 23656
rect 5632 23647 5684 23656
rect 5632 23613 5641 23647
rect 5641 23613 5675 23647
rect 5675 23613 5684 23647
rect 5632 23604 5684 23613
rect 6828 23647 6880 23656
rect 6828 23613 6837 23647
rect 6837 23613 6871 23647
rect 6871 23613 6880 23647
rect 6828 23604 6880 23613
rect 8208 23604 8260 23656
rect 10048 23604 10100 23656
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 13084 23604 13136 23656
rect 4252 23536 4304 23588
rect 6184 23536 6236 23588
rect 8392 23536 8444 23588
rect 3424 23468 3476 23520
rect 4712 23468 4764 23520
rect 7104 23468 7156 23520
rect 8024 23511 8076 23520
rect 8024 23477 8033 23511
rect 8033 23477 8067 23511
rect 8067 23477 8076 23511
rect 8024 23468 8076 23477
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 4436 23307 4488 23316
rect 4436 23273 4445 23307
rect 4445 23273 4479 23307
rect 4479 23273 4488 23307
rect 4436 23264 4488 23273
rect 7840 23307 7892 23316
rect 7840 23273 7849 23307
rect 7849 23273 7883 23307
rect 7883 23273 7892 23307
rect 7840 23264 7892 23273
rect 1676 23196 1728 23248
rect 4988 23196 5040 23248
rect 5540 23196 5592 23248
rect 6644 23239 6696 23248
rect 6644 23205 6647 23239
rect 6647 23205 6681 23239
rect 6681 23205 6696 23239
rect 6644 23196 6696 23205
rect 7104 23196 7156 23248
rect 8208 23239 8260 23248
rect 8208 23205 8217 23239
rect 8217 23205 8251 23239
rect 8251 23205 8260 23239
rect 8208 23196 8260 23205
rect 8852 23196 8904 23248
rect 9312 23196 9364 23248
rect 9772 23239 9824 23248
rect 9772 23205 9781 23239
rect 9781 23205 9815 23239
rect 9815 23205 9824 23239
rect 9772 23196 9824 23205
rect 9864 23239 9916 23248
rect 9864 23205 9873 23239
rect 9873 23205 9907 23239
rect 9907 23205 9916 23239
rect 9864 23196 9916 23205
rect 3148 23128 3200 23180
rect 4712 23171 4764 23180
rect 4712 23137 4721 23171
rect 4721 23137 4755 23171
rect 4755 23137 4764 23171
rect 4712 23128 4764 23137
rect 5632 23128 5684 23180
rect 7196 23128 7248 23180
rect 7288 23128 7340 23180
rect 7932 23128 7984 23180
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 6184 23060 6236 23112
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 8116 23060 8168 23069
rect 6736 22992 6788 23044
rect 8024 22992 8076 23044
rect 2964 22924 3016 22976
rect 3516 22924 3568 22976
rect 4344 22924 4396 22976
rect 5908 22924 5960 22976
rect 6828 22924 6880 22976
rect 8576 22924 8628 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 1676 22763 1728 22772
rect 1676 22729 1685 22763
rect 1685 22729 1719 22763
rect 1719 22729 1728 22763
rect 1676 22720 1728 22729
rect 4068 22720 4120 22772
rect 4712 22763 4764 22772
rect 4712 22729 4721 22763
rect 4721 22729 4755 22763
rect 4755 22729 4764 22763
rect 4712 22720 4764 22729
rect 6644 22763 6696 22772
rect 6644 22729 6653 22763
rect 6653 22729 6687 22763
rect 6687 22729 6696 22763
rect 6644 22720 6696 22729
rect 8392 22720 8444 22772
rect 9772 22720 9824 22772
rect 2964 22584 3016 22636
rect 3976 22584 4028 22636
rect 5448 22584 5500 22636
rect 7472 22584 7524 22636
rect 8668 22652 8720 22704
rect 9864 22584 9916 22636
rect 3332 22516 3384 22568
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 5632 22559 5684 22568
rect 5632 22525 5641 22559
rect 5641 22525 5675 22559
rect 5675 22525 5684 22559
rect 5632 22516 5684 22525
rect 5908 22559 5960 22568
rect 5908 22525 5917 22559
rect 5917 22525 5951 22559
rect 5951 22525 5960 22559
rect 5908 22516 5960 22525
rect 9588 22516 9640 22568
rect 10784 22559 10836 22568
rect 10784 22525 10793 22559
rect 10793 22525 10827 22559
rect 10827 22525 10836 22559
rect 10784 22516 10836 22525
rect 4344 22448 4396 22500
rect 7104 22448 7156 22500
rect 7932 22448 7984 22500
rect 8576 22448 8628 22500
rect 9496 22491 9548 22500
rect 2780 22380 2832 22432
rect 2964 22423 3016 22432
rect 2964 22389 2973 22423
rect 2973 22389 3007 22423
rect 3007 22389 3016 22423
rect 2964 22380 3016 22389
rect 3976 22380 4028 22432
rect 4712 22380 4764 22432
rect 6644 22380 6696 22432
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 9496 22457 9505 22491
rect 9505 22457 9539 22491
rect 9539 22457 9548 22491
rect 9496 22448 9548 22457
rect 8668 22380 8720 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 6184 22176 6236 22228
rect 7472 22219 7524 22228
rect 7472 22185 7481 22219
rect 7481 22185 7515 22219
rect 7515 22185 7524 22219
rect 7472 22176 7524 22185
rect 8116 22176 8168 22228
rect 13820 22176 13872 22228
rect 3332 22108 3384 22160
rect 3056 22083 3108 22092
rect 2412 21972 2464 22024
rect 3056 22049 3065 22083
rect 3065 22049 3099 22083
rect 3099 22049 3108 22083
rect 3056 22040 3108 22049
rect 4068 22040 4120 22092
rect 4620 22040 4672 22092
rect 6552 22108 6604 22160
rect 7932 22108 7984 22160
rect 8208 22151 8260 22160
rect 8208 22117 8217 22151
rect 8217 22117 8251 22151
rect 8251 22117 8260 22151
rect 8208 22108 8260 22117
rect 9864 22151 9916 22160
rect 9864 22117 9873 22151
rect 9873 22117 9907 22151
rect 9907 22117 9916 22151
rect 9864 22108 9916 22117
rect 5632 22040 5684 22092
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 112 21904 164 21956
rect 3148 21904 3200 21956
rect 4160 21904 4212 21956
rect 6368 21972 6420 22024
rect 6736 21972 6788 22024
rect 8852 21972 8904 22024
rect 10048 22015 10100 22024
rect 1400 21836 1452 21888
rect 2320 21836 2372 21888
rect 5172 21879 5224 21888
rect 5172 21845 5181 21879
rect 5181 21845 5215 21879
rect 5215 21845 5224 21879
rect 5172 21836 5224 21845
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 5632 21836 5684 21845
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 8760 21904 8812 21956
rect 9496 21904 9548 21956
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 9956 21836 10008 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 3056 21632 3108 21684
rect 4160 21675 4212 21684
rect 4160 21641 4169 21675
rect 4169 21641 4203 21675
rect 4203 21641 4212 21675
rect 4804 21675 4856 21684
rect 4160 21632 4212 21641
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 8208 21632 8260 21684
rect 8852 21632 8904 21684
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 4712 21564 4764 21616
rect 2044 21496 2096 21548
rect 9864 21564 9916 21616
rect 1216 21428 1268 21480
rect 1860 21428 1912 21480
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 3332 21471 3384 21480
rect 2228 21403 2280 21412
rect 2228 21369 2237 21403
rect 2237 21369 2271 21403
rect 2271 21369 2280 21403
rect 2228 21360 2280 21369
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 4068 21360 4120 21412
rect 4436 21360 4488 21412
rect 2964 21335 3016 21344
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 6368 21496 6420 21548
rect 4804 21428 4856 21480
rect 6920 21428 6972 21480
rect 7840 21428 7892 21480
rect 7104 21360 7156 21412
rect 8116 21360 8168 21412
rect 10324 21360 10376 21412
rect 11244 21360 11296 21412
rect 5816 21292 5868 21344
rect 9496 21335 9548 21344
rect 9496 21301 9505 21335
rect 9505 21301 9539 21335
rect 9539 21301 9548 21335
rect 9496 21292 9548 21301
rect 9588 21292 9640 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 1860 21131 1912 21140
rect 1860 21097 1869 21131
rect 1869 21097 1903 21131
rect 1903 21097 1912 21131
rect 1860 21088 1912 21097
rect 2228 21131 2280 21140
rect 2228 21097 2237 21131
rect 2237 21097 2271 21131
rect 2271 21097 2280 21131
rect 2228 21088 2280 21097
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 2412 20995 2464 21004
rect 2412 20961 2421 20995
rect 2421 20961 2455 20995
rect 2455 20961 2464 20995
rect 2412 20952 2464 20961
rect 3332 21088 3384 21140
rect 4896 21131 4948 21140
rect 4896 21097 4905 21131
rect 4905 21097 4939 21131
rect 4939 21097 4948 21131
rect 4896 21088 4948 21097
rect 6736 21088 6788 21140
rect 8116 21131 8168 21140
rect 8116 21097 8125 21131
rect 8125 21097 8159 21131
rect 8159 21097 8168 21131
rect 8116 21088 8168 21097
rect 8668 21131 8720 21140
rect 8668 21097 8677 21131
rect 8677 21097 8711 21131
rect 8711 21097 8720 21131
rect 8668 21088 8720 21097
rect 3240 21020 3292 21072
rect 6920 21063 6972 21072
rect 6920 21029 6929 21063
rect 6929 21029 6963 21063
rect 6963 21029 6972 21063
rect 6920 21020 6972 21029
rect 9496 21020 9548 21072
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 3056 20952 3108 21004
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 6184 20995 6236 21004
rect 4620 20884 4672 20936
rect 2228 20816 2280 20868
rect 4528 20859 4580 20868
rect 4528 20825 4537 20859
rect 4537 20825 4571 20859
rect 4571 20825 4580 20859
rect 4528 20816 4580 20825
rect 4436 20748 4488 20800
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 7196 20952 7248 21004
rect 9588 20952 9640 21004
rect 6000 20748 6052 20800
rect 7564 20791 7616 20800
rect 7564 20757 7573 20791
rect 7573 20757 7607 20791
rect 7607 20757 7616 20791
rect 10324 20859 10376 20868
rect 10324 20825 10333 20859
rect 10333 20825 10367 20859
rect 10367 20825 10376 20859
rect 10324 20816 10376 20825
rect 7564 20748 7616 20757
rect 8208 20748 8260 20800
rect 9772 20748 9824 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 3148 20544 3200 20596
rect 4068 20587 4120 20596
rect 4068 20553 4077 20587
rect 4077 20553 4111 20587
rect 4111 20553 4120 20587
rect 4068 20544 4120 20553
rect 4528 20544 4580 20596
rect 5632 20544 5684 20596
rect 7196 20544 7248 20596
rect 8116 20587 8168 20596
rect 8116 20553 8125 20587
rect 8125 20553 8159 20587
rect 8159 20553 8168 20587
rect 8116 20544 8168 20553
rect 9496 20544 9548 20596
rect 15476 20544 15528 20596
rect 4252 20476 4304 20528
rect 4620 20476 4672 20528
rect 5080 20476 5132 20528
rect 9864 20476 9916 20528
rect 1584 20408 1636 20460
rect 8208 20451 8260 20460
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 1676 20383 1728 20392
rect 1676 20349 1685 20383
rect 1685 20349 1719 20383
rect 1719 20349 1728 20383
rect 1676 20340 1728 20349
rect 2964 20340 3016 20392
rect 4068 20340 4120 20392
rect 4252 20383 4304 20392
rect 4252 20349 4261 20383
rect 4261 20349 4295 20383
rect 4295 20349 4304 20383
rect 4252 20340 4304 20349
rect 2136 20272 2188 20324
rect 2688 20272 2740 20324
rect 3424 20315 3476 20324
rect 3424 20281 3433 20315
rect 3433 20281 3467 20315
rect 3467 20281 3476 20315
rect 3424 20272 3476 20281
rect 2228 20247 2280 20256
rect 2228 20213 2237 20247
rect 2237 20213 2271 20247
rect 2271 20213 2280 20247
rect 2228 20204 2280 20213
rect 3148 20204 3200 20256
rect 4160 20204 4212 20256
rect 5172 20340 5224 20392
rect 6184 20383 6236 20392
rect 6184 20349 6193 20383
rect 6193 20349 6227 20383
rect 6227 20349 6236 20383
rect 6184 20340 6236 20349
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 8116 20340 8168 20392
rect 10784 20340 10836 20392
rect 4712 20272 4764 20324
rect 8024 20272 8076 20324
rect 6644 20204 6696 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 3424 20043 3476 20052
rect 3424 20009 3433 20043
rect 3433 20009 3467 20043
rect 3467 20009 3476 20043
rect 3424 20000 3476 20009
rect 4804 20043 4856 20052
rect 4804 20009 4813 20043
rect 4813 20009 4847 20043
rect 4847 20009 4856 20043
rect 4804 20000 4856 20009
rect 7196 20043 7248 20052
rect 7196 20009 7205 20043
rect 7205 20009 7239 20043
rect 7239 20009 7248 20043
rect 7196 20000 7248 20009
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 1676 19932 1728 19984
rect 3332 19932 3384 19984
rect 3516 19932 3568 19984
rect 4620 19932 4672 19984
rect 4896 19932 4948 19984
rect 8024 19932 8076 19984
rect 2596 19864 2648 19916
rect 4528 19864 4580 19916
rect 2228 19796 2280 19848
rect 3976 19796 4028 19848
rect 5816 19864 5868 19916
rect 6736 19864 6788 19916
rect 9404 19864 9456 19916
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 9496 19796 9548 19848
rect 4712 19728 4764 19780
rect 4804 19728 4856 19780
rect 1768 19660 1820 19712
rect 3240 19660 3292 19712
rect 4252 19660 4304 19712
rect 4436 19703 4488 19712
rect 4436 19669 4445 19703
rect 4445 19669 4479 19703
rect 4479 19669 4488 19703
rect 4436 19660 4488 19669
rect 5540 19660 5592 19712
rect 6000 19660 6052 19712
rect 7104 19660 7156 19712
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 4528 19456 4580 19508
rect 2596 19388 2648 19440
rect 3056 19388 3108 19440
rect 5816 19456 5868 19508
rect 10600 19456 10652 19508
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 1492 19295 1544 19304
rect 1492 19261 1501 19295
rect 1501 19261 1535 19295
rect 1535 19261 1544 19295
rect 1492 19252 1544 19261
rect 2872 19252 2924 19304
rect 1768 19184 1820 19236
rect 2320 19184 2372 19236
rect 3424 19252 3476 19304
rect 5264 19388 5316 19440
rect 6920 19388 6972 19440
rect 8024 19388 8076 19440
rect 8760 19388 8812 19440
rect 3700 19320 3752 19372
rect 4436 19320 4488 19372
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 3884 19252 3936 19304
rect 4804 19295 4856 19304
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 6000 19252 6052 19304
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 7196 19252 7248 19304
rect 4160 19184 4212 19236
rect 4988 19184 5040 19236
rect 8392 19184 8444 19236
rect 9496 19184 9548 19236
rect 3332 19116 3384 19168
rect 3976 19116 4028 19168
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 4712 19116 4764 19168
rect 5540 19116 5592 19168
rect 6736 19116 6788 19168
rect 8208 19116 8260 19168
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 9680 19116 9732 19125
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 1400 18912 1452 18964
rect 3056 18912 3108 18964
rect 6000 18955 6052 18964
rect 6000 18921 6009 18955
rect 6009 18921 6043 18955
rect 6043 18921 6052 18955
rect 6000 18912 6052 18921
rect 8392 18912 8444 18964
rect 9772 18955 9824 18964
rect 9772 18921 9781 18955
rect 9781 18921 9815 18955
rect 9815 18921 9824 18955
rect 9772 18912 9824 18921
rect 1584 18776 1636 18828
rect 5264 18844 5316 18896
rect 5540 18844 5592 18896
rect 2872 18776 2924 18828
rect 2964 18776 3016 18828
rect 6460 18776 6512 18828
rect 7472 18844 7524 18896
rect 7196 18776 7248 18828
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 8116 18776 8168 18785
rect 9496 18776 9548 18828
rect 10140 18819 10192 18828
rect 10140 18785 10149 18819
rect 10149 18785 10183 18819
rect 10183 18785 10192 18819
rect 10140 18776 10192 18785
rect 2320 18708 2372 18760
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 3424 18708 3476 18717
rect 3516 18708 3568 18760
rect 4344 18708 4396 18760
rect 5264 18708 5316 18760
rect 664 18572 716 18624
rect 1492 18572 1544 18624
rect 4068 18640 4120 18692
rect 4712 18640 4764 18692
rect 10140 18640 10192 18692
rect 4252 18572 4304 18624
rect 4988 18572 5040 18624
rect 10416 18572 10468 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 1952 18368 2004 18420
rect 2688 18368 2740 18420
rect 4068 18411 4120 18420
rect 2872 18300 2924 18352
rect 3240 18300 3292 18352
rect 4068 18377 4077 18411
rect 4077 18377 4111 18411
rect 4111 18377 4120 18411
rect 4068 18368 4120 18377
rect 4252 18368 4304 18420
rect 4804 18300 4856 18352
rect 1952 18164 2004 18216
rect 2780 18164 2832 18216
rect 3056 18164 3108 18216
rect 3976 18164 4028 18216
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 5356 18368 5408 18420
rect 8116 18411 8168 18420
rect 5448 18300 5500 18352
rect 6644 18300 6696 18352
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 10140 18411 10192 18420
rect 10140 18377 10149 18411
rect 10149 18377 10183 18411
rect 10183 18377 10192 18411
rect 10140 18368 10192 18377
rect 6460 18232 6512 18284
rect 9496 18232 9548 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 5540 18164 5592 18216
rect 5080 18096 5132 18148
rect 5264 18139 5316 18148
rect 5264 18105 5273 18139
rect 5273 18105 5307 18139
rect 5307 18105 5316 18139
rect 5264 18096 5316 18105
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 8852 18139 8904 18148
rect 8852 18105 8861 18139
rect 8861 18105 8895 18139
rect 8895 18105 8904 18139
rect 8852 18096 8904 18105
rect 7196 18028 7248 18080
rect 8300 18028 8352 18080
rect 10692 18096 10744 18148
rect 10600 18028 10652 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3056 17824 3108 17876
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 7380 17824 7432 17876
rect 9772 17824 9824 17876
rect 1768 17756 1820 17808
rect 2228 17756 2280 17808
rect 4988 17756 5040 17808
rect 5080 17756 5132 17808
rect 6000 17756 6052 17808
rect 6092 17756 6144 17808
rect 3148 17688 3200 17740
rect 9496 17756 9548 17808
rect 10140 17756 10192 17808
rect 7840 17731 7892 17740
rect 7840 17697 7849 17731
rect 7849 17697 7883 17731
rect 7883 17697 7892 17731
rect 7840 17688 7892 17697
rect 10508 17688 10560 17740
rect 11704 17688 11756 17740
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 4068 17620 4120 17672
rect 4896 17620 4948 17672
rect 4988 17620 5040 17672
rect 7012 17620 7064 17672
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 9864 17620 9916 17672
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 5356 17552 5408 17604
rect 6644 17552 6696 17604
rect 10692 17595 10744 17604
rect 2228 17484 2280 17536
rect 5816 17484 5868 17536
rect 6000 17484 6052 17536
rect 10692 17561 10701 17595
rect 10701 17561 10735 17595
rect 10735 17561 10744 17595
rect 10692 17552 10744 17561
rect 8852 17527 8904 17536
rect 8852 17493 8861 17527
rect 8861 17493 8895 17527
rect 8895 17493 8904 17527
rect 8852 17484 8904 17493
rect 10784 17484 10836 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 2320 17280 2372 17332
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 4988 17323 5040 17332
rect 4988 17289 4997 17323
rect 4997 17289 5031 17323
rect 5031 17289 5040 17323
rect 4988 17280 5040 17289
rect 8852 17280 8904 17332
rect 2136 17212 2188 17264
rect 2596 17144 2648 17196
rect 10324 17212 10376 17264
rect 11704 17255 11756 17264
rect 11704 17221 11713 17255
rect 11713 17221 11747 17255
rect 11747 17221 11756 17255
rect 11704 17212 11756 17221
rect 6644 17144 6696 17196
rect 6920 17144 6972 17196
rect 7380 17187 7432 17196
rect 4068 17076 4120 17128
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 6184 17076 6236 17128
rect 1400 17008 1452 17060
rect 2320 16940 2372 16992
rect 5356 17051 5408 17060
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 6092 17008 6144 17060
rect 6828 17008 6880 17060
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 9312 17144 9364 17196
rect 10416 17144 10468 17196
rect 11980 17076 12032 17128
rect 13084 17280 13136 17332
rect 13636 17323 13688 17332
rect 13636 17289 13645 17323
rect 13645 17289 13679 17323
rect 13679 17289 13688 17323
rect 13636 17280 13688 17289
rect 7472 17008 7524 17060
rect 7840 17008 7892 17060
rect 9864 17051 9916 17060
rect 3148 16940 3200 16992
rect 4252 16940 4304 16992
rect 4988 16940 5040 16992
rect 6000 16940 6052 16992
rect 8300 16983 8352 16992
rect 8300 16949 8309 16983
rect 8309 16949 8343 16983
rect 8343 16949 8352 16983
rect 8300 16940 8352 16949
rect 8484 16940 8536 16992
rect 9864 17017 9873 17051
rect 9873 17017 9907 17051
rect 9907 17017 9916 17051
rect 9864 17008 9916 17017
rect 10416 17008 10468 17060
rect 10600 17008 10652 17060
rect 9956 16940 10008 16992
rect 10140 16983 10192 16992
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 10968 17008 11020 17060
rect 10508 16940 10560 16949
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 1400 16779 1452 16788
rect 1400 16745 1409 16779
rect 1409 16745 1443 16779
rect 1443 16745 1452 16779
rect 1400 16736 1452 16745
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 10140 16736 10192 16788
rect 10600 16736 10652 16788
rect 3148 16668 3200 16720
rect 4252 16711 4304 16720
rect 4252 16677 4261 16711
rect 4261 16677 4295 16711
rect 4295 16677 4304 16711
rect 4252 16668 4304 16677
rect 5448 16668 5500 16720
rect 5908 16711 5960 16720
rect 5908 16677 5917 16711
rect 5917 16677 5951 16711
rect 5951 16677 5960 16711
rect 5908 16668 5960 16677
rect 6092 16668 6144 16720
rect 8300 16668 8352 16720
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 9956 16668 10008 16720
rect 11704 16668 11756 16720
rect 6644 16600 6696 16652
rect 9404 16600 9456 16652
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 2136 16532 2188 16584
rect 2596 16464 2648 16516
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4804 16575 4856 16584
rect 4160 16532 4212 16541
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 8576 16532 8628 16584
rect 4896 16464 4948 16516
rect 1584 16396 1636 16448
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 9312 16396 9364 16448
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 10784 16464 10836 16516
rect 12072 16396 12124 16448
rect 12256 16396 12308 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 5908 16192 5960 16244
rect 7472 16192 7524 16244
rect 8484 16192 8536 16244
rect 10508 16192 10560 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 11704 16235 11756 16244
rect 11704 16201 11713 16235
rect 11713 16201 11747 16235
rect 11747 16201 11756 16235
rect 11704 16192 11756 16201
rect 12256 16192 12308 16244
rect 3424 16056 3476 16108
rect 4804 16056 4856 16108
rect 8024 16056 8076 16108
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 9312 16124 9364 16176
rect 9496 16056 9548 16108
rect 9864 16056 9916 16108
rect 2872 15988 2924 16040
rect 9956 15988 10008 16040
rect 11336 15988 11388 16040
rect 1584 15963 1636 15972
rect 1584 15929 1593 15963
rect 1593 15929 1627 15963
rect 1627 15929 1636 15963
rect 1584 15920 1636 15929
rect 2320 15852 2372 15904
rect 4804 15963 4856 15972
rect 4804 15929 4813 15963
rect 4813 15929 4847 15963
rect 4847 15929 4856 15963
rect 4804 15920 4856 15929
rect 3056 15852 3108 15904
rect 4252 15852 4304 15904
rect 4436 15852 4488 15904
rect 7472 15920 7524 15972
rect 8116 15920 8168 15972
rect 9496 15963 9548 15972
rect 6092 15852 6144 15904
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 9496 15929 9499 15963
rect 9499 15929 9533 15963
rect 9533 15929 9548 15963
rect 9496 15920 9548 15929
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 3424 15648 3476 15700
rect 8852 15691 8904 15700
rect 8852 15657 8861 15691
rect 8861 15657 8895 15691
rect 8895 15657 8904 15691
rect 8852 15648 8904 15657
rect 12072 15648 12124 15700
rect 2320 15580 2372 15632
rect 4252 15580 4304 15632
rect 4988 15580 5040 15632
rect 7472 15580 7524 15632
rect 9128 15623 9180 15632
rect 9128 15589 9137 15623
rect 9137 15589 9171 15623
rect 9171 15589 9180 15623
rect 9128 15580 9180 15589
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 10416 15623 10468 15632
rect 10416 15589 10425 15623
rect 10425 15589 10459 15623
rect 10459 15589 10468 15623
rect 10416 15580 10468 15589
rect 11152 15580 11204 15632
rect 1584 15512 1636 15564
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 2412 15444 2464 15496
rect 2780 15444 2832 15496
rect 5724 15512 5776 15564
rect 6276 15555 6328 15564
rect 6276 15521 6320 15555
rect 6320 15521 6328 15555
rect 11244 15555 11296 15564
rect 6276 15512 6328 15521
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 12624 15512 12676 15564
rect 4896 15376 4948 15428
rect 6920 15376 6972 15428
rect 8208 15444 8260 15496
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10232 15376 10284 15428
rect 3516 15308 3568 15360
rect 4160 15308 4212 15360
rect 4528 15308 4580 15360
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 8668 15308 8720 15360
rect 9404 15308 9456 15360
rect 10784 15308 10836 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 2320 15147 2372 15156
rect 2320 15113 2329 15147
rect 2329 15113 2363 15147
rect 2363 15113 2372 15147
rect 2320 15104 2372 15113
rect 5264 15104 5316 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 8116 15104 8168 15156
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 9864 15147 9916 15156
rect 8668 15104 8720 15113
rect 9864 15113 9873 15147
rect 9873 15113 9907 15147
rect 9907 15113 9916 15147
rect 9864 15104 9916 15113
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 12624 15147 12676 15156
rect 12624 15113 12633 15147
rect 12633 15113 12667 15147
rect 12667 15113 12676 15147
rect 12624 15104 12676 15113
rect 4252 15036 4304 15088
rect 5172 15036 5224 15088
rect 7472 15036 7524 15088
rect 8852 15036 8904 15088
rect 4896 15011 4948 15020
rect 4896 14977 4905 15011
rect 4905 14977 4939 15011
rect 4939 14977 4948 15011
rect 4896 14968 4948 14977
rect 9680 15036 9732 15088
rect 11244 15036 11296 15088
rect 10600 14968 10652 15020
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 1676 14900 1728 14952
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 3424 14943 3476 14952
rect 3424 14909 3433 14943
rect 3433 14909 3467 14943
rect 3467 14909 3476 14943
rect 3424 14900 3476 14909
rect 1860 14832 1912 14884
rect 2504 14832 2556 14884
rect 2964 14832 3016 14884
rect 4160 14900 4212 14952
rect 7196 14900 7248 14952
rect 7472 14900 7524 14952
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 3148 14764 3200 14816
rect 5816 14832 5868 14884
rect 7656 14832 7708 14884
rect 8668 14832 8720 14884
rect 10324 14832 10376 14884
rect 3976 14764 4028 14816
rect 4252 14764 4304 14816
rect 5172 14764 5224 14816
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 10232 14764 10284 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 3516 14560 3568 14612
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 5264 14560 5316 14612
rect 6092 14603 6144 14612
rect 6092 14569 6101 14603
rect 6101 14569 6135 14603
rect 6135 14569 6144 14603
rect 6092 14560 6144 14569
rect 8576 14560 8628 14612
rect 8760 14560 8812 14612
rect 9772 14560 9824 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 10324 14560 10376 14612
rect 4436 14492 4488 14544
rect 5172 14492 5224 14544
rect 5724 14492 5776 14544
rect 8208 14492 8260 14544
rect 2044 14424 2096 14476
rect 2412 14424 2464 14476
rect 3056 14424 3108 14476
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 3976 14424 4028 14476
rect 6828 14424 6880 14476
rect 1860 14356 1912 14408
rect 2688 14356 2740 14408
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 7012 14424 7064 14476
rect 8116 14424 8168 14476
rect 7196 14356 7248 14408
rect 8852 14356 8904 14408
rect 7932 14288 7984 14340
rect 10140 14467 10192 14476
rect 10140 14433 10149 14467
rect 10149 14433 10183 14467
rect 10183 14433 10192 14467
rect 10140 14424 10192 14433
rect 9680 14288 9732 14340
rect 2228 14220 2280 14272
rect 2872 14220 2924 14272
rect 4804 14263 4856 14272
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 7196 14220 7248 14272
rect 8484 14220 8536 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 2688 14059 2740 14068
rect 2688 14025 2697 14059
rect 2697 14025 2731 14059
rect 2731 14025 2740 14059
rect 2688 14016 2740 14025
rect 4436 14016 4488 14068
rect 4988 14016 5040 14068
rect 5356 14016 5408 14068
rect 5448 14016 5500 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 2044 13991 2096 14000
rect 2044 13957 2053 13991
rect 2053 13957 2087 13991
rect 2087 13957 2096 13991
rect 2044 13948 2096 13957
rect 3148 13948 3200 14000
rect 4804 13948 4856 14000
rect 3424 13880 3476 13932
rect 1676 13812 1728 13864
rect 2136 13812 2188 13864
rect 3608 13855 3660 13864
rect 2780 13744 2832 13796
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 5632 13948 5684 14000
rect 7288 13948 7340 14000
rect 5356 13812 5408 13864
rect 7012 13880 7064 13932
rect 7472 14016 7524 14068
rect 7932 14059 7984 14068
rect 7932 14025 7941 14059
rect 7941 14025 7975 14059
rect 7975 14025 7984 14059
rect 7932 14016 7984 14025
rect 8116 14016 8168 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 9772 14016 9824 14068
rect 9496 13880 9548 13932
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 3424 13744 3476 13796
rect 6184 13787 6236 13796
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 3516 13676 3568 13728
rect 3976 13676 4028 13728
rect 6184 13753 6193 13787
rect 6193 13753 6227 13787
rect 6227 13753 6236 13787
rect 6184 13744 6236 13753
rect 4804 13719 4856 13728
rect 4804 13685 4813 13719
rect 4813 13685 4847 13719
rect 4847 13685 4856 13719
rect 4804 13676 4856 13685
rect 5356 13676 5408 13728
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 3056 13472 3108 13524
rect 3240 13472 3292 13524
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 4252 13472 4304 13524
rect 5172 13515 5224 13524
rect 2228 13404 2280 13456
rect 3332 13404 3384 13456
rect 2596 13336 2648 13388
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 6000 13472 6052 13524
rect 7196 13472 7248 13524
rect 7288 13472 7340 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 5080 13404 5132 13456
rect 5448 13404 5500 13456
rect 5908 13404 5960 13456
rect 7932 13404 7984 13456
rect 4804 13336 4856 13388
rect 9588 13336 9640 13388
rect 11980 13336 12032 13388
rect 3424 13268 3476 13320
rect 3608 13268 3660 13320
rect 4712 13268 4764 13320
rect 5356 13311 5408 13320
rect 4988 13200 5040 13252
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 8852 13268 8904 13320
rect 6828 13200 6880 13252
rect 8760 13200 8812 13252
rect 9404 13132 9456 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 4436 12928 4488 12980
rect 2412 12860 2464 12912
rect 4160 12860 4212 12912
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 3148 12588 3200 12640
rect 4436 12792 4488 12844
rect 5356 12928 5408 12980
rect 6920 12928 6972 12980
rect 5172 12860 5224 12912
rect 6736 12860 6788 12912
rect 9588 12860 9640 12912
rect 4896 12724 4948 12776
rect 4528 12656 4580 12708
rect 5724 12792 5776 12844
rect 7840 12792 7892 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9680 12792 9732 12844
rect 6184 12724 6236 12776
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 10324 12724 10376 12776
rect 11520 12928 11572 12980
rect 5908 12588 5960 12640
rect 6000 12588 6052 12640
rect 7288 12588 7340 12640
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 8024 12588 8076 12640
rect 9772 12588 9824 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 4528 12384 4580 12436
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 8852 12427 8904 12436
rect 8852 12393 8861 12427
rect 8861 12393 8895 12427
rect 8895 12393 8904 12427
rect 8852 12384 8904 12393
rect 5908 12316 5960 12368
rect 7012 12316 7064 12368
rect 9772 12359 9824 12368
rect 9772 12325 9781 12359
rect 9781 12325 9815 12359
rect 9815 12325 9824 12359
rect 9772 12316 9824 12325
rect 9864 12359 9916 12368
rect 9864 12325 9873 12359
rect 9873 12325 9907 12359
rect 9907 12325 9916 12359
rect 9864 12316 9916 12325
rect 2412 12248 2464 12300
rect 2872 12248 2924 12300
rect 4712 12248 4764 12300
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 5632 12248 5684 12257
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 11428 12248 11480 12300
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 1676 12112 1728 12164
rect 5632 12112 5684 12164
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 7932 12155 7984 12164
rect 7932 12121 7941 12155
rect 7941 12121 7975 12155
rect 7975 12121 7984 12155
rect 7932 12112 7984 12121
rect 9864 12112 9916 12164
rect 3056 12044 3108 12096
rect 4712 12044 4764 12096
rect 6460 12087 6512 12096
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 10600 12044 10652 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2412 11883 2464 11892
rect 2412 11849 2421 11883
rect 2421 11849 2455 11883
rect 2455 11849 2464 11883
rect 2412 11840 2464 11849
rect 3424 11883 3476 11892
rect 3424 11849 3433 11883
rect 3433 11849 3467 11883
rect 3467 11849 3476 11883
rect 3424 11840 3476 11849
rect 4068 11840 4120 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5080 11704 5132 11756
rect 6000 11840 6052 11892
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 6460 11704 6512 11756
rect 8944 11704 8996 11756
rect 6184 11636 6236 11688
rect 6920 11568 6972 11620
rect 2964 11500 3016 11552
rect 3424 11500 3476 11552
rect 4160 11543 4212 11552
rect 4160 11509 4169 11543
rect 4169 11509 4203 11543
rect 4203 11509 4212 11543
rect 4160 11500 4212 11509
rect 7012 11500 7064 11552
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8760 11500 8812 11552
rect 8944 11611 8996 11620
rect 8944 11577 8953 11611
rect 8953 11577 8987 11611
rect 8987 11577 8996 11611
rect 8944 11568 8996 11577
rect 10232 11568 10284 11620
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 11520 11568 11572 11620
rect 11428 11543 11480 11552
rect 10140 11500 10192 11509
rect 11428 11509 11437 11543
rect 11437 11509 11471 11543
rect 11471 11509 11480 11543
rect 11428 11500 11480 11509
rect 12624 11500 12676 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 3516 11296 3568 11348
rect 5080 11296 5132 11348
rect 5632 11339 5684 11348
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 8944 11296 8996 11348
rect 9772 11296 9824 11348
rect 3148 11271 3200 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2780 11160 2832 11212
rect 3148 11237 3157 11271
rect 3157 11237 3191 11271
rect 3191 11237 3200 11271
rect 3148 11228 3200 11237
rect 7012 11228 7064 11280
rect 7932 11228 7984 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 11428 11271 11480 11280
rect 11428 11237 11437 11271
rect 11437 11237 11471 11271
rect 11471 11237 11480 11271
rect 11428 11228 11480 11237
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 4160 11203 4212 11212
rect 4160 11169 4169 11203
rect 4169 11169 4203 11203
rect 4203 11169 4212 11203
rect 4344 11203 4396 11212
rect 4160 11160 4212 11169
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 6000 11160 6052 11212
rect 2964 11092 3016 11144
rect 7196 11092 7248 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 10232 11135 10284 11144
rect 2504 11067 2556 11076
rect 2504 11033 2513 11067
rect 2513 11033 2547 11067
rect 2547 11033 2556 11067
rect 2504 11024 2556 11033
rect 3056 11024 3108 11076
rect 7104 11024 7156 11076
rect 7656 11024 7708 11076
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10600 11024 10652 11076
rect 4252 10956 4304 11008
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 9680 10956 9732 11008
rect 11520 11092 11572 11144
rect 11612 10956 11664 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 4988 10795 5040 10804
rect 4988 10761 4997 10795
rect 4997 10761 5031 10795
rect 5031 10761 5040 10795
rect 4988 10752 5040 10761
rect 6000 10752 6052 10804
rect 7288 10752 7340 10804
rect 8852 10752 8904 10804
rect 9864 10752 9916 10804
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 11612 10795 11664 10804
rect 11612 10761 11621 10795
rect 11621 10761 11655 10795
rect 11655 10761 11664 10795
rect 11612 10752 11664 10761
rect 3056 10684 3108 10736
rect 3976 10684 4028 10736
rect 10140 10684 10192 10736
rect 2504 10616 2556 10668
rect 4252 10616 4304 10668
rect 8208 10616 8260 10668
rect 11428 10616 11480 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 2780 10523 2832 10532
rect 2780 10489 2789 10523
rect 2789 10489 2823 10523
rect 2823 10489 2832 10523
rect 2780 10480 2832 10489
rect 3976 10548 4028 10600
rect 4344 10548 4396 10600
rect 5540 10548 5592 10600
rect 6000 10548 6052 10600
rect 7104 10548 7156 10600
rect 5908 10523 5960 10532
rect 5908 10489 5917 10523
rect 5917 10489 5951 10523
rect 5951 10489 5960 10523
rect 5908 10480 5960 10489
rect 7012 10480 7064 10532
rect 8116 10480 8168 10532
rect 9220 10523 9272 10532
rect 9220 10489 9229 10523
rect 9229 10489 9263 10523
rect 9263 10489 9272 10523
rect 9220 10480 9272 10489
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 8852 10412 8904 10464
rect 9680 10480 9732 10532
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 2412 10208 2464 10260
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 5540 10208 5592 10260
rect 5724 10208 5776 10260
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 9220 10251 9272 10260
rect 9220 10217 9229 10251
rect 9229 10217 9263 10251
rect 9263 10217 9272 10251
rect 9220 10208 9272 10217
rect 1400 10140 1452 10192
rect 4068 10140 4120 10192
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 8116 10140 8168 10192
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 4252 10115 4304 10124
rect 2688 10072 2740 10081
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 4436 10072 4488 10124
rect 5172 10072 5224 10124
rect 6000 10072 6052 10124
rect 7196 10072 7248 10124
rect 3976 10004 4028 10056
rect 4160 10004 4212 10056
rect 5356 10004 5408 10056
rect 6920 10004 6972 10056
rect 9588 10004 9640 10056
rect 3148 9936 3200 9988
rect 5448 9936 5500 9988
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 2412 9664 2464 9716
rect 2504 9664 2556 9716
rect 3148 9707 3200 9716
rect 3148 9673 3157 9707
rect 3157 9673 3191 9707
rect 3191 9673 3200 9707
rect 3148 9664 3200 9673
rect 3976 9664 4028 9716
rect 4252 9664 4304 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 6000 9707 6052 9716
rect 6000 9673 6009 9707
rect 6009 9673 6043 9707
rect 6043 9673 6052 9707
rect 6000 9664 6052 9673
rect 7196 9664 7248 9716
rect 8760 9664 8812 9716
rect 9588 9707 9640 9716
rect 9588 9673 9597 9707
rect 9597 9673 9631 9707
rect 9631 9673 9640 9707
rect 9588 9664 9640 9673
rect 10324 9707 10376 9716
rect 10324 9673 10333 9707
rect 10333 9673 10367 9707
rect 10367 9673 10376 9707
rect 10324 9664 10376 9673
rect 10968 9664 11020 9716
rect 4068 9639 4120 9648
rect 4068 9605 4077 9639
rect 4077 9605 4111 9639
rect 4111 9605 4120 9639
rect 4068 9596 4120 9605
rect 8300 9596 8352 9648
rect 2688 9528 2740 9580
rect 3240 9528 3292 9580
rect 4436 9528 4488 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5264 9528 5316 9580
rect 2964 9503 3016 9512
rect 2964 9469 2973 9503
rect 2973 9469 3007 9503
rect 3007 9469 3016 9503
rect 2964 9460 3016 9469
rect 3516 9324 3568 9376
rect 4344 9460 4396 9512
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 7196 9528 7248 9580
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 7748 9435 7800 9444
rect 7748 9401 7757 9435
rect 7757 9401 7791 9435
rect 7791 9401 7800 9435
rect 7748 9392 7800 9401
rect 10324 9460 10376 9512
rect 10968 9460 11020 9512
rect 9496 9392 9548 9444
rect 10692 9392 10744 9444
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 9680 9324 9732 9376
rect 10508 9324 10560 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 9588 9120 9640 9172
rect 2780 9052 2832 9104
rect 4804 9095 4856 9104
rect 3516 8984 3568 9036
rect 3976 8848 4028 8900
rect 4252 8984 4304 9036
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 6644 9052 6696 9104
rect 10232 9052 10284 9104
rect 4988 8984 5040 9036
rect 11244 9027 11296 9036
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 6736 8916 6788 8968
rect 3332 8780 3384 8832
rect 7840 8848 7892 8900
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 7564 8780 7616 8832
rect 11244 8993 11288 9027
rect 11288 8993 11296 9027
rect 11244 8984 11296 8993
rect 11428 8984 11480 9036
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 10416 8848 10468 8900
rect 10600 8780 10652 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 2872 8576 2924 8628
rect 3516 8576 3568 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 11428 8576 11480 8628
rect 3056 8508 3108 8560
rect 4068 8508 4120 8560
rect 5816 8551 5868 8560
rect 5816 8517 5825 8551
rect 5825 8517 5859 8551
rect 5859 8517 5868 8551
rect 5816 8508 5868 8517
rect 112 8440 164 8492
rect 3332 8440 3384 8492
rect 7288 8440 7340 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9680 8440 9732 8492
rect 4620 8372 4672 8424
rect 10784 8415 10836 8424
rect 10784 8381 10802 8415
rect 10802 8381 10836 8415
rect 10784 8372 10836 8381
rect 3792 8304 3844 8356
rect 9036 8347 9088 8356
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 9864 8347 9916 8356
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 6644 8236 6696 8245
rect 7104 8236 7156 8288
rect 7472 8236 7524 8288
rect 10232 8279 10284 8288
rect 10232 8245 10241 8279
rect 10241 8245 10275 8279
rect 10275 8245 10284 8279
rect 10232 8236 10284 8245
rect 10600 8236 10652 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 3332 8032 3384 8084
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 6000 8032 6052 8084
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 8116 8032 8168 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 4620 8007 4672 8016
rect 4620 7973 4629 8007
rect 4629 7973 4663 8007
rect 4663 7973 4672 8007
rect 4620 7964 4672 7973
rect 5448 7964 5500 8016
rect 9036 7964 9088 8016
rect 9588 7964 9640 8016
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 2136 7896 2188 7948
rect 2964 7939 3016 7948
rect 2964 7905 3008 7939
rect 3008 7905 3016 7939
rect 2964 7896 3016 7905
rect 4436 7896 4488 7948
rect 6828 7939 6880 7948
rect 6828 7905 6837 7939
rect 6837 7905 6871 7939
rect 6871 7905 6880 7939
rect 6828 7896 6880 7905
rect 7748 7896 7800 7948
rect 11520 7896 11572 7948
rect 12072 7896 12124 7948
rect 5172 7828 5224 7880
rect 9496 7828 9548 7880
rect 10508 7828 10560 7880
rect 10232 7760 10284 7812
rect 4068 7692 4120 7744
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 6184 7692 6236 7744
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 6552 7692 6604 7744
rect 7472 7692 7524 7744
rect 10692 7692 10744 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 6276 7488 6328 7540
rect 9588 7488 9640 7540
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 2596 7420 2648 7472
rect 6828 7420 6880 7472
rect 9864 7420 9916 7472
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5908 7352 5960 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 8208 7352 8260 7404
rect 9036 7352 9088 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4068 7284 4120 7336
rect 4896 7284 4948 7336
rect 2964 7216 3016 7268
rect 8668 7284 8720 7336
rect 5448 7148 5500 7200
rect 7932 7191 7984 7200
rect 7932 7157 7941 7191
rect 7941 7157 7975 7191
rect 7975 7157 7984 7191
rect 7932 7148 7984 7157
rect 8116 7148 8168 7200
rect 10232 7216 10284 7268
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 3424 6987 3476 6996
rect 3424 6953 3433 6987
rect 3433 6953 3467 6987
rect 3467 6953 3476 6987
rect 3424 6944 3476 6953
rect 4068 6808 4120 6860
rect 5264 6944 5316 6996
rect 7012 6987 7064 6996
rect 7012 6953 7021 6987
rect 7021 6953 7055 6987
rect 7055 6953 7064 6987
rect 7012 6944 7064 6953
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 8116 6944 8168 6996
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 10600 6944 10652 6996
rect 5172 6919 5224 6928
rect 5172 6885 5181 6919
rect 5181 6885 5215 6919
rect 5215 6885 5224 6919
rect 5172 6876 5224 6885
rect 6184 6919 6236 6928
rect 6184 6885 6193 6919
rect 6193 6885 6227 6919
rect 6227 6885 6236 6919
rect 6184 6876 6236 6885
rect 6736 6919 6788 6928
rect 6736 6885 6745 6919
rect 6745 6885 6779 6919
rect 6779 6885 6788 6919
rect 6736 6876 6788 6885
rect 9312 6876 9364 6928
rect 10416 6919 10468 6928
rect 10416 6885 10425 6919
rect 10425 6885 10459 6919
rect 10459 6885 10468 6919
rect 10416 6876 10468 6885
rect 4896 6851 4948 6860
rect 4896 6817 4905 6851
rect 4905 6817 4939 6851
rect 4939 6817 4948 6851
rect 4896 6808 4948 6817
rect 12624 6808 12676 6860
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 10692 6740 10744 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 3056 6672 3108 6724
rect 7748 6672 7800 6724
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9496 6604 9548 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 1860 6400 1912 6452
rect 4068 6375 4120 6384
rect 4068 6341 4077 6375
rect 4077 6341 4111 6375
rect 4111 6341 4120 6375
rect 4068 6332 4120 6341
rect 6092 6400 6144 6452
rect 7656 6400 7708 6452
rect 8300 6400 8352 6452
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 10692 6400 10744 6452
rect 11428 6400 11480 6452
rect 6184 6332 6236 6384
rect 15108 6332 15160 6384
rect 4896 6196 4948 6248
rect 7840 6264 7892 6316
rect 9496 6264 9548 6316
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 10508 6196 10560 6248
rect 112 6128 164 6180
rect 2044 6128 2096 6180
rect 7012 6128 7064 6180
rect 9312 6171 9364 6180
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9864 6171 9916 6180
rect 9312 6128 9364 6137
rect 9864 6137 9873 6171
rect 9873 6137 9907 6171
rect 9907 6137 9916 6171
rect 9864 6128 9916 6137
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 8116 6060 8168 6112
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 6092 5856 6144 5908
rect 9496 5856 9548 5908
rect 7932 5788 7984 5840
rect 10048 5788 10100 5840
rect 10508 5788 10560 5840
rect 5632 5720 5684 5772
rect 7196 5720 7248 5772
rect 7472 5720 7524 5772
rect 8484 5720 8536 5772
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 11244 5652 11296 5704
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4620 5312 4672 5364
rect 5632 5312 5684 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 5908 5244 5960 5296
rect 6736 5176 6788 5228
rect 4712 5108 4764 5160
rect 8484 5108 8536 5160
rect 10232 5108 10284 5160
rect 5448 5040 5500 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 6092 4972 6144 5024
rect 6828 4972 6880 5024
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 5356 4768 5408 4820
rect 5816 4768 5868 4820
rect 6092 4743 6144 4752
rect 6092 4709 6101 4743
rect 6101 4709 6135 4743
rect 6135 4709 6144 4743
rect 6092 4700 6144 4709
rect 6736 4768 6788 4820
rect 7196 4768 7248 4820
rect 8208 4768 8260 4820
rect 10416 4768 10468 4820
rect 7656 4743 7708 4752
rect 7656 4709 7665 4743
rect 7665 4709 7699 4743
rect 7699 4709 7708 4743
rect 7656 4700 7708 4709
rect 4712 4632 4764 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 10968 4632 11020 4684
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 7288 4564 7340 4616
rect 4988 4496 5040 4548
rect 5816 4496 5868 4548
rect 4160 4428 4212 4480
rect 8392 4428 8444 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 3424 4224 3476 4276
rect 4160 4224 4212 4276
rect 6000 4224 6052 4276
rect 8300 4224 8352 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 4896 4156 4948 4208
rect 4988 4199 5040 4208
rect 4988 4165 4997 4199
rect 4997 4165 5031 4199
rect 5031 4165 5040 4199
rect 4988 4156 5040 4165
rect 6092 4156 6144 4208
rect 7656 4156 7708 4208
rect 7288 4088 7340 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 10416 4224 10468 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 5448 3952 5500 4004
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 7380 3952 7432 4004
rect 10140 3995 10192 4004
rect 6644 3884 6696 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 10140 3961 10149 3995
rect 10149 3961 10183 3995
rect 10183 3961 10192 3995
rect 10140 3952 10192 3961
rect 9128 3927 9180 3936
rect 8116 3884 8168 3893
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 5080 3680 5132 3732
rect 6184 3680 6236 3732
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 4896 3587 4948 3596
rect 4528 3476 4580 3528
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 8484 3680 8536 3732
rect 10140 3680 10192 3732
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 9128 3612 9180 3664
rect 9496 3612 9548 3664
rect 6552 3476 6604 3528
rect 8024 3476 8076 3528
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10048 3476 10100 3528
rect 8300 3408 8352 3460
rect 10324 3451 10376 3460
rect 10324 3417 10333 3451
rect 10333 3417 10367 3451
rect 10367 3417 10376 3451
rect 10324 3408 10376 3417
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 5540 3340 5592 3392
rect 12624 3340 12676 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 112 3136 164 3188
rect 3976 3136 4028 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 5448 3136 5500 3188
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 9496 3179 9548 3188
rect 9496 3145 9505 3179
rect 9505 3145 9539 3179
rect 9539 3145 9548 3179
rect 9496 3136 9548 3145
rect 9772 3136 9824 3188
rect 4896 3000 4948 3052
rect 5080 3000 5132 3052
rect 5724 3068 5776 3120
rect 7196 3000 7248 3052
rect 8024 3000 8076 3052
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 6736 2932 6788 2984
rect 6920 2932 6972 2984
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 10784 2932 10836 2984
rect 6184 2907 6236 2916
rect 1768 2796 1820 2848
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 6184 2873 6193 2907
rect 6193 2873 6227 2907
rect 6227 2873 6236 2907
rect 6184 2864 6236 2873
rect 8024 2839 8076 2848
rect 4804 2796 4856 2805
rect 8024 2805 8033 2839
rect 8033 2805 8067 2839
rect 8067 2805 8076 2839
rect 8024 2796 8076 2805
rect 10324 2864 10376 2916
rect 11060 2864 11112 2916
rect 12348 2796 12400 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 3976 2592 4028 2644
rect 4896 2592 4948 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 6644 2524 6696 2576
rect 7196 2567 7248 2576
rect 7196 2533 7205 2567
rect 7205 2533 7239 2567
rect 7239 2533 7248 2567
rect 7196 2524 7248 2533
rect 6736 2456 6788 2508
rect 8852 2456 8904 2508
rect 7012 2388 7064 2440
rect 11060 2456 11112 2508
rect 5540 2320 5592 2372
rect 5908 2363 5960 2372
rect 5908 2329 5917 2363
rect 5917 2329 5951 2363
rect 5951 2329 5960 2363
rect 5908 2320 5960 2329
rect 10784 2320 10836 2372
rect 13360 2320 13412 2372
rect 4528 2252 4580 2304
rect 6184 2252 6236 2304
rect 7196 2252 7248 2304
rect 8024 2252 8076 2304
rect 9772 2252 9824 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 11060 2252 11112 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
<< metal2 >>
rect 570 39636 626 40000
rect 1674 39658 1730 40000
rect 570 39584 572 39636
rect 624 39584 626 39636
rect 570 39520 626 39584
rect 1216 39636 1268 39642
rect 1216 39578 1268 39584
rect 1674 39630 1808 39658
rect 112 21956 164 21962
rect 112 21898 164 21904
rect 124 18601 152 21898
rect 1228 21486 1256 39578
rect 1674 39520 1730 39630
rect 1674 38040 1730 38049
rect 1674 37975 1730 37984
rect 1582 29472 1638 29481
rect 1582 29407 1638 29416
rect 1596 28762 1624 29407
rect 1584 28756 1636 28762
rect 1584 28698 1636 28704
rect 1400 28620 1452 28626
rect 1400 28562 1452 28568
rect 1412 28014 1440 28562
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1582 24032 1638 24041
rect 1582 23967 1638 23976
rect 1596 23322 1624 23967
rect 1688 23866 1716 37975
rect 1780 25906 1808 39630
rect 2778 39636 2834 40000
rect 3974 39658 4030 40000
rect 5078 39658 5134 40000
rect 6274 39658 6330 40000
rect 7378 39658 7434 40000
rect 2778 39584 2780 39636
rect 2832 39584 2834 39636
rect 2778 39520 2834 39584
rect 3516 39636 3568 39642
rect 3516 39578 3568 39584
rect 3974 39630 4200 39658
rect 2502 35184 2558 35193
rect 2502 35119 2558 35128
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 2056 25974 2084 26386
rect 2044 25968 2096 25974
rect 2044 25910 2096 25916
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 2412 25832 2464 25838
rect 2412 25774 2464 25780
rect 2424 25226 2452 25774
rect 2412 25220 2464 25226
rect 2412 25162 2464 25168
rect 2228 24676 2280 24682
rect 2228 24618 2280 24624
rect 2240 24274 2268 24618
rect 2516 24410 2544 35119
rect 3424 32020 3476 32026
rect 3424 31962 3476 31968
rect 2688 28620 2740 28626
rect 2688 28562 2740 28568
rect 2596 27940 2648 27946
rect 2596 27882 2648 27888
rect 2504 24404 2556 24410
rect 2504 24346 2556 24352
rect 2228 24268 2280 24274
rect 2228 24210 2280 24216
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1780 23662 1808 24006
rect 1768 23656 1820 23662
rect 1768 23598 1820 23604
rect 2056 23526 2084 24142
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1676 23248 1728 23254
rect 1676 23190 1728 23196
rect 1688 22778 1716 23190
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 2056 22001 2084 23462
rect 2412 22024 2464 22030
rect 2042 21992 2098 22001
rect 2412 21966 2464 21972
rect 2042 21927 2098 21936
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 1216 21480 1268 21486
rect 1216 21422 1268 21428
rect 1412 21010 1440 21830
rect 2056 21554 2084 21927
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 1860 21480 1912 21486
rect 1860 21422 1912 21428
rect 1872 21146 1900 21422
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 2240 21146 2268 21354
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 2228 21140 2280 21146
rect 2228 21082 2280 21088
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 18970 1440 20946
rect 1872 20505 1900 21082
rect 2228 20868 2280 20874
rect 2228 20810 2280 20816
rect 1858 20496 1914 20505
rect 1584 20460 1636 20466
rect 1858 20431 1914 20440
rect 1584 20402 1636 20408
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1504 18630 1532 19246
rect 1596 18834 1624 20402
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1688 19990 1716 20334
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1780 19242 1808 19654
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1674 18864 1730 18873
rect 1584 18828 1636 18834
rect 1674 18799 1730 18808
rect 1584 18770 1636 18776
rect 664 18624 716 18630
rect 110 18592 166 18601
rect 664 18566 716 18572
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 110 18527 166 18536
rect 124 8498 152 18527
rect 112 8492 164 8498
rect 112 8434 164 8440
rect 110 7168 166 7177
rect 110 7103 166 7112
rect 124 6186 152 7103
rect 112 6180 164 6186
rect 112 6122 164 6128
rect 112 3188 164 3194
rect 112 3130 164 3136
rect 124 1465 152 3130
rect 110 1456 166 1465
rect 110 1391 166 1400
rect 478 82 534 480
rect 676 82 704 18566
rect 1596 17882 1624 18770
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1400 17060 1452 17066
rect 1400 17002 1452 17008
rect 1412 16794 1440 17002
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 15978 1624 16390
rect 1584 15972 1636 15978
rect 1584 15914 1636 15920
rect 1596 15570 1624 15914
rect 1688 15706 1716 18799
rect 1872 18408 1900 20431
rect 1950 20360 2006 20369
rect 1950 20295 2006 20304
rect 2136 20324 2188 20330
rect 1964 20058 1992 20295
rect 2136 20266 2188 20272
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1952 18420 2004 18426
rect 1872 18380 1952 18408
rect 1952 18362 2004 18368
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17882 1992 18158
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1582 15192 1638 15201
rect 1582 15127 1638 15136
rect 1596 14074 1624 15127
rect 1688 14958 1716 15642
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1780 13814 1808 17750
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1872 14414 1900 14826
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1964 13814 1992 17818
rect 2148 17270 2176 20266
rect 2240 20262 2268 20810
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 2240 19854 2268 20198
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2332 19334 2360 21830
rect 2424 21010 2452 21966
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2424 19417 2452 20946
rect 2410 19408 2466 19417
rect 2410 19343 2466 19352
rect 2240 19306 2360 19334
rect 2240 17814 2268 19306
rect 2320 19236 2372 19242
rect 2320 19178 2372 19184
rect 2332 18766 2360 19178
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2148 15706 2176 16526
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2240 15586 2268 17478
rect 2332 17338 2360 17614
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2332 16998 2360 17274
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 15638 2360 15846
rect 2148 15558 2268 15586
rect 2320 15632 2372 15638
rect 2320 15574 2372 15580
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2056 14006 2084 14418
rect 2044 14000 2096 14006
rect 2044 13942 2096 13948
rect 2148 13870 2176 15558
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2240 14278 2268 15438
rect 2332 15162 2360 15574
rect 2424 15502 2452 19343
rect 2516 18986 2544 23598
rect 2608 20210 2636 27882
rect 2700 27402 2728 28562
rect 2688 27396 2740 27402
rect 2688 27338 2740 27344
rect 2700 20330 2728 27338
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 2884 23866 2912 24210
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2792 20584 2820 22374
rect 2884 21593 2912 23802
rect 2976 23474 3004 25842
rect 3068 25702 3096 26386
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3068 24177 3096 25638
rect 3054 24168 3110 24177
rect 3054 24103 3110 24112
rect 3056 23520 3108 23526
rect 2976 23468 3056 23474
rect 2976 23462 3108 23468
rect 2976 23446 3096 23462
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2976 22642 3004 22918
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 2976 22438 3004 22578
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2870 21584 2926 21593
rect 2870 21519 2926 21528
rect 2976 21350 3004 22374
rect 3068 22098 3096 23446
rect 3160 23186 3188 27066
rect 3436 27062 3464 31962
rect 3424 27056 3476 27062
rect 3424 26998 3476 27004
rect 3436 26586 3464 26998
rect 3424 26580 3476 26586
rect 3424 26522 3476 26528
rect 3332 26240 3384 26246
rect 3332 26182 3384 26188
rect 3344 25906 3372 26182
rect 3332 25900 3384 25906
rect 3332 25842 3384 25848
rect 3240 25356 3292 25362
rect 3240 25298 3292 25304
rect 3252 24614 3280 25298
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3148 23180 3200 23186
rect 3148 23122 3200 23128
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3068 21690 3096 22034
rect 3160 21962 3188 23122
rect 3148 21956 3200 21962
rect 3148 21898 3200 21904
rect 3056 21684 3108 21690
rect 3108 21644 3188 21672
rect 3056 21626 3108 21632
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2792 20556 2912 20584
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2608 20182 2820 20210
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 19446 2636 19858
rect 2596 19440 2648 19446
rect 2648 19400 2728 19428
rect 2596 19382 2648 19388
rect 2516 18958 2636 18986
rect 2608 17202 2636 18958
rect 2700 18426 2728 19400
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2792 18222 2820 20182
rect 2884 19394 2912 20556
rect 2976 20398 3004 21286
rect 3068 21010 3096 21422
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 3068 19446 3096 20946
rect 3160 20602 3188 21644
rect 3252 21078 3280 24550
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 3436 23662 3464 24006
rect 3528 23798 3556 39578
rect 3974 39520 4030 39630
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 4068 33584 4120 33590
rect 4068 33526 4120 33532
rect 3976 33380 4028 33386
rect 3976 33322 4028 33328
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3988 31278 4016 33322
rect 4080 32366 4108 33526
rect 4172 33134 4200 39630
rect 5078 39630 5396 39658
rect 5078 39520 5134 39630
rect 5368 35562 5396 39630
rect 6196 39630 6330 39658
rect 5540 35624 5592 35630
rect 5540 35566 5592 35572
rect 5356 35556 5408 35562
rect 5356 35498 5408 35504
rect 5552 34746 5580 35566
rect 6196 35154 6224 39630
rect 6274 39520 6330 39630
rect 7116 39630 7434 39658
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6736 35556 6788 35562
rect 6736 35498 6788 35504
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6184 35148 6236 35154
rect 6184 35090 6236 35096
rect 6196 34746 6224 35090
rect 6748 34746 6776 35498
rect 6828 35488 6880 35494
rect 6828 35430 6880 35436
rect 6840 35290 6868 35430
rect 6828 35284 6880 35290
rect 6828 35226 6880 35232
rect 5540 34740 5592 34746
rect 5540 34682 5592 34688
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 6184 34740 6236 34746
rect 6184 34682 6236 34688
rect 6736 34740 6788 34746
rect 6736 34682 6788 34688
rect 5552 34542 5580 34682
rect 5540 34536 5592 34542
rect 5540 34478 5592 34484
rect 4804 33992 4856 33998
rect 4804 33934 4856 33940
rect 4620 33380 4672 33386
rect 4620 33322 4672 33328
rect 4172 33106 4568 33134
rect 4632 33114 4660 33322
rect 4712 33312 4764 33318
rect 4712 33254 4764 33260
rect 4344 32836 4396 32842
rect 4344 32778 4396 32784
rect 4160 32496 4212 32502
rect 4160 32438 4212 32444
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 4080 32026 4108 32302
rect 4068 32020 4120 32026
rect 4068 31962 4120 31968
rect 3976 31272 4028 31278
rect 3976 31214 4028 31220
rect 3988 30938 4016 31214
rect 3976 30932 4028 30938
rect 4028 30892 4108 30920
rect 3976 30874 4028 30880
rect 3976 30796 4028 30802
rect 3976 30738 4028 30744
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3988 30394 4016 30738
rect 4080 30394 4108 30892
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4172 30274 4200 32438
rect 4356 32434 4384 32778
rect 4344 32428 4396 32434
rect 4344 32370 4396 32376
rect 4250 32328 4306 32337
rect 4250 32263 4306 32272
rect 4344 32292 4396 32298
rect 4264 30870 4292 32263
rect 4344 32234 4396 32240
rect 4252 30864 4304 30870
rect 4252 30806 4304 30812
rect 4080 30246 4200 30274
rect 4080 29714 4108 30246
rect 4356 30190 4384 32234
rect 4344 30184 4396 30190
rect 4344 30126 4396 30132
rect 4436 30116 4488 30122
rect 4436 30058 4488 30064
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3884 28960 3936 28966
rect 4080 28948 4108 29650
rect 4172 29170 4200 29786
rect 4448 29714 4476 30058
rect 4436 29708 4488 29714
rect 4540 29696 4568 33106
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 4724 32892 4752 33254
rect 4816 32994 4844 33934
rect 4988 33380 5040 33386
rect 4988 33322 5040 33328
rect 5000 33046 5028 33322
rect 4988 33040 5040 33046
rect 4816 32966 4936 32994
rect 4988 32982 5040 32988
rect 4804 32904 4856 32910
rect 4724 32864 4804 32892
rect 4804 32846 4856 32852
rect 4816 32026 4844 32846
rect 4908 32434 4936 32966
rect 4896 32428 4948 32434
rect 4896 32370 4948 32376
rect 5000 32230 5028 32982
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5368 32298 5396 32710
rect 5356 32292 5408 32298
rect 5356 32234 5408 32240
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 4804 32020 4856 32026
rect 4804 31962 4856 31968
rect 5000 31958 5028 32166
rect 4988 31952 5040 31958
rect 4988 31894 5040 31900
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4632 31142 4660 31758
rect 5000 31346 5028 31894
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 5000 31210 5028 31282
rect 4988 31204 5040 31210
rect 4988 31146 5040 31152
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4632 30054 4660 31078
rect 5000 30598 5028 31146
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 4988 30592 5040 30598
rect 4988 30534 5040 30540
rect 5000 30326 5028 30534
rect 4988 30320 5040 30326
rect 4988 30262 5040 30268
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4620 29708 4672 29714
rect 4540 29668 4620 29696
rect 4436 29650 4488 29656
rect 4620 29650 4672 29656
rect 4160 29164 4212 29170
rect 4160 29106 4212 29112
rect 3936 28920 4108 28948
rect 3884 28902 3936 28908
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3700 27872 3752 27878
rect 3700 27814 3752 27820
rect 3712 27402 3740 27814
rect 3988 27674 4016 28358
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 3700 27396 3752 27402
rect 3700 27338 3752 27344
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3988 26926 4016 27610
rect 4080 27606 4108 28920
rect 4448 28762 4476 29650
rect 5000 29034 5028 30262
rect 5368 30054 5396 30670
rect 5356 30048 5408 30054
rect 5356 29990 5408 29996
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 5000 28762 5028 28970
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4436 28756 4488 28762
rect 4436 28698 4488 28704
rect 4988 28756 5040 28762
rect 4988 28698 5040 28704
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 4252 27872 4304 27878
rect 4252 27814 4304 27820
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4264 26994 4292 27814
rect 4356 27674 4384 28494
rect 4448 28422 4476 28698
rect 5092 28694 5120 28902
rect 5080 28688 5132 28694
rect 5080 28630 5132 28636
rect 4436 28416 4488 28422
rect 4436 28358 4488 28364
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4620 28144 4672 28150
rect 4620 28086 4672 28092
rect 4344 27668 4396 27674
rect 4344 27610 4396 27616
rect 4436 27396 4488 27402
rect 4436 27338 4488 27344
rect 4448 27130 4476 27338
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 4252 26988 4304 26994
rect 4252 26930 4304 26936
rect 3976 26920 4028 26926
rect 4028 26880 4108 26908
rect 3976 26862 4028 26868
rect 3976 26580 4028 26586
rect 3976 26522 4028 26528
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3988 25956 4016 26522
rect 3896 25928 4016 25956
rect 3896 25838 3924 25928
rect 3884 25832 3936 25838
rect 3884 25774 3936 25780
rect 3896 25498 3924 25774
rect 3976 25764 4028 25770
rect 3976 25706 4028 25712
rect 3884 25492 3936 25498
rect 3884 25434 3936 25440
rect 3988 25294 4016 25706
rect 3976 25288 4028 25294
rect 3976 25230 4028 25236
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3896 24614 3924 24686
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 24154 3924 24550
rect 3988 24274 4016 25230
rect 4080 24886 4108 26880
rect 4344 26852 4396 26858
rect 4344 26794 4396 26800
rect 4158 26616 4214 26625
rect 4158 26551 4214 26560
rect 4252 26580 4304 26586
rect 4172 24954 4200 26551
rect 4252 26522 4304 26528
rect 4264 25702 4292 26522
rect 4356 26382 4384 26794
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4344 26376 4396 26382
rect 4344 26318 4396 26324
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4356 25498 4384 26318
rect 4540 26042 4568 26454
rect 4632 26042 4660 28086
rect 5000 28082 5028 28358
rect 5092 28218 5120 28630
rect 5368 28558 5396 29990
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5080 28212 5132 28218
rect 5080 28154 5132 28160
rect 4988 28076 5040 28082
rect 4988 28018 5040 28024
rect 5092 27946 5120 28154
rect 5080 27940 5132 27946
rect 5080 27882 5132 27888
rect 5092 27674 5120 27882
rect 5080 27668 5132 27674
rect 5080 27610 5132 27616
rect 4988 27600 5040 27606
rect 4988 27542 5040 27548
rect 4804 27532 4856 27538
rect 4804 27474 4856 27480
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4344 25492 4396 25498
rect 4344 25434 4396 25440
rect 4540 25430 4568 25978
rect 4724 25838 4752 27406
rect 4816 27062 4844 27474
rect 4804 27056 4856 27062
rect 4804 26998 4856 27004
rect 4816 26790 4844 26998
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4528 25424 4580 25430
rect 4528 25366 4580 25372
rect 4540 24954 4568 25366
rect 4724 25294 4752 25638
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4436 24880 4488 24886
rect 4436 24822 4488 24828
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 3976 24268 4028 24274
rect 3976 24210 4028 24216
rect 3896 24126 4016 24154
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3516 23792 3568 23798
rect 3516 23734 3568 23740
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3344 22166 3372 22510
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 3344 21486 3372 22102
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3344 21146 3372 21422
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3240 21072 3292 21078
rect 3240 21014 3292 21020
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3436 20448 3464 23462
rect 3528 22982 3556 23734
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3988 22642 4016 24126
rect 4080 22778 4108 24686
rect 4448 24206 4476 24822
rect 4436 24200 4488 24206
rect 4436 24142 4488 24148
rect 4252 23588 4304 23594
rect 4252 23530 4304 23536
rect 4264 22964 4292 23530
rect 4448 23322 4476 24142
rect 4540 24138 4568 24890
rect 4632 24410 4660 25230
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4540 23730 4568 24074
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 4724 23526 4752 24210
rect 4816 23866 4844 26726
rect 4896 25220 4948 25226
rect 4896 25162 4948 25168
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4724 23186 4752 23462
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4344 22976 4396 22982
rect 4264 22936 4344 22964
rect 4344 22918 4396 22924
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 4356 22506 4384 22918
rect 4724 22778 4752 23122
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3344 20420 3464 20448
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3056 19440 3108 19446
rect 2884 19366 3004 19394
rect 3056 19382 3108 19388
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2884 18834 2912 19246
rect 2976 18834 3004 19366
rect 3068 18970 3096 19382
rect 3160 19378 3188 20198
rect 3344 19990 3372 20420
rect 3424 20324 3476 20330
rect 3424 20266 3476 20272
rect 3436 20058 3464 20266
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3146 19136 3202 19145
rect 3146 19071 3202 19080
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2884 18358 2912 18770
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 3068 18222 3096 18906
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 3056 18216 3108 18222
rect 3160 18204 3188 19071
rect 3252 18358 3280 19654
rect 3436 19310 3464 19994
rect 3516 19984 3568 19990
rect 3988 19961 4016 22374
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4080 21418 4108 22034
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 4172 21690 4200 21898
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 4250 20632 4306 20641
rect 4068 20596 4120 20602
rect 4250 20567 4306 20576
rect 4068 20538 4120 20544
rect 4080 20482 4108 20538
rect 4264 20534 4292 20567
rect 4252 20528 4304 20534
rect 4080 20454 4200 20482
rect 4252 20470 4304 20476
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3516 19926 3568 19932
rect 3974 19952 4030 19961
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3160 18176 3280 18204
rect 3056 18158 3108 18164
rect 3068 17882 3096 18158
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16522 2636 17138
rect 3160 16998 3188 17682
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3160 16726 3188 16934
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2792 14958 2820 15438
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2136 13864 2188 13870
rect 1688 13530 1716 13806
rect 1780 13786 1900 13814
rect 1964 13786 2084 13814
rect 2136 13806 2188 13812
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1596 11898 1624 12271
rect 1688 12170 1716 12718
rect 1872 12646 1900 13786
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10198 1440 11154
rect 1400 10192 1452 10198
rect 1400 10134 1452 10140
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1596 8634 1624 9415
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1872 6458 1900 12582
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 2056 6186 2084 13786
rect 2148 7954 2176 13806
rect 2424 13530 2452 14418
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2240 12986 2268 13398
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2424 12306 2452 12854
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11898 2452 12242
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2412 11212 2464 11218
rect 2516 11200 2544 14826
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 14074 2728 14350
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2792 13802 2820 14894
rect 2884 14822 2912 15982
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2884 13734 2912 14214
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 12986 2636 13330
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2780 11212 2832 11218
rect 2516 11172 2636 11200
rect 2412 11154 2464 11160
rect 2424 10266 2452 11154
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2516 10674 2544 11018
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2424 10130 2452 10202
rect 2516 10130 2544 10610
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2424 9722 2452 10066
rect 2516 9722 2544 10066
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2608 7478 2636 11172
rect 2780 11154 2832 11160
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 10130 2728 10542
rect 2792 10538 2820 11154
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 9586 2728 10066
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2792 9110 2820 10474
rect 2884 10266 2912 12242
rect 2976 11558 3004 14826
rect 3068 14482 3096 15846
rect 3160 15706 3188 16662
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 3054 14376 3110 14385
rect 3054 14311 3110 14320
rect 3068 13530 3096 14311
rect 3160 14006 3188 14758
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 3252 13814 3280 18176
rect 3160 13786 3280 13814
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3160 12730 3188 13786
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3252 12832 3280 13466
rect 3344 13462 3372 19110
rect 3528 18766 3556 19926
rect 4080 19938 4108 20334
rect 4172 20262 4200 20454
rect 4252 20392 4304 20398
rect 4356 20380 4384 22442
rect 4724 22438 4752 22714
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4448 21010 4476 21354
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4448 20806 4476 20946
rect 4632 20942 4660 22034
rect 4816 21690 4844 23666
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4712 21616 4764 21622
rect 4712 21558 4764 21564
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4528 20868 4580 20874
rect 4528 20810 4580 20816
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 4304 20352 4384 20380
rect 4252 20334 4304 20340
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4080 19910 4200 19938
rect 3974 19887 4030 19896
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3790 19408 3846 19417
rect 3700 19372 3752 19378
rect 3790 19343 3846 19352
rect 3700 19314 3752 19320
rect 3712 18873 3740 19314
rect 3804 19292 3832 19343
rect 3884 19304 3936 19310
rect 3804 19264 3884 19292
rect 3884 19246 3936 19252
rect 3988 19174 4016 19790
rect 4172 19334 4200 19910
rect 4264 19718 4292 20334
rect 4448 19718 4476 20742
rect 4540 20602 4568 20810
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4540 19922 4568 20538
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4632 19990 4660 20470
rect 4724 20330 4752 21558
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4436 19712 4488 19718
rect 4436 19654 4488 19660
rect 4448 19378 4476 19654
rect 4540 19514 4568 19858
rect 4724 19786 4752 20266
rect 4816 20058 4844 21422
rect 4908 21146 4936 25162
rect 5000 24614 5028 27542
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 5276 27130 5304 27474
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5368 26858 5396 28494
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 5356 26852 5408 26858
rect 5356 26794 5408 26800
rect 5184 26246 5212 26794
rect 5264 26784 5316 26790
rect 5264 26726 5316 26732
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 5184 25770 5212 26182
rect 5276 25974 5304 26726
rect 5460 26518 5488 27066
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5264 25968 5316 25974
rect 5264 25910 5316 25916
rect 5080 25764 5132 25770
rect 5080 25706 5132 25712
rect 5172 25764 5224 25770
rect 5172 25706 5224 25712
rect 5092 25498 5120 25706
rect 5080 25492 5132 25498
rect 5080 25434 5132 25440
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5276 24682 5304 25298
rect 5552 24682 5580 31078
rect 5644 28082 5672 31418
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5644 25974 5672 28018
rect 5736 26194 5764 34682
rect 6000 34536 6052 34542
rect 6000 34478 6052 34484
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 5920 30870 5948 31622
rect 5908 30864 5960 30870
rect 5908 30806 5960 30812
rect 5920 30394 5948 30806
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 5920 29306 5948 29650
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 5828 26994 5856 27270
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5736 26166 5856 26194
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 5632 25968 5684 25974
rect 5632 25910 5684 25916
rect 5644 24818 5672 25910
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5172 24676 5224 24682
rect 5172 24618 5224 24624
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 5184 24342 5212 24618
rect 5276 24410 5304 24618
rect 5356 24608 5408 24614
rect 5356 24550 5408 24556
rect 5264 24404 5316 24410
rect 5264 24346 5316 24352
rect 5172 24336 5224 24342
rect 5172 24278 5224 24284
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4080 19306 4200 19334
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4816 19310 4844 19722
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3698 18864 3754 18873
rect 3698 18799 3754 18808
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3436 16538 3464 18702
rect 4080 18698 4108 19306
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4172 19145 4200 19178
rect 4252 19168 4304 19174
rect 4158 19136 4214 19145
rect 4712 19168 4764 19174
rect 4252 19110 4304 19116
rect 4632 19128 4712 19156
rect 4158 19071 4214 19080
rect 4068 18692 4120 18698
rect 4068 18634 4120 18640
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 4080 18426 4108 18634
rect 4264 18630 4292 19110
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18426 4292 18566
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3436 16510 3556 16538
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16114 3464 16390
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15706 3464 16050
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3528 15586 3556 16510
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3436 15558 3556 15586
rect 3436 14958 3464 15558
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 14482 3464 14894
rect 3528 14618 3556 15302
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3988 14822 4016 18158
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 17338 4108 17614
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3436 13938 3464 14418
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 13530 3464 13738
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3252 12804 3372 12832
rect 3160 12702 3280 12730
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2976 9518 3004 11086
rect 3068 11082 3096 12038
rect 3160 11286 3188 12582
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 9178 3004 9454
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 478 54 704 82
rect 1490 82 1546 480
rect 1780 82 1808 2790
rect 1490 54 1808 82
rect 2594 82 2650 480
rect 2884 82 2912 8570
rect 3068 8566 3096 10678
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3160 9722 3188 9930
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3252 9586 3280 12702
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3344 8838 3372 12804
rect 3436 11898 3464 13262
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 10452 3464 11494
rect 3528 11354 3556 13670
rect 3620 13326 3648 13806
rect 3988 13734 4016 14418
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 4080 12050 4108 17070
rect 4264 16998 4292 18362
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 15366 4200 16526
rect 4264 16250 4292 16662
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4264 15910 4292 16186
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4264 15094 4292 15574
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4172 12918 4200 14894
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 13530 4292 14758
rect 4356 14618 4384 18702
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4448 14550 4476 15846
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4448 12986 4476 14010
rect 4540 13841 4568 15302
rect 4526 13832 4582 13841
rect 4526 13767 4582 13776
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 3988 12022 4108 12050
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3988 10742 4016 12022
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4080 11218 4108 11834
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 11218 4200 11494
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3516 10464 3568 10470
rect 3436 10424 3516 10452
rect 3516 10406 3568 10412
rect 3528 9382 3556 10406
rect 3988 10062 4016 10542
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10198 4108 10406
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4172 10062 4200 11154
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10674 4292 10950
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4264 10130 4292 10610
rect 4356 10606 4384 11154
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4448 10130 4476 12786
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12442 4568 12650
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 3976 10056 4028 10062
rect 3974 10024 3976 10033
rect 4160 10056 4212 10062
rect 4028 10024 4030 10033
rect 3974 9959 4030 9968
rect 4080 10004 4160 10010
rect 4080 9998 4212 10004
rect 4080 9982 4200 9998
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3988 9722 4016 9959
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4080 9654 4108 9982
rect 4264 9722 4292 10066
rect 4342 10024 4398 10033
rect 4342 9959 4398 9968
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3528 9042 3556 9318
rect 4264 9042 4292 9658
rect 4356 9518 4384 9959
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 3332 8832 3384 8838
rect 3384 8780 3464 8786
rect 3332 8774 3464 8780
rect 3344 8758 3464 8774
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7546 3004 7890
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2976 7274 3004 7482
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 3068 6730 3096 8502
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 8090 3372 8434
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3436 7342 3464 8758
rect 3528 8634 3556 8978
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 8090 3832 8298
rect 3988 8294 4016 8842
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 7002 3464 7278
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 2594 54 2912 82
rect 3436 82 3464 4218
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3988 3194 4016 8230
rect 4080 7750 4108 8502
rect 4448 7954 4476 9522
rect 4632 8430 4660 19128
rect 4712 19110 4764 19116
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4724 18222 4752 18634
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4816 18068 4844 18294
rect 4724 18040 4844 18068
rect 4724 13326 4752 18040
rect 4908 17678 4936 19926
rect 5000 19242 5028 23190
rect 5092 20534 5120 23598
rect 5172 22568 5224 22574
rect 5368 22556 5396 24550
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5552 23254 5580 23802
rect 5644 23662 5672 24006
rect 5632 23656 5684 23662
rect 5632 23598 5684 23604
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5644 23186 5672 23598
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22642 5488 23054
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5644 22574 5672 23122
rect 5224 22528 5396 22556
rect 5632 22568 5684 22574
rect 5172 22510 5224 22516
rect 5632 22510 5684 22516
rect 5184 21894 5212 22510
rect 5644 22098 5672 22510
rect 5632 22092 5684 22098
rect 5632 22034 5684 22040
rect 5644 21894 5672 22034
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 20602 5672 21830
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5080 20528 5132 20534
rect 5080 20470 5132 20476
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 5000 17814 5028 18566
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5092 17814 5120 18090
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 5000 17678 5028 17750
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4988 17672 5040 17678
rect 5184 17660 5212 20334
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5276 18902 5304 19382
rect 5552 19174 5580 19654
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18902 5580 19110
rect 5264 18896 5316 18902
rect 5540 18896 5592 18902
rect 5316 18856 5488 18884
rect 5264 18838 5316 18844
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5276 18154 5304 18702
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5276 17882 5304 18090
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 4988 17614 5040 17620
rect 5092 17632 5212 17660
rect 5000 17338 5028 17614
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 16114 4844 16526
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4804 15972 4856 15978
rect 4908 15960 4936 16458
rect 4856 15932 4936 15960
rect 4804 15914 4856 15920
rect 5000 15638 5028 16934
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4908 15026 4936 15370
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14006 4844 14214
rect 5000 14074 5028 15574
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4802 13832 4858 13841
rect 5092 13814 5120 17632
rect 5368 17610 5396 18362
rect 5460 18358 5488 18856
rect 5540 18838 5592 18844
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5552 18222 5580 18838
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5356 17604 5408 17610
rect 5408 17564 5488 17592
rect 5356 17546 5408 17552
rect 5356 17060 5408 17066
rect 5276 17020 5356 17048
rect 5276 16454 5304 17020
rect 5356 17002 5408 17008
rect 5460 16726 5488 17564
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5276 15162 5304 16390
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5184 14822 5212 15030
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14550 5212 14758
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 4802 13767 4858 13776
rect 4908 13786 5120 13814
rect 4816 13734 4844 13767
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4816 13190 4844 13330
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4724 12102 4752 12242
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 9586 4752 12038
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4816 9110 4844 13126
rect 4908 12782 4936 13786
rect 5184 13530 5212 14350
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4632 8022 4660 8366
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7342 4108 7686
rect 4448 7546 4476 7890
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4908 7426 4936 12718
rect 5000 11898 5028 13194
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5000 10810 5028 11834
rect 5092 11762 5120 13398
rect 5184 12918 5212 13466
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 11354 5120 11698
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9178 5212 10066
rect 5276 9586 5304 14554
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5368 13870 5396 14010
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 13734 5396 13806
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5460 13462 5488 14010
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5368 12986 5396 13262
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5552 10606 5580 18158
rect 5736 15570 5764 25978
rect 5828 25838 5856 26166
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 5828 24886 5856 25774
rect 5816 24880 5868 24886
rect 5816 24822 5868 24828
rect 5920 24274 5948 29242
rect 6012 27402 6040 34478
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6276 34060 6328 34066
rect 6276 34002 6328 34008
rect 6104 33318 6132 34002
rect 6288 33658 6316 34002
rect 6276 33652 6328 33658
rect 6276 33594 6328 33600
rect 6288 33386 6316 33594
rect 6644 33448 6696 33454
rect 6644 33390 6696 33396
rect 6276 33380 6328 33386
rect 6276 33322 6328 33328
rect 6092 33312 6144 33318
rect 6092 33254 6144 33260
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6656 32774 6684 33390
rect 6644 32768 6696 32774
rect 6644 32710 6696 32716
rect 6656 32230 6684 32710
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6748 30274 6776 34682
rect 6840 34610 6868 35226
rect 7012 35216 7064 35222
rect 7012 35158 7064 35164
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 7024 34474 7052 35158
rect 7116 34678 7144 39630
rect 7378 39520 7434 39630
rect 8574 39658 8630 40000
rect 9678 39658 9734 40000
rect 10782 39658 10838 40000
rect 11978 39658 12034 40000
rect 13082 39658 13138 40000
rect 14278 39658 14334 40000
rect 8574 39630 8800 39658
rect 8574 39520 8630 39630
rect 8300 35556 8352 35562
rect 8300 35498 8352 35504
rect 8392 35556 8444 35562
rect 8392 35498 8444 35504
rect 8312 35290 8340 35498
rect 8300 35284 8352 35290
rect 8300 35226 8352 35232
rect 8300 34944 8352 34950
rect 8404 34932 8432 35498
rect 8352 34904 8432 34932
rect 8300 34886 8352 34892
rect 7104 34672 7156 34678
rect 7104 34614 7156 34620
rect 7564 34672 7616 34678
rect 7564 34614 7616 34620
rect 7012 34468 7064 34474
rect 7012 34410 7064 34416
rect 7024 33862 7052 34410
rect 7472 34128 7524 34134
rect 7472 34070 7524 34076
rect 7012 33856 7064 33862
rect 7012 33798 7064 33804
rect 7024 33658 7052 33798
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 7484 33386 7512 34070
rect 6920 33380 6972 33386
rect 6920 33322 6972 33328
rect 7472 33380 7524 33386
rect 7472 33322 7524 33328
rect 6932 32774 6960 33322
rect 7484 33114 7512 33322
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6932 32434 6960 32710
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 7012 32292 7064 32298
rect 7012 32234 7064 32240
rect 6920 31952 6972 31958
rect 6920 31894 6972 31900
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6840 31482 6868 31758
rect 6828 31476 6880 31482
rect 6828 31418 6880 31424
rect 6932 31414 6960 31894
rect 7024 31822 7052 32234
rect 7116 31958 7144 32846
rect 7484 32570 7512 33050
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7104 31952 7156 31958
rect 7104 31894 7156 31900
rect 7012 31816 7064 31822
rect 7012 31758 7064 31764
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 7024 30870 7052 31758
rect 7012 30864 7064 30870
rect 7012 30806 7064 30812
rect 6656 30246 6776 30274
rect 7012 30252 7064 30258
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6092 28552 6144 28558
rect 6092 28494 6144 28500
rect 6104 27946 6132 28494
rect 6196 28218 6224 28698
rect 6656 28370 6684 30246
rect 7012 30194 7064 30200
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6748 28490 6776 30126
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6840 29782 6868 29990
rect 6828 29776 6880 29782
rect 6828 29718 6880 29724
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6932 29170 6960 29446
rect 7024 29238 7052 30194
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 7012 29232 7064 29238
rect 7012 29174 7064 29180
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 6932 28762 6960 29106
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6736 28484 6788 28490
rect 6736 28426 6788 28432
rect 6656 28342 6776 28370
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6092 27940 6144 27946
rect 6092 27882 6144 27888
rect 6104 27606 6132 27882
rect 6196 27606 6224 28154
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6092 27600 6144 27606
rect 6092 27542 6144 27548
rect 6184 27600 6236 27606
rect 6184 27542 6236 27548
rect 6000 27396 6052 27402
rect 6000 27338 6052 27344
rect 6196 27130 6224 27542
rect 6184 27124 6236 27130
rect 6184 27066 6236 27072
rect 6644 26852 6696 26858
rect 6644 26794 6696 26800
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 6012 25294 6040 26726
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6276 26512 6328 26518
rect 6276 26454 6328 26460
rect 6288 26042 6316 26454
rect 6656 26382 6684 26794
rect 6644 26376 6696 26382
rect 6644 26318 6696 26324
rect 6460 26308 6512 26314
rect 6460 26250 6512 26256
rect 6472 26042 6500 26250
rect 6276 26036 6328 26042
rect 6196 25996 6276 26024
rect 6196 25362 6224 25996
rect 6276 25978 6328 25984
rect 6460 26036 6512 26042
rect 6460 25978 6512 25984
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 6012 24886 6040 25230
rect 6748 25226 6776 28342
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6736 25220 6788 25226
rect 6736 25162 6788 25168
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 6840 24818 6868 25094
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5920 22574 5948 22918
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 5906 21584 5962 21593
rect 5906 21519 5962 21528
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 19922 5856 21286
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5828 17542 5856 19450
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5920 17134 5948 21519
rect 6012 20992 6040 24618
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6840 24410 6868 24754
rect 6932 24614 6960 25298
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 6288 23866 6316 24210
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6184 23588 6236 23594
rect 6184 23530 6236 23536
rect 6196 23118 6224 23530
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6196 22234 6224 23054
rect 6656 22778 6684 23190
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6552 22160 6604 22166
rect 6656 22148 6684 22374
rect 6604 22120 6684 22148
rect 6552 22102 6604 22108
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6380 21554 6408 21966
rect 6564 21690 6592 22102
rect 6748 22030 6776 22986
rect 6840 22982 6868 23598
rect 6828 22976 6880 22982
rect 6828 22918 6880 22924
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6368 21548 6420 21554
rect 6368 21490 6420 21496
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6748 21146 6776 21966
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6932 21078 6960 21422
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6184 21004 6236 21010
rect 6012 20964 6184 20992
rect 6184 20946 6236 20952
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 6012 19718 6040 20742
rect 6090 20632 6146 20641
rect 6090 20567 6146 20576
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6012 19310 6040 19654
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 18970 6040 19246
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 6104 17814 6132 20567
rect 6196 20398 6224 20946
rect 7024 20584 7052 29174
rect 7116 28966 7144 29718
rect 7576 29170 7604 34614
rect 7932 34400 7984 34406
rect 7932 34342 7984 34348
rect 7944 34066 7972 34342
rect 8312 34202 8340 34886
rect 8576 34604 8628 34610
rect 8576 34546 8628 34552
rect 8588 34202 8616 34546
rect 8668 34468 8720 34474
rect 8668 34410 8720 34416
rect 8300 34196 8352 34202
rect 8300 34138 8352 34144
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 7932 34060 7984 34066
rect 7932 34002 7984 34008
rect 8392 33856 8444 33862
rect 8392 33798 8444 33804
rect 8116 31136 8168 31142
rect 8116 31078 8168 31084
rect 8128 30938 8156 31078
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 7840 30728 7892 30734
rect 7840 30670 7892 30676
rect 7852 29782 7880 30670
rect 8128 30326 8156 30874
rect 8116 30320 8168 30326
rect 8116 30262 8168 30268
rect 8128 30122 8156 30262
rect 8116 30116 8168 30122
rect 8116 30058 8168 30064
rect 7840 29776 7892 29782
rect 7840 29718 7892 29724
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8116 29028 8168 29034
rect 8116 28970 8168 28976
rect 7104 28960 7156 28966
rect 7104 28902 7156 28908
rect 7116 28626 7144 28902
rect 8128 28694 8156 28970
rect 8116 28688 8168 28694
rect 8116 28630 8168 28636
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7748 28416 7800 28422
rect 7748 28358 7800 28364
rect 7760 28218 7788 28358
rect 7748 28212 7800 28218
rect 7748 28154 7800 28160
rect 8128 27674 8156 28630
rect 8312 28558 8340 29106
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 8404 27606 8432 33798
rect 8680 33658 8708 34410
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8576 33448 8628 33454
rect 8576 33390 8628 33396
rect 8588 32842 8616 33390
rect 8668 33312 8720 33318
rect 8668 33254 8720 33260
rect 8576 32836 8628 32842
rect 8576 32778 8628 32784
rect 8680 32366 8708 33254
rect 8668 32360 8720 32366
rect 8668 32302 8720 32308
rect 8484 32224 8536 32230
rect 8484 32166 8536 32172
rect 8496 30258 8524 32166
rect 8680 31686 8708 32302
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8496 29850 8524 30194
rect 8484 29844 8536 29850
rect 8484 29786 8536 29792
rect 8668 29708 8720 29714
rect 8772 29696 8800 39630
rect 9678 39630 9996 39658
rect 9678 39520 9734 39630
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9324 34610 9352 35566
rect 9680 35148 9732 35154
rect 9680 35090 9732 35096
rect 9692 34746 9720 35090
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9312 34604 9364 34610
rect 9312 34546 9364 34552
rect 9324 33930 9352 34546
rect 9588 34128 9640 34134
rect 9588 34070 9640 34076
rect 9312 33924 9364 33930
rect 9312 33866 9364 33872
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9312 33584 9364 33590
rect 9312 33526 9364 33532
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8720 29668 8800 29696
rect 8668 29650 8720 29656
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29170 8524 29446
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8680 28966 8708 29650
rect 9324 29646 9352 33526
rect 9600 33318 9628 34070
rect 9784 33998 9812 35022
rect 9968 34746 9996 39630
rect 10520 39630 10838 39658
rect 10046 38312 10102 38321
rect 10046 38247 10102 38256
rect 10060 35834 10088 38247
rect 10048 35828 10100 35834
rect 10048 35770 10100 35776
rect 10520 35290 10548 39630
rect 10782 39520 10838 39630
rect 11532 39630 12034 39658
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 11058 35048 11114 35057
rect 11058 34983 11114 34992
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9784 33658 9812 33934
rect 10060 33862 10088 34478
rect 10048 33856 10100 33862
rect 10048 33798 10100 33804
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 9588 33312 9640 33318
rect 9588 33254 9640 33260
rect 9600 33114 9628 33254
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32366 10088 32710
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 10048 32360 10100 32366
rect 10048 32302 10100 32308
rect 9692 32230 9720 32302
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 10048 32224 10100 32230
rect 10048 32166 10100 32172
rect 9692 31890 9720 32166
rect 9772 32020 9824 32026
rect 9772 31962 9824 31968
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9496 31680 9548 31686
rect 9496 31622 9548 31628
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9324 29170 9352 29582
rect 9312 29164 9364 29170
rect 9312 29106 9364 29112
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8760 28008 8812 28014
rect 8760 27950 8812 27956
rect 8392 27600 8444 27606
rect 8392 27542 8444 27548
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7944 27130 7972 27406
rect 8404 27130 8432 27542
rect 8772 27402 8800 27950
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 8760 27396 8812 27402
rect 8760 27338 8812 27344
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 7932 27124 7984 27130
rect 7932 27066 7984 27072
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 7656 26852 7708 26858
rect 7656 26794 7708 26800
rect 7668 25906 7696 26794
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7760 25786 7788 26998
rect 8864 26994 8892 27270
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8668 26852 8720 26858
rect 8668 26794 8720 26800
rect 8680 26586 8708 26794
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 7932 26512 7984 26518
rect 7932 26454 7984 26460
rect 7840 26376 7892 26382
rect 7840 26318 7892 26324
rect 7668 25758 7788 25786
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 24138 7144 25094
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 7116 23526 7144 24074
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7116 23254 7144 23462
rect 7104 23248 7156 23254
rect 7104 23190 7156 23196
rect 7116 22506 7144 23190
rect 7208 23186 7236 25638
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7116 21418 7144 22442
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7208 20602 7236 20946
rect 7196 20596 7248 20602
rect 7024 20556 7144 20584
rect 7010 20496 7066 20505
rect 7010 20431 7066 20440
rect 7024 20398 7052 20431
rect 6184 20392 6236 20398
rect 7012 20392 7064 20398
rect 6184 20334 6236 20340
rect 6642 20360 6698 20369
rect 7012 20334 7064 20340
rect 6642 20295 6698 20304
rect 6656 20262 6684 20295
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6748 19174 6776 19858
rect 7116 19718 7144 20556
rect 7196 20538 7248 20544
rect 7208 20058 7236 20538
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6472 18290 6500 18770
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6092 17808 6144 17814
rect 6092 17750 6144 17756
rect 6012 17542 6040 17750
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 6012 16998 6040 17478
rect 6104 17066 6132 17750
rect 6656 17610 6684 18294
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6656 17202 6684 17546
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5920 16250 5948 16662
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5736 14074 5764 14486
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5644 12306 5672 13942
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5644 12170 5672 12242
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11354 5672 12106
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5736 11218 5764 12786
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10266 5580 10542
rect 5736 10266 5764 11154
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9722 5396 9998
rect 5448 9988 5500 9994
rect 5552 9976 5580 10202
rect 5500 9948 5580 9976
rect 5448 9930 5500 9936
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4724 7398 4936 7426
rect 5000 7410 5028 7686
rect 4988 7404 5040 7410
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 6390 4108 6802
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5370 4660 6054
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5166 4752 7398
rect 4988 7346 5040 7352
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4908 6866 4936 7278
rect 5184 6934 5212 7822
rect 5276 7002 5304 9522
rect 5552 9518 5580 9948
rect 5828 9674 5856 14826
rect 6012 13530 6040 16934
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6104 15910 6132 16662
rect 6196 16590 6224 17070
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6656 16658 6684 17138
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 14618 6132 15846
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15162 6316 15506
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5920 12646 5948 13398
rect 6196 12782 6224 13738
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6748 12918 6776 19110
rect 6932 17202 6960 19382
rect 7116 19310 7144 19654
rect 7208 19310 7236 19994
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7024 17678 7052 18090
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6840 14482 6868 17002
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 14822 6960 15370
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7024 13938 7052 14418
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6840 12782 6868 13194
rect 6932 12986 6960 13670
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5920 12374 5948 12582
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 6012 12306 6040 12582
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6840 12442 6868 12718
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11898 6040 12242
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6012 11218 6040 11834
rect 6196 11694 6224 12174
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11762 6500 12038
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6012 10810 6040 11154
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 10606 6040 10746
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5644 9646 5856 9674
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5552 9178 5580 9454
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5460 7206 5488 7958
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6254 4936 6802
rect 5460 6662 5488 7142
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4690 4752 5102
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4282 4200 4422
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 3194 4568 3470
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 2650 4016 2926
rect 4816 2854 4844 4966
rect 4908 4690 4936 5850
rect 5460 5098 5488 6598
rect 5644 5778 5672 9646
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5644 5370 5672 5714
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4214 4936 4626
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5000 4214 5028 4490
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4908 3602 4936 4150
rect 5092 3738 5120 4558
rect 5264 4004 5316 4010
rect 5368 3992 5396 4762
rect 5644 4729 5672 5306
rect 5828 4826 5856 8502
rect 5920 7410 5948 10474
rect 6012 10130 6040 10542
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9722 6040 10066
rect 6932 10062 6960 11562
rect 7024 11558 7052 12310
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11286 7052 11494
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 7024 11014 7052 11222
rect 7116 11082 7144 19246
rect 7208 18834 7236 19246
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7208 18086 7236 18770
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7300 16946 7328 23122
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7484 22234 7512 22578
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7484 18902 7512 19790
rect 7576 19378 7604 20742
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17202 7420 17818
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7300 16918 7420 16946
rect 7392 15745 7420 16918
rect 7484 16794 7512 17002
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7484 16250 7512 16730
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7484 15978 7512 16186
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7378 15736 7434 15745
rect 7378 15671 7434 15680
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 14958 7236 15302
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7208 14414 7236 14894
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 13530 7236 14214
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7300 13530 7328 13942
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 11150 7328 12582
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10538 7052 10950
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7116 10198 7144 10542
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7208 10130 7236 11086
rect 7300 10810 7328 11086
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 7208 9722 7236 10066
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 8090 6040 8910
rect 6656 8294 6684 9046
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6196 7750 6224 8230
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6552 7744 6604 7750
rect 6656 7732 6684 8230
rect 6604 7704 6684 7732
rect 6552 7686 6604 7692
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6196 6934 6224 7686
rect 6288 7546 6316 7686
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6748 6934 6776 8910
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8294 7144 8774
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7478 6868 7890
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 7002 7052 7346
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6458 6132 6734
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6104 5914 6132 6394
rect 6196 6390 6224 6870
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5630 4720 5686 4729
rect 5630 4655 5686 4664
rect 5828 4554 5856 4762
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5920 4010 5948 5238
rect 6748 5234 6776 6870
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4758 6132 4966
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6748 4826 6776 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4282 6040 4558
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4214 6132 4694
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 5316 3964 5396 3992
rect 5448 4004 5500 4010
rect 5264 3946 5316 3952
rect 5448 3946 5500 3952
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4908 3058 4936 3538
rect 5092 3058 5120 3674
rect 5460 3398 5488 3946
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5460 3194 5488 3334
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4908 2650 4936 2994
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5552 2378 5580 3334
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3606 82 3662 480
rect 3436 54 3662 82
rect 4540 82 4568 2246
rect 4710 82 4766 480
rect 4540 54 4766 82
rect 5736 82 5764 3062
rect 5920 2378 5948 3946
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6196 2922 6224 3674
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 3194 6592 3470
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 6196 2310 6224 2858
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 2582 6684 3878
rect 6840 3738 6868 4966
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 6748 2514 6776 2926
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 5814 82 5870 480
rect 5736 54 5870 82
rect 478 0 534 54
rect 1490 0 1546 54
rect 2594 0 2650 54
rect 3606 0 3662 54
rect 4710 0 4766 54
rect 5814 0 5870 54
rect 6826 82 6882 480
rect 6932 82 6960 2926
rect 7024 2446 7052 6122
rect 7208 5778 7236 9522
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 8090 7328 8434
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 4826 7236 5714
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7208 3058 7236 4762
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4146 7328 4558
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3738 7328 4082
rect 7392 4010 7420 15671
rect 7484 15638 7512 15914
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7484 15094 7512 15574
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14074 7512 14894
rect 7668 14890 7696 25758
rect 7852 25430 7880 26318
rect 7944 25702 7972 26454
rect 8680 26042 8708 26522
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 7944 25158 7972 25638
rect 8864 25498 8892 26930
rect 9416 26586 9444 27406
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8944 25900 8996 25906
rect 8944 25842 8996 25848
rect 8956 25498 8984 25842
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9416 25430 9444 25638
rect 9404 25424 9456 25430
rect 9404 25366 9456 25372
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 8404 24682 8432 25298
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 7748 24676 7800 24682
rect 7748 24618 7800 24624
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 7760 22488 7788 24618
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23798 7880 24142
rect 7840 23792 7892 23798
rect 7840 23734 7892 23740
rect 7852 23322 7880 23734
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7944 23186 7972 24618
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 8036 24342 8064 24550
rect 8024 24336 8076 24342
rect 8024 24278 8076 24284
rect 8036 23526 8064 24278
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 8036 23050 8064 23462
rect 8220 23254 8248 23598
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8024 23044 8076 23050
rect 8024 22986 8076 22992
rect 7932 22500 7984 22506
rect 7760 22460 7932 22488
rect 7932 22442 7984 22448
rect 7944 22166 7972 22442
rect 8128 22234 8156 23054
rect 8220 22438 8248 23190
rect 8404 22778 8432 23530
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21486 7880 21830
rect 8220 21690 8248 22102
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 7840 21480 7892 21486
rect 7840 21422 7892 21428
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8128 21146 8156 21354
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8128 20602 8156 21082
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20596 8168 20602
rect 8036 20556 8116 20584
rect 8036 20330 8064 20556
rect 8116 20538 8168 20544
rect 8220 20466 8248 20742
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 8036 19990 8064 20266
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 8036 19446 8064 19926
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 8128 18834 8156 20334
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19242 8432 19654
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 8128 18426 8156 18770
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7852 17066 7880 17682
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7656 14884 7708 14890
rect 7656 14826 7708 14832
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7852 12850 7880 17002
rect 8036 16114 8064 17614
rect 8220 16572 8248 19110
rect 8404 18970 8432 19178
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8496 18612 8524 24686
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8680 23730 8708 24006
rect 8864 23730 8892 24142
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8588 22506 8616 22918
rect 8680 22710 8708 23666
rect 8864 23254 8892 23666
rect 9324 23254 9352 24618
rect 9508 23474 9536 31622
rect 9692 31278 9720 31826
rect 9784 31346 9812 31962
rect 10060 31958 10088 32166
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 10244 31890 10272 32234
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10968 31884 11020 31890
rect 10968 31826 11020 31832
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 10152 31346 10180 31622
rect 10416 31408 10468 31414
rect 10416 31350 10468 31356
rect 9772 31340 9824 31346
rect 9772 31282 9824 31288
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 9680 31272 9732 31278
rect 9680 31214 9732 31220
rect 9954 31240 10010 31249
rect 9954 31175 10010 31184
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9600 30054 9628 31078
rect 9864 30864 9916 30870
rect 9864 30806 9916 30812
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9784 30394 9812 30670
rect 9876 30394 9904 30806
rect 9772 30388 9824 30394
rect 9772 30330 9824 30336
rect 9864 30388 9916 30394
rect 9864 30330 9916 30336
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9968 29832 9996 31175
rect 10152 30240 10180 31282
rect 10232 31204 10284 31210
rect 10232 31146 10284 31152
rect 10244 30938 10272 31146
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 10428 30870 10456 31350
rect 10980 31142 11008 31826
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10416 30864 10468 30870
rect 10416 30806 10468 30812
rect 10428 30258 10456 30806
rect 10416 30252 10468 30258
rect 10152 30212 10272 30240
rect 10140 30116 10192 30122
rect 10140 30058 10192 30064
rect 10152 29850 10180 30058
rect 9784 29804 9996 29832
rect 10140 29844 10192 29850
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9692 29238 9720 29650
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9416 23446 9536 23474
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8680 21146 8708 22374
rect 8864 22030 8892 23190
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8760 21956 8812 21962
rect 8760 21898 8812 21904
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8772 19446 8800 21898
rect 8864 21690 8892 21966
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9416 19922 9444 23446
rect 9600 22574 9628 28902
rect 9784 28744 9812 29804
rect 10140 29786 10192 29792
rect 9864 29708 9916 29714
rect 9864 29650 9916 29656
rect 9876 28966 9904 29650
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9692 28716 9812 28744
rect 9692 24177 9720 28716
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9784 28218 9812 28562
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9876 26858 9904 28902
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9968 28082 9996 28358
rect 10152 28082 10180 29786
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10060 27606 10088 27882
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 9956 27396 10008 27402
rect 9956 27338 10008 27344
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9968 26790 9996 27338
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26512 9916 26518
rect 9864 26454 9916 26460
rect 9876 25430 9904 26454
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 10060 25770 10088 25978
rect 10152 25906 10180 28018
rect 10244 27470 10272 30212
rect 10416 30194 10468 30200
rect 10980 29714 11008 31078
rect 10968 29708 11020 29714
rect 10968 29650 11020 29656
rect 11072 28626 11100 34983
rect 11244 34536 11296 34542
rect 11244 34478 11296 34484
rect 11060 28620 11112 28626
rect 10980 28580 11060 28608
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 26994 10272 27406
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10244 26518 10272 26930
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10888 26042 10916 26318
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10140 25900 10192 25906
rect 10140 25842 10192 25848
rect 9956 25764 10008 25770
rect 9956 25706 10008 25712
rect 10048 25764 10100 25770
rect 10048 25706 10100 25712
rect 9968 25498 9996 25706
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9864 25424 9916 25430
rect 9864 25366 9916 25372
rect 10152 25294 10180 25842
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 9784 24954 9812 25230
rect 10428 24954 10456 25366
rect 10508 25220 10560 25226
rect 10508 25162 10560 25168
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 9678 24168 9734 24177
rect 9678 24103 9734 24112
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9496 22500 9548 22506
rect 9496 22442 9548 22448
rect 9508 21962 9536 22442
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9508 21078 9536 21286
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9508 20602 9536 21014
rect 9600 21010 9628 21286
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9692 20040 9720 24103
rect 10060 23662 10088 24686
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9784 22778 9812 23190
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9876 22642 9904 23190
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9876 21622 9904 22102
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21690 9996 21830
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9864 21616 9916 21622
rect 10060 21593 10088 21966
rect 9864 21558 9916 21564
rect 10046 21584 10102 21593
rect 10046 21519 10102 21528
rect 10324 21412 10376 21418
rect 10324 21354 10376 21360
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 20058 9812 20742
rect 9876 20534 9904 21014
rect 10336 20874 10364 21354
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 9864 20528 9916 20534
rect 9864 20470 9916 20476
rect 9600 20012 9720 20040
rect 9772 20052 9824 20058
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8404 18584 8524 18612
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8312 16998 8340 18022
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16726 8340 16934
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8220 16544 8340 16572
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8128 15162 8156 15914
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8128 14482 8156 15098
rect 8220 14822 8248 15438
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14550 8248 14758
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7944 14074 7972 14282
rect 8128 14074 8156 14418
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7944 12646 7972 13398
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7944 12170 7972 12582
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7932 11552 7984 11558
rect 8036 11540 8064 12582
rect 7984 11512 8064 11540
rect 7932 11494 7984 11500
rect 7944 11286 7972 11494
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7484 8537 7512 9959
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 8838 7604 9454
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7470 8528 7526 8537
rect 7470 8463 7526 8472
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 7750 7512 8230
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6254 7512 7686
rect 7668 6458 7696 11018
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 10198 8156 10474
rect 8220 10266 8248 10610
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7760 7954 7788 9386
rect 8128 9382 8156 10134
rect 8312 9654 8340 16544
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7852 8634 7880 8842
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8128 8090 8156 9318
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7002 7788 7890
rect 8128 7206 8156 8026
rect 8220 7410 8248 8910
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7484 5778 7512 6190
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7668 4214 7696 4694
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7392 2990 7420 3946
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7208 2310 7236 2518
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6826 54 6960 82
rect 7760 82 7788 6666
rect 7852 6322 7880 6734
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7944 5846 7972 7142
rect 8128 7002 8156 7142
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8128 6118 8156 6938
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 3534 8064 5646
rect 8128 3942 8156 6054
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8220 4146 8248 4762
rect 8312 4282 8340 6394
rect 8404 4486 8432 18584
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16250 8524 16934
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8588 15910 8616 16526
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8588 14770 8616 15846
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8680 15162 8708 15302
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8680 14890 8708 15098
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8588 14742 8708 14770
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 12850 8524 14214
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8496 12442 8524 12786
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8588 8956 8616 14554
rect 8680 13734 8708 14742
rect 8772 14618 8800 19382
rect 9508 19242 9536 19790
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9508 18834 9536 19178
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9508 18290 9536 18770
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8864 17542 8892 18090
rect 9508 17814 9536 18226
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17338 8892 17478
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 16454 9352 17138
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9324 16182 9352 16390
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8864 15094 8892 15642
rect 9140 15638 9168 16050
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9416 15366 9444 16594
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 15978 9536 16050
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 15088 8904 15094
rect 9600 15076 9628 20012
rect 9772 19994 9824 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9692 19174 9720 19858
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9784 17882 9812 18906
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10152 18698 10180 18770
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10152 18426 10180 18634
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9876 17066 9904 17614
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 10152 16998 10180 17750
rect 10336 17660 10364 20810
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 18290 10456 18566
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10520 17746 10548 25162
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10612 19514 10640 23598
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10796 20398 10824 22510
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10416 17672 10468 17678
rect 10336 17632 10416 17660
rect 10416 17614 10468 17620
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9968 16726 9996 16934
rect 10152 16794 10180 16934
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9876 16114 9904 16662
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 15088 9732 15094
rect 9600 15048 9680 15076
rect 8852 15030 8904 15036
rect 9680 15030 9732 15036
rect 9784 14618 9812 15438
rect 9876 15162 9904 15574
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9968 14618 9996 15982
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10244 15162 10272 15370
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 14822 10272 15098
rect 10336 14890 10364 17206
rect 10428 17202 10456 17614
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10612 17066 10640 18022
rect 10704 17610 10732 18090
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10428 16590 10456 17002
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 15638 10456 16526
rect 10520 16250 10548 16934
rect 10612 16794 10640 17002
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10612 15026 10640 16730
rect 10796 16522 10824 17478
rect 10980 17066 11008 28580
rect 11060 28562 11112 28568
rect 11060 27600 11112 27606
rect 11060 27542 11112 27548
rect 11072 27130 11100 27542
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11256 25362 11284 34478
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 11440 31482 11468 31826
rect 11428 31476 11480 31482
rect 11428 31418 11480 31424
rect 11334 27976 11390 27985
rect 11334 27911 11390 27920
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 11256 24954 11284 25298
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11256 21418 11284 22034
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 16250 10824 16458
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 15026 10824 15302
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10336 14618 10364 14826
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8864 13870 8892 14350
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9692 14074 9720 14282
rect 9784 14074 9812 14554
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12850 8800 13194
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8864 12442 8892 13262
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 11626 8984 11698
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8772 11014 8800 11494
rect 8956 11354 8984 11562
rect 8944 11348 8996 11354
rect 8864 11308 8944 11336
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 9722 8800 10950
rect 8864 10810 8892 11308
rect 8944 11290 8996 11296
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8864 10470 8892 10746
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 9232 10266 9260 10474
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8588 8928 8892 8956
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8496 5574 8524 5714
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5166 8524 5510
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3670 8156 3878
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8036 3058 8064 3470
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8024 2848 8076 2854
rect 8128 2836 8156 3606
rect 8312 3466 8340 4218
rect 8496 3738 8524 4966
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8076 2808 8156 2836
rect 8024 2790 8076 2796
rect 8036 2310 8064 2790
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 7930 82 7986 480
rect 7760 54 7986 82
rect 8680 82 8708 7278
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6458 8800 6598
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8864 2514 8892 8928
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 8022 9076 8298
rect 9232 8090 9260 8434
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 7002 9076 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6458 9352 6870
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9324 6186 9352 6394
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9416 4593 9444 13126
rect 9508 9450 9536 13874
rect 10152 13530 10180 14418
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9600 12918 9628 13330
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 11014 9720 12786
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12374 9812 12582
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9784 11354 9812 12310
rect 9876 12170 9904 12310
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11898 9904 12106
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10244 11626 10272 12174
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10538 9720 10950
rect 9876 10810 9904 11222
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10152 10742 10180 11494
rect 10244 11150 10272 11562
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9722 9628 9998
rect 10336 9722 10364 12718
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11082 10640 12038
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10612 10810 10640 11018
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10980 9722 11008 17002
rect 11348 16250 11376 27911
rect 11532 27674 11560 39630
rect 11978 39520 12034 39630
rect 12820 39630 13138 39658
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12820 34746 12848 39630
rect 13082 39520 13138 39630
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 14016 39630 14334 39658
rect 12808 34740 12860 34746
rect 12808 34682 12860 34688
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11520 27668 11572 27674
rect 11520 27610 11572 27616
rect 11428 27532 11480 27538
rect 11428 27474 11480 27480
rect 11440 26790 11468 27474
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 11440 26518 11468 26726
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11428 26512 11480 26518
rect 11428 26454 11480 26460
rect 11440 25702 11468 26454
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17270 11744 17682
rect 11704 17264 11756 17270
rect 11532 17224 11704 17252
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11348 16046 11376 16186
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11150 15736 11206 15745
rect 11150 15671 11206 15680
rect 11164 15638 11192 15671
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 15094 11284 15506
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9600 9178 9628 9658
rect 10336 9518 10364 9658
rect 10980 9518 11008 9658
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10692 9444 10744 9450
rect 10744 9404 10824 9432
rect 10692 9386 10744 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 8498 9720 9318
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9508 7002 9536 7822
rect 9600 7546 9628 7958
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9876 7478 9904 8298
rect 10244 8294 10272 9046
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 7818 10272 8230
rect 10428 8022 10456 8842
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6322 9536 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9508 5914 9536 6258
rect 9876 6186 9904 7414
rect 10244 7274 10272 7754
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10428 6934 10456 7958
rect 10520 7886 10548 9318
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8634 10640 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10796 8430 10824 9404
rect 11256 9042 11284 15030
rect 11348 13814 11376 15982
rect 11348 13786 11468 13814
rect 11440 12306 11468 13786
rect 11532 12986 11560 17224
rect 11704 17206 11756 17212
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 16250 11744 16662
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11992 13394 12020 17070
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 15706 12112 16390
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12176 13814 12204 25638
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 13096 17338 13124 23598
rect 13832 22234 13860 39578
rect 14016 32026 14044 39630
rect 14278 39520 14334 39630
rect 15382 39636 15438 40000
rect 15382 39584 15384 39636
rect 15436 39584 15438 39636
rect 15382 39520 15438 39584
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14004 32020 14056 32026
rect 14004 31962 14056 31968
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 15474 24984 15530 24993
rect 15474 24919 15530 24928
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 15488 23866 15516 24919
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 15474 21720 15530 21729
rect 15474 21655 15530 21664
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 15488 20602 15516 21655
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 13634 18320 13690 18329
rect 13634 18255 13690 18264
rect 13648 17338 13676 18255
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16250 12296 16390
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12820 15910 12848 16594
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12636 15162 12664 15506
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12820 15065 12848 15846
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 12806 15056 12862 15065
rect 12806 14991 12862 15000
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 12084 13786 12204 13814
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11440 11558 11468 12242
rect 12084 11665 12112 13786
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 12070 11656 12126 11665
rect 11520 11620 11572 11626
rect 12070 11591 12126 11600
rect 11520 11562 11572 11568
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11440 10674 11468 11222
rect 11532 11150 11560 11562
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8634 11468 8978
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 10784 8424 10836 8430
rect 10782 8392 10784 8401
rect 10836 8392 10838 8401
rect 10782 8327 10838 8336
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10612 7410 10640 8230
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10612 7002 10640 7346
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5370 9812 5646
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9402 4584 9458 4593
rect 9402 4519 9458 4528
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9692 4282 9720 4626
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9876 4154 9904 6122
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10060 5370 10088 5782
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4690 10272 5102
rect 10428 4826 10456 6870
rect 10704 6798 10732 7686
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6458 10732 6734
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5846 10548 6190
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10428 4282 10456 4762
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10796 4154 10824 8327
rect 11532 8106 11560 11086
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10810 11652 10950
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11440 8078 11560 8106
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 5710 11284 6734
rect 11440 6458 11468 8078
rect 12084 7954 12112 11591
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11532 7546 11560 7890
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 12636 6866 12664 11494
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 13910 8528 13966 8537
rect 13910 8463 13966 8472
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 12636 6118 12664 6802
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10980 4282 11008 4626
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 9784 4126 9904 4154
rect 10324 4140 10376 4146
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3670 9168 3878
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 9508 3194 9536 3606
rect 9784 3534 9812 4126
rect 10324 4082 10376 4088
rect 10428 4126 10824 4154
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3738 10180 3946
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9784 3194 9812 3470
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 10060 3058 10088 3470
rect 10336 3466 10364 4082
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10336 2922 10364 3402
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10428 2650 10456 4126
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 12636 3398 12664 6054
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 10796 2378 10824 2926
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11072 2514 11100 2858
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 9784 2009 9812 2246
rect 9770 2000 9826 2009
rect 9770 1935 9826 1944
rect 8942 82 8998 480
rect 8680 54 8998 82
rect 9968 82 9996 2246
rect 10046 82 10102 480
rect 9968 54 10102 82
rect 11072 82 11100 2246
rect 11150 82 11206 480
rect 11072 54 11206 82
rect 6826 0 6882 54
rect 7930 0 7986 54
rect 8942 0 8998 54
rect 10046 0 10102 54
rect 11150 0 11206 54
rect 12162 82 12218 480
rect 12360 82 12388 2790
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 12162 54 12388 82
rect 13266 82 13322 480
rect 13372 82 13400 2314
rect 13924 1737 13952 8463
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14094 2000 14150 2009
rect 14094 1935 14150 1944
rect 13910 1728 13966 1737
rect 13910 1663 13966 1672
rect 13266 54 13400 82
rect 14108 82 14136 1935
rect 14278 82 14334 480
rect 14108 54 14334 82
rect 15120 82 15148 6326
rect 15382 82 15438 480
rect 15120 54 15438 82
rect 12162 0 12218 54
rect 13266 0 13322 54
rect 14278 0 14334 54
rect 15382 0 15438 54
<< via2 >>
rect 1674 37984 1730 38040
rect 1582 29416 1638 29472
rect 1582 23976 1638 24032
rect 2502 35128 2558 35184
rect 2042 21936 2098 21992
rect 1858 20440 1914 20496
rect 1674 18808 1730 18864
rect 110 18536 166 18592
rect 110 7112 166 7168
rect 110 1400 166 1456
rect 1950 20304 2006 20360
rect 1582 15136 1638 15192
rect 2410 19352 2466 19408
rect 3054 24112 3110 24168
rect 2870 21528 2926 21584
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 4250 32272 4306 32328
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 4158 26560 4214 26616
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3146 19080 3202 19136
rect 4250 20576 4306 20632
rect 1582 12280 1638 12336
rect 1582 9424 1638 9480
rect 3054 14320 3110 14376
rect 3974 19896 4030 19952
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3790 19352 3846 19408
rect 3698 18808 3754 18864
rect 4158 19080 4214 19136
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 4526 13776 4582 13832
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3974 10004 3976 10024
rect 3976 10004 4028 10024
rect 4028 10004 4030 10024
rect 3974 9968 4030 10004
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 4342 9968 4398 10024
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4802 13776 4858 13832
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 5906 21528 5962 21584
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6090 20576 6146 20632
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 10046 38256 10102 38312
rect 11058 34992 11114 35048
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 7010 20440 7066 20496
rect 6642 20304 6698 20360
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 7378 15680 7434 15736
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 5630 4664 5686 4720
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 9954 31184 10010 31240
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 9678 24112 9734 24168
rect 10046 21528 10102 21584
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 7470 9968 7526 10024
rect 7470 8472 7526 8528
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 11334 27920 11390 27976
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11150 15680 11206 15736
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 15474 24928 15530 24984
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 15474 21664 15530 21720
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 13634 18264 13690 18320
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 12806 15000 12862 15056
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 12070 11600 12126 11656
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 10782 8372 10784 8392
rect 10784 8372 10836 8392
rect 10836 8372 10838 8392
rect 10782 8336 10838 8372
rect 9402 4528 9458 4584
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 13910 8472 13966 8528
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9770 1944 9826 2000
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14094 1944 14150 2000
rect 13910 1672 13966 1728
<< metal3 >>
rect 0 38496 480 38616
rect 62 38042 122 38496
rect 10041 38314 10107 38317
rect 15520 38314 16000 38344
rect 10041 38312 16000 38314
rect 10041 38256 10046 38312
rect 10102 38256 16000 38312
rect 10041 38254 16000 38256
rect 10041 38251 10107 38254
rect 15520 38224 16000 38254
rect 1669 38042 1735 38045
rect 62 38040 1735 38042
rect 62 37984 1674 38040
rect 1730 37984 1735 38040
rect 62 37982 1735 37984
rect 1669 37979 1735 37982
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 0 35640 480 35760
rect 62 35186 122 35640
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2497 35186 2563 35189
rect 62 35184 2563 35186
rect 62 35128 2502 35184
rect 2558 35128 2563 35184
rect 62 35126 2563 35128
rect 2497 35123 2563 35126
rect 11053 35050 11119 35053
rect 15520 35050 16000 35080
rect 11053 35048 16000 35050
rect 11053 34992 11058 35048
rect 11114 34992 16000 35048
rect 11053 34990 16000 34992
rect 11053 34987 11119 34990
rect 15520 34960 16000 34990
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 0 32784 480 32904
rect 62 32330 122 32784
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 4245 32330 4311 32333
rect 62 32328 4311 32330
rect 62 32272 4250 32328
rect 4306 32272 4311 32328
rect 62 32270 4311 32272
rect 4245 32267 4311 32270
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 15520 31650 16000 31680
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 15518 31560 16000 31650
rect 9949 31242 10015 31245
rect 15518 31242 15578 31560
rect 9949 31240 15578 31242
rect 9949 31184 9954 31240
rect 10010 31184 15578 31240
rect 9949 31182 15578 31184
rect 9949 31179 10015 31182
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 0 29928 480 30048
rect 6277 29952 6597 29953
rect 62 29474 122 29928
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 1577 29474 1643 29477
rect 62 29472 1643 29474
rect 62 29416 1582 29472
rect 1638 29416 1643 29472
rect 62 29414 1643 29416
rect 1577 29411 1643 29414
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 15520 28386 16000 28416
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 15518 28296 16000 28386
rect 11329 27978 11395 27981
rect 15518 27978 15578 28296
rect 11329 27976 15578 27978
rect 11329 27920 11334 27976
rect 11390 27920 15578 27976
rect 11329 27918 15578 27920
rect 11329 27915 11395 27918
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 3610 27232 3930 27233
rect 0 27072 480 27192
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 62 26618 122 27072
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 4153 26618 4219 26621
rect 62 26616 4219 26618
rect 62 26560 4158 26616
rect 4214 26560 4219 26616
rect 62 26558 4219 26560
rect 4153 26555 4219 26558
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 15520 24989 16000 25016
rect 15469 24986 16000 24989
rect 15388 24984 16000 24986
rect 15388 24928 15474 24984
rect 15530 24928 16000 24984
rect 15388 24926 16000 24928
rect 15469 24923 16000 24926
rect 15520 24896 16000 24923
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 0 24216 480 24336
rect 62 24034 122 24216
rect 3049 24170 3115 24173
rect 9673 24170 9739 24173
rect 3049 24168 9739 24170
rect 3049 24112 3054 24168
rect 3110 24112 9678 24168
rect 9734 24112 9739 24168
rect 3049 24110 9739 24112
rect 3049 24107 3115 24110
rect 9673 24107 9739 24110
rect 1577 24034 1643 24037
rect 62 24032 1643 24034
rect 62 23976 1582 24032
rect 1638 23976 1643 24032
rect 62 23974 1643 23976
rect 1577 23971 1643 23974
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 2037 21994 2103 21997
rect 62 21992 2103 21994
rect 62 21936 2042 21992
rect 2098 21936 2103 21992
rect 62 21934 2103 21936
rect 62 21480 122 21934
rect 2037 21931 2103 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 15520 21725 16000 21752
rect 15469 21722 16000 21725
rect 15388 21720 16000 21722
rect 15388 21664 15474 21720
rect 15530 21664 16000 21720
rect 15388 21662 16000 21664
rect 15469 21659 16000 21662
rect 15520 21632 16000 21659
rect 2865 21586 2931 21589
rect 5901 21586 5967 21589
rect 10041 21586 10107 21589
rect 2865 21584 10107 21586
rect 2865 21528 2870 21584
rect 2926 21528 5906 21584
rect 5962 21528 10046 21584
rect 10102 21528 10107 21584
rect 2865 21526 10107 21528
rect 2865 21523 2931 21526
rect 5901 21523 5967 21526
rect 10041 21523 10107 21526
rect 0 21360 480 21480
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 4245 20634 4311 20637
rect 6085 20634 6151 20637
rect 4245 20632 6151 20634
rect 4245 20576 4250 20632
rect 4306 20576 6090 20632
rect 6146 20576 6151 20632
rect 4245 20574 6151 20576
rect 4245 20571 4311 20574
rect 6085 20571 6151 20574
rect 1853 20498 1919 20501
rect 7005 20498 7071 20501
rect 1853 20496 7071 20498
rect 1853 20440 1858 20496
rect 1914 20440 7010 20496
rect 7066 20440 7071 20496
rect 1853 20438 7071 20440
rect 1853 20435 1919 20438
rect 7005 20435 7071 20438
rect 1945 20362 2011 20365
rect 6637 20362 6703 20365
rect 1945 20360 6703 20362
rect 1945 20304 1950 20360
rect 2006 20304 6642 20360
rect 6698 20304 6703 20360
rect 1945 20302 6703 20304
rect 1945 20299 2011 20302
rect 6637 20299 6703 20302
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 3182 19892 3188 19956
rect 3252 19954 3258 19956
rect 3969 19954 4035 19957
rect 3252 19952 4035 19954
rect 3252 19896 3974 19952
rect 4030 19896 4035 19952
rect 3252 19894 4035 19896
rect 3252 19892 3258 19894
rect 3969 19891 4035 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 2405 19410 2471 19413
rect 3785 19410 3851 19413
rect 2405 19408 3851 19410
rect 2405 19352 2410 19408
rect 2466 19352 3790 19408
rect 3846 19352 3851 19408
rect 2405 19350 3851 19352
rect 2405 19347 2471 19350
rect 3785 19347 3851 19350
rect 3141 19138 3207 19141
rect 4153 19138 4219 19141
rect 3141 19136 4219 19138
rect 3141 19080 3146 19136
rect 3202 19080 4158 19136
rect 4214 19080 4219 19136
rect 3141 19078 4219 19080
rect 3141 19075 3207 19078
rect 4153 19075 4219 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 1669 18866 1735 18869
rect 3693 18866 3759 18869
rect 1669 18864 3759 18866
rect 1669 18808 1674 18864
rect 1730 18808 3698 18864
rect 3754 18808 3759 18864
rect 1669 18806 3759 18808
rect 1669 18803 1735 18806
rect 3693 18803 3759 18806
rect 0 18592 480 18624
rect 0 18536 110 18592
rect 166 18536 480 18592
rect 0 18504 480 18536
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 13629 18322 13695 18325
rect 15520 18322 16000 18352
rect 13629 18320 16000 18322
rect 13629 18264 13634 18320
rect 13690 18264 16000 18320
rect 13629 18262 16000 18264
rect 13629 18259 13695 18262
rect 15520 18232 16000 18262
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 6277 15808 6597 15809
rect 0 15648 480 15768
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 7373 15738 7439 15741
rect 11145 15738 11211 15741
rect 7373 15736 11211 15738
rect 7373 15680 7378 15736
rect 7434 15680 11150 15736
rect 11206 15680 11211 15736
rect 7373 15678 11211 15680
rect 7373 15675 7439 15678
rect 11145 15675 11211 15678
rect 62 15194 122 15648
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1577 15194 1643 15197
rect 62 15192 1643 15194
rect 62 15136 1582 15192
rect 1638 15136 1643 15192
rect 62 15134 1643 15136
rect 1577 15131 1643 15134
rect 12801 15058 12867 15061
rect 15520 15058 16000 15088
rect 12801 15056 16000 15058
rect 12801 15000 12806 15056
rect 12862 15000 16000 15056
rect 12801 14998 16000 15000
rect 12801 14995 12867 14998
rect 15520 14968 16000 14998
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3049 14378 3115 14381
rect 3182 14378 3188 14380
rect 3049 14376 3188 14378
rect 3049 14320 3054 14376
rect 3110 14320 3188 14376
rect 3049 14318 3188 14320
rect 3049 14315 3115 14318
rect 3182 14316 3188 14318
rect 3252 14316 3258 14380
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 4521 13834 4587 13837
rect 4797 13834 4863 13837
rect 4521 13832 4863 13834
rect 4521 13776 4526 13832
rect 4582 13776 4802 13832
rect 4858 13776 4863 13832
rect 4521 13774 4863 13776
rect 4521 13771 4587 13774
rect 4797 13771 4863 13774
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12792 480 12912
rect 62 12338 122 12792
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 1577 12338 1643 12341
rect 62 12336 1643 12338
rect 62 12280 1582 12336
rect 1638 12280 1643 12336
rect 62 12278 1643 12280
rect 1577 12275 1643 12278
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 12065 11658 12131 11661
rect 15520 11658 16000 11688
rect 12065 11656 16000 11658
rect 12065 11600 12070 11656
rect 12126 11600 16000 11656
rect 12065 11598 16000 11600
rect 12065 11595 12131 11598
rect 15520 11568 16000 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 0 9936 480 10056
rect 3969 10026 4035 10029
rect 4337 10026 4403 10029
rect 7465 10026 7531 10029
rect 3969 10024 7531 10026
rect 3969 9968 3974 10024
rect 4030 9968 4342 10024
rect 4398 9968 7470 10024
rect 7526 9968 7531 10024
rect 3969 9966 7531 9968
rect 3969 9963 4035 9966
rect 4337 9963 4403 9966
rect 7465 9963 7531 9966
rect 62 9482 122 9936
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 1577 9482 1643 9485
rect 62 9480 1643 9482
rect 62 9424 1582 9480
rect 1638 9424 1643 9480
rect 62 9422 1643 9424
rect 1577 9419 1643 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 7465 8530 7531 8533
rect 13905 8530 13971 8533
rect 7465 8528 13971 8530
rect 7465 8472 7470 8528
rect 7526 8472 13910 8528
rect 13966 8472 13971 8528
rect 7465 8470 13971 8472
rect 7465 8467 7531 8470
rect 13905 8467 13971 8470
rect 10777 8394 10843 8397
rect 15520 8394 16000 8424
rect 10777 8392 16000 8394
rect 10777 8336 10782 8392
rect 10838 8336 16000 8392
rect 10777 8334 16000 8336
rect 10777 8331 10843 8334
rect 15520 8304 16000 8334
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 0 7168 480 7200
rect 0 7112 110 7168
rect 166 7112 480 7168
rect 0 7080 480 7112
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 15520 4994 16000 5024
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 15518 4904 16000 4994
rect 5625 4722 5691 4725
rect 62 4720 5691 4722
rect 62 4664 5630 4720
rect 5686 4664 5691 4720
rect 62 4662 5691 4664
rect 62 4344 122 4662
rect 5625 4659 5691 4662
rect 9397 4586 9463 4589
rect 15518 4586 15578 4904
rect 9397 4584 15578 4586
rect 9397 4528 9402 4584
rect 9458 4528 15578 4584
rect 9397 4526 15578 4528
rect 9397 4523 9463 4526
rect 3610 4384 3930 4385
rect 0 4224 480 4344
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 9765 2002 9831 2005
rect 14089 2002 14155 2005
rect 9765 2000 14155 2002
rect 9765 1944 9770 2000
rect 9826 1944 14094 2000
rect 14150 1944 14155 2000
rect 9765 1942 14155 1944
rect 9765 1939 9831 1942
rect 14089 1939 14155 1942
rect 13905 1730 13971 1733
rect 15520 1730 16000 1760
rect 13905 1728 16000 1730
rect 13905 1672 13910 1728
rect 13966 1672 16000 1728
rect 13905 1670 16000 1672
rect 13905 1667 13971 1670
rect 15520 1640 16000 1670
rect 0 1456 480 1488
rect 0 1400 110 1456
rect 166 1400 480 1456
rect 0 1368 480 1400
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3188 19892 3252 19956
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3188 14316 3252 14380
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3187 19956 3253 19957
rect 3187 19892 3188 19956
rect 3252 19892 3253 19956
rect 3187 19891 3253 19892
rect 3190 14381 3250 19891
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3187 14380 3253 14381
rect 3187 14316 3188 14380
rect 3252 14316 3253 14380
rect 3187 14315 3253 14316
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_nor2_4  _070_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _188_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_70 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_48
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_63
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_69
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_conb_1  _175_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_25
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _172_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_65
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_130
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_38
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_42
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_52
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_124
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_35
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _103_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use scs8hd_or3_4  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_113
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_9
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _150_
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _167_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _147_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _157_
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_buf_1  _063_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 590 592
use scs8hd_or3_4  _161_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_85
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_119
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_121
timestamp 1586364061
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _073_
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_8
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_12
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_39
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_9
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_12
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_16
timestamp 1586364061
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_20
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_24
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_31
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_38
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_100
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_112
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use scs8hd_nor3_4  _143_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_48
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_92
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_103
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_21_115
timestamp 1586364061
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_130
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 406 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 682 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_nor3_4  _144_
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_14
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_37
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_139
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_145
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_48
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_52
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_85
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_113
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_12
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7360 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_102
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_129
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_9
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_46
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_50
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_70
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_82
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_130
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_138
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_142
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 2300 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_63
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_79
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_8  _152_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_or4_4  _135_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_16
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_20
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 130 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_49
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 314 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_10
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_38
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_48
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_52
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_114
timestamp 1586364061
transform 1 0 11592 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_138
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_10
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_9
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_13
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_or3_4  _082_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_8  _126_
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_26
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 866 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_49
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 866 592
use scs8hd_or2_4  _100_
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_87
timestamp 1586364061
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_114
timestamp 1586364061
transform 1 0 11592 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_138
timestamp 1586364061
transform 1 0 13800 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 1472 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_13
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_17
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4876 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_30
timestamp 1586364061
transform 1 0 3864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_60
timestamp 1586364061
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_68
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7728 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_83
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  _119_
timestamp 1586364061
transform 1 0 10488 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_105
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_10
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 4140 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_42
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_50
timestamp 1586364061
transform 1 0 5704 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_67
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_71
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_14
timestamp 1586364061
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_18
timestamp 1586364061
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  FILLER_37_41
timestamp 1586364061
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_79
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_103
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_107
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_119
timestamp 1586364061
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_37
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_48
timestamp 1586364061
transform 1 0 5520 0 -1 23392
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_67
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_88
timestamp 1586364061
transform 1 0 9200 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_114
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_12
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 774 592
use scs8hd_or3_4  _154_
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_23
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_48
timestamp 1586364061
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_52
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_59
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_64
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_73
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_76
timestamp 1586364061
transform 1 0 8096 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_83
timestamp 1586364061
transform 1 0 8740 0 -1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_117
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_138
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 2944 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_19
timestamp 1586364061
transform 1 0 2852 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_35
timestamp 1586364061
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_52
timestamp 1586364061
transform 1 0 5888 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_57
timestamp 1586364061
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_73
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_77
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_84
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_88
timestamp 1586364061
transform 1 0 9200 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_95
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_99
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_103
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_109
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_112
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_120
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 2944 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2392 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_16
timestamp 1586364061
transform 1 0 2576 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_37
timestamp 1586364061
transform 1 0 4508 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_49
timestamp 1586364061
transform 1 0 5612 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_53
timestamp 1586364061
transform 1 0 5980 0 -1 25568
box -38 -48 774 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_72
timestamp 1586364061
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_76
timestamp 1586364061
transform 1 0 8096 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_83
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_102
timestamp 1586364061
transform 1 0 10488 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_113
timestamp 1586364061
transform 1 0 11500 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 590 592
use scs8hd_decap_3  FILLER_43_11
timestamp 1586364061
transform 1 0 2116 0 1 25568
box -38 -48 314 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 3404 0 1 25568
box -38 -48 866 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 2392 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_17
timestamp 1586364061
transform 1 0 2668 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_22
timestamp 1586364061
transform 1 0 3128 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_34
timestamp 1586364061
transform 1 0 4232 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_38
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_56
timestamp 1586364061
transform 1 0 6256 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_60
timestamp 1586364061
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_65
timestamp 1586364061
transform 1 0 7084 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_69
timestamp 1586364061
transform 1 0 7452 0 1 25568
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8096 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_73
timestamp 1586364061
transform 1 0 7820 0 1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_87
timestamp 1586364061
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_91
timestamp 1586364061
transform 1 0 9476 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_104
timestamp 1586364061
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_108
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_43_112
timestamp 1586364061
transform 1 0 11408 0 1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_43_120
timestamp 1586364061
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_6  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_8  FILLER_44_12
timestamp 1586364061
transform 1 0 2208 0 -1 26656
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 3404 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_23
timestamp 1586364061
transform 1 0 3220 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 26656
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_46
timestamp 1586364061
transform 1 0 5336 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_50
timestamp 1586364061
transform 1 0 5704 0 -1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 7084 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_63
timestamp 1586364061
transform 1 0 6900 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_67
timestamp 1586364061
transform 1 0 7268 0 -1 26656
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 26656
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_84
timestamp 1586364061
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_102
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_12  FILLER_44_113
timestamp 1586364061
transform 1 0 11500 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_125
timestamp 1586364061
transform 1 0 12604 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_44_137
timestamp 1586364061
transform 1 0 13708 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 3404 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 3220 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_34
timestamp 1586364061
transform 1 0 4232 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_38
timestamp 1586364061
transform 1 0 4600 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_55
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 6900 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_72
timestamp 1586364061
transform 1 0 7728 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_76
timestamp 1586364061
transform 1 0 8096 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 9476 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_89
timestamp 1586364061
transform 1 0 9292 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_93
timestamp 1586364061
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 10028 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_106
timestamp 1586364061
transform 1 0 10856 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_114
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 774 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 1564 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_7
timestamp 1586364061
transform 1 0 1748 0 1 27744
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2852 0 1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 3404 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_22
timestamp 1586364061
transform 1 0 3128 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_26
timestamp 1586364061
transform 1 0 3496 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_33
timestamp 1586364061
transform 1 0 4140 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_37
timestamp 1586364061
transform 1 0 4508 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_36
timestamp 1586364061
transform 1 0 4416 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 27744
box -38 -48 866 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 4784 0 -1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_49
timestamp 1586364061
transform 1 0 5612 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_53
timestamp 1586364061
transform 1 0 5980 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_4  FILLER_47_50
timestamp 1586364061
transform 1 0 5704 0 1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_47_54
timestamp 1586364061
transform 1 0 6072 0 1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 27744
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_57
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_65
timestamp 1586364061
transform 1 0 7084 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_69
timestamp 1586364061
transform 1 0 7452 0 1 27744
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_76
timestamp 1586364061
transform 1 0 8096 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_81
timestamp 1586364061
transform 1 0 8556 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_73
timestamp 1586364061
transform 1 0 7820 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_87
timestamp 1586364061
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_89
timestamp 1586364061
transform 1 0 9292 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_85
timestamp 1586364061
transform 1 0 8924 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_91
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_8  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_110
timestamp 1586364061
transform 1 0 11224 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_104
timestamp 1586364061
transform 1 0 10672 0 1 27744
box -38 -48 1142 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 11408 0 -1 27744
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_116
timestamp 1586364061
transform 1 0 11776 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_47_116
timestamp 1586364061
transform 1 0 11776 0 1 27744
box -38 -48 590 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_128
timestamp 1586364061
transform 1 0 12880 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_decap_6  FILLER_46_140
timestamp 1586364061
transform 1 0 13984 0 -1 27744
box -38 -48 590 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_7
timestamp 1586364061
transform 1 0 1748 0 -1 28832
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_19
timestamp 1586364061
transform 1 0 2852 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_23
timestamp 1586364061
transform 1 0 3220 0 -1 28832
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 4232 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_36
timestamp 1586364061
transform 1 0 4416 0 -1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6164 0 -1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_47
timestamp 1586364061
transform 1 0 5428 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_51
timestamp 1586364061
transform 1 0 5796 0 -1 28832
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_66
timestamp 1586364061
transform 1 0 7176 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_70
timestamp 1586364061
transform 1 0 7544 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_83
timestamp 1586364061
transform 1 0 8740 0 -1 28832
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_87
timestamp 1586364061
transform 1 0 9108 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_91
timestamp 1586364061
transform 1 0 9476 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_96
timestamp 1586364061
transform 1 0 9936 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_100
timestamp 1586364061
transform 1 0 10304 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_112
timestamp 1586364061
transform 1 0 11408 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_124
timestamp 1586364061
transform 1 0 12512 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_136
timestamp 1586364061
transform 1 0 13616 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_144
timestamp 1586364061
transform 1 0 14352 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_25
timestamp 1586364061
transform 1 0 3404 0 1 28832
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4140 0 1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_29
timestamp 1586364061
transform 1 0 3772 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_44
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 774 592
use scs8hd_decap_4  FILLER_49_54
timestamp 1586364061
transform 1 0 6072 0 1 28832
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_58
timestamp 1586364061
transform 1 0 6440 0 1 28832
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_75
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_88
timestamp 1586364061
transform 1 0 9200 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_92
timestamp 1586364061
transform 1 0 9568 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_95
timestamp 1586364061
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_99
timestamp 1586364061
transform 1 0 10212 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_111
timestamp 1586364061
transform 1 0 11316 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  FILLER_49_119
timestamp 1586364061
transform 1 0 12052 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_41
timestamp 1586364061
transform 1 0 4876 0 -1 29920
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_49
timestamp 1586364061
transform 1 0 5612 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_50_55
timestamp 1586364061
transform 1 0 6164 0 -1 29920
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 29920
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_72
timestamp 1586364061
transform 1 0 7728 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_76
timestamp 1586364061
transform 1 0 8096 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_83
timestamp 1586364061
transform 1 0 8740 0 -1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_87
timestamp 1586364061
transform 1 0 9108 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_91
timestamp 1586364061
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_102
timestamp 1586364061
transform 1 0 10488 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_50_106
timestamp 1586364061
transform 1 0 10856 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_118
timestamp 1586364061
transform 1 0 11960 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_130
timestamp 1586364061
transform 1 0 13064 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_142
timestamp 1586364061
transform 1 0 14168 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4508 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4140 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_31
timestamp 1586364061
transform 1 0 3956 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_35
timestamp 1586364061
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_48
timestamp 1586364061
transform 1 0 5520 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_52
timestamp 1586364061
transform 1 0 5888 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_56
timestamp 1586364061
transform 1 0 6256 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_60
timestamp 1586364061
transform 1 0 6624 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_65
timestamp 1586364061
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_51_69
timestamp 1586364061
transform 1 0 7452 0 1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8280 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_89
timestamp 1586364061
transform 1 0 9292 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_95
timestamp 1586364061
transform 1 0 9844 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_106
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 3312 0 1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 3128 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 3312 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_1  FILLER_52_23
timestamp 1586364061
transform 1 0 3220 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_26
timestamp 1586364061
transform 1 0 3496 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_6  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_21
timestamp 1586364061
transform 1 0 3036 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_33
timestamp 1586364061
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_30
timestamp 1586364061
transform 1 0 3864 0 -1 31008
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_37
timestamp 1586364061
transform 1 0 4508 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_38
timestamp 1586364061
transform 1 0 4600 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 31008
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4876 0 1 31008
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5428 0 -1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_52
timestamp 1586364061
transform 1 0 5888 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_4  FILLER_53_56
timestamp 1586364061
transform 1 0 6256 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_60
timestamp 1586364061
transform 1 0 6624 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_66
timestamp 1586364061
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 31008
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8280 0 1 31008
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_72
timestamp 1586364061
transform 1 0 7728 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_70
timestamp 1586364061
transform 1 0 7544 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_84
timestamp 1586364061
transform 1 0 8832 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_4  FILLER_53_89
timestamp 1586364061
transform 1 0 9292 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_95
timestamp 1586364061
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 11224 0 -1 31008
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 31008
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 11040 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_102
timestamp 1586364061
transform 1 0 10488 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_106
timestamp 1586364061
transform 1 0 10856 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_106
timestamp 1586364061
transform 1 0 10856 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_113
timestamp 1586364061
transform 1 0 11500 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_114
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 774 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_125
timestamp 1586364061
transform 1 0 12604 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_52_137
timestamp 1586364061
transform 1 0 13708 0 -1 31008
box -38 -48 774 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4784 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_29
timestamp 1586364061
transform 1 0 3772 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 32096
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_54_53
timestamp 1586364061
transform 1 0 5980 0 -1 32096
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_70
timestamp 1586364061
transform 1 0 7544 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_74
timestamp 1586364061
transform 1 0 7912 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_78
timestamp 1586364061
transform 1 0 8280 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_81
timestamp 1586364061
transform 1 0 8556 0 -1 32096
box -38 -48 774 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_89
timestamp 1586364061
transform 1 0 9292 0 -1 32096
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_102
timestamp 1586364061
transform 1 0 10488 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_106
timestamp 1586364061
transform 1 0 10856 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_113
timestamp 1586364061
transform 1 0 11500 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_125
timestamp 1586364061
transform 1 0 12604 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_54_137
timestamp 1586364061
transform 1 0 13708 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3404 0 1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_55_23
timestamp 1586364061
transform 1 0 3220 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_36
timestamp 1586364061
transform 1 0 4416 0 1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_42
timestamp 1586364061
transform 1 0 4968 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_53
timestamp 1586364061
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_57
timestamp 1586364061
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 8372 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8188 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_71
timestamp 1586364061
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_75
timestamp 1586364061
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 9936 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_55_88
timestamp 1586364061
transform 1 0 9200 0 1 32096
box -38 -48 590 592
use scs8hd_decap_12  FILLER_55_105
timestamp 1586364061
transform 1 0 10764 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_55_117
timestamp 1586364061
transform 1 0 11868 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_121
timestamp 1586364061
transform 1 0 12236 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 4600 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_6  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_51
timestamp 1586364061
transform 1 0 5796 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_55
timestamp 1586364061
transform 1 0 6164 0 -1 33184
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 6808 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_60
timestamp 1586364061
transform 1 0 6624 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_64
timestamp 1586364061
transform 1 0 6992 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_76
timestamp 1586364061
transform 1 0 8096 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_83
timestamp 1586364061
transform 1 0 8740 0 -1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 9936 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_91
timestamp 1586364061
transform 1 0 9476 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_98
timestamp 1586364061
transform 1 0 10120 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_110
timestamp 1586364061
transform 1 0 11224 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_122
timestamp 1586364061
transform 1 0 12328 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_134
timestamp 1586364061
transform 1 0 13432 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 4600 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 4416 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_35
timestamp 1586364061
transform 1 0 4324 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_47
timestamp 1586364061
transform 1 0 5428 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_53
timestamp 1586364061
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_57
timestamp 1586364061
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8556 0 1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_73
timestamp 1586364061
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_77
timestamp 1586364061
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_92
timestamp 1586364061
transform 1 0 9568 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_96
timestamp 1586364061
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_100
timestamp 1586364061
transform 1 0 10304 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_57_112
timestamp 1586364061
transform 1 0 11408 0 1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_57_120
timestamp 1586364061
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 4784 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 5796 0 -1 34272
box -38 -48 866 592
use scs8hd_decap_8  FILLER_58_43
timestamp 1586364061
transform 1 0 5060 0 -1 34272
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_60
timestamp 1586364061
transform 1 0 6624 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_3  FILLER_58_65
timestamp 1586364061
transform 1 0 7084 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_79
timestamp 1586364061
transform 1 0 8372 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_83
timestamp 1586364061
transform 1 0 8740 0 -1 34272
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_58_91
timestamp 1586364061
transform 1 0 9476 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_102
timestamp 1586364061
transform 1 0 10488 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_114
timestamp 1586364061
transform 1 0 11592 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_126
timestamp 1586364061
transform 1 0 12696 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_58_138
timestamp 1586364061
transform 1 0 13800 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 5612 0 1 34272
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5888 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_53
timestamp 1586364061
transform 1 0 5980 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_60_55
timestamp 1586364061
transform 1 0 6164 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_59
timestamp 1586364061
transform 1 0 6532 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_76
timestamp 1586364061
transform 1 0 8096 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_72
timestamp 1586364061
transform 1 0 7728 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_76
timestamp 1586364061
transform 1 0 8096 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_72
timestamp 1586364061
transform 1 0 7728 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_79
timestamp 1586364061
transform 1 0 8372 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 34272
box -38 -48 222 592
use scs8hd_conb_1  _173_
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_8  FILLER_60_83
timestamp 1586364061
transform 1 0 8740 0 -1 35360
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 34272
box -38 -48 866 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_89
timestamp 1586364061
transform 1 0 9292 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_91
timestamp 1586364061
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 10580 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_101
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_105
timestamp 1586364061
transform 1 0 10764 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_97
timestamp 1586364061
transform 1 0 10028 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_109
timestamp 1586364061
transform 1 0 11132 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_59_117
timestamp 1586364061
transform 1 0 11868 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_121
timestamp 1586364061
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 12972 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_127
timestamp 1586364061
transform 1 0 12788 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_131
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_133
timestamp 1586364061
transform 1 0 13340 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_65
timestamp 1586364061
transform 1 0 7084 0 1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_61_69
timestamp 1586364061
transform 1 0 7452 0 1 35360
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 35360
box -38 -48 314 592
use scs8hd_decap_8  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_97
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_101
timestamp 1586364061
transform 1 0 10396 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_61_113
timestamp 1586364061
transform 1 0 11500 0 1 35360
box -38 -48 774 592
use scs8hd_fill_1  FILLER_61_121
timestamp 1586364061
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 2594 0 2650 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 15520 1640 16000 1760 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 1368 480 1488 6 address[2]
port 2 nsew default input
rlabel metal3 s 15520 4904 16000 5024 6 address[3]
port 3 nsew default input
rlabel metal2 s 570 39520 626 40000 6 address[4]
port 4 nsew default input
rlabel metal2 s 1674 39520 1730 40000 6 address[5]
port 5 nsew default input
rlabel metal2 s 2778 39520 2834 40000 6 address[6]
port 6 nsew default input
rlabel metal3 s 15520 8304 16000 8424 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 3974 39520 4030 40000 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 5078 39520 5134 40000 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal3 s 15520 11568 16000 11688 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 6274 39520 6330 40000 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal3 s 15520 14968 16000 15088 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal3 s 15520 18232 16000 18352 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal3 s 15520 21632 16000 21752 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal3 s 15520 24896 16000 25016 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal3 s 15520 28296 16000 28416 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_top_in[1]
port 26 nsew default input
rlabel metal3 s 0 18504 480 18624 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 7930 0 7986 480 6 chany_top_in[3]
port 28 nsew default input
rlabel metal3 s 15520 31560 16000 31680 6 chany_top_in[4]
port 29 nsew default input
rlabel metal3 s 15520 34960 16000 35080 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal3 s 0 21360 480 21480 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 9678 39520 9734 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 10782 39520 10838 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 11978 39520 12034 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 13082 39520 13138 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal3 s 0 29928 480 30048 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 data_in
port 43 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 44 nsew default input
rlabel metal2 s 12162 0 12218 480 6 left_grid_pin_0_
port 45 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 left_grid_pin_10_
port 46 nsew default tristate
rlabel metal3 s 0 35640 480 35760 6 left_grid_pin_12_
port 47 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 left_grid_pin_14_
port 48 nsew default tristate
rlabel metal3 s 15520 38224 16000 38344 6 left_grid_pin_2_
port 49 nsew default tristate
rlabel metal3 s 0 32784 480 32904 6 left_grid_pin_4_
port 50 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 left_grid_pin_6_
port 51 nsew default tristate
rlabel metal2 s 14278 39520 14334 40000 6 left_grid_pin_8_
port 52 nsew default tristate
rlabel metal2 s 15382 39520 15438 40000 6 right_grid_pin_3_
port 53 nsew default tristate
rlabel metal3 s 0 38496 480 38616 6 right_grid_pin_7_
port 54 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 55 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 56 nsew default input
<< end >>
