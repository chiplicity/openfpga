magic
tech EFS8A
magscale 1 2
timestamp 1602269000
<< locali >>
rect 11103 25313 11138 25347
rect 11253 24735 11287 24769
rect 11253 24701 11414 24735
rect 14841 24667 14875 24837
rect 23063 24225 23098 24259
rect 18003 22117 18048 22151
rect 22511 20961 22546 20995
rect 3341 20383 3375 20553
rect 19435 20009 19441 20043
rect 19435 19941 19469 20009
rect 1443 19873 1478 19907
rect 7757 18887 7791 18921
rect 7665 18853 7791 18887
rect 3709 18615 3743 18785
rect 7475 17833 7481 17867
rect 12167 17833 12173 17867
rect 7475 17765 7509 17833
rect 12167 17765 12201 17833
rect 24075 17697 24110 17731
rect 19251 16983 19285 17051
rect 19251 16949 19257 16983
rect 4439 16745 4445 16779
rect 4439 16677 4473 16745
rect 17267 16609 17302 16643
rect 7107 15657 7113 15691
rect 12811 15657 12817 15691
rect 7107 15589 7141 15657
rect 12811 15589 12845 15657
rect 11287 15521 11322 15555
rect 22419 14909 22454 14943
rect 13829 13855 13863 14025
rect 23811 14025 23949 14059
rect 24823 14025 24961 14059
rect 14105 13855 14139 13957
rect 16405 13855 16439 14025
rect 4019 13345 4110 13379
rect 16031 12631 16065 12699
rect 16031 12597 16037 12631
rect 19251 12393 19257 12427
rect 19251 12325 19285 12393
rect 17819 12257 17854 12291
rect 17693 11611 17727 11781
rect 23765 11543 23799 11849
rect 13363 11305 13369 11339
rect 13363 11237 13397 11305
rect 12023 11169 12058 11203
rect 1443 9469 1570 9503
rect 10051 9129 10057 9163
rect 10051 9061 10085 9129
rect 11471 8993 11506 9027
rect 2881 8279 2915 8585
rect 10603 8041 10609 8075
rect 10603 7973 10637 8041
rect 17693 6171 17727 6341
rect 12115 5729 12150 5763
rect 16899 4641 16934 4675
rect 9321 3995 9355 4233
rect 7067 3961 7205 3995
rect 12265 3995 12299 4233
rect 10149 3553 10310 3587
rect 10149 3383 10183 3553
rect 12391 2941 12518 2975
rect 13093 2839 13127 3009
<< viali >>
rect 10124 25313 10158 25347
rect 11069 25313 11103 25347
rect 13436 25313 13470 25347
rect 14448 25313 14482 25347
rect 10195 25109 10229 25143
rect 11207 25109 11241 25143
rect 12817 25109 12851 25143
rect 13507 25109 13541 25143
rect 14519 25109 14553 25143
rect 15393 24905 15427 24939
rect 10609 24837 10643 24871
rect 14841 24837 14875 24871
rect 11253 24769 11287 24803
rect 12725 24769 12759 24803
rect 8712 24701 8746 24735
rect 9137 24701 9171 24735
rect 9756 24701 9790 24735
rect 10241 24701 10275 24735
rect 11805 24701 11839 24735
rect 13737 24701 13771 24735
rect 14232 24701 14266 24735
rect 15209 24701 15243 24735
rect 15761 24701 15795 24735
rect 11161 24633 11195 24667
rect 12817 24633 12851 24667
rect 13369 24633 13403 24667
rect 14657 24633 14691 24667
rect 14841 24633 14875 24667
rect 8815 24565 8849 24599
rect 9827 24565 9861 24599
rect 11483 24565 11517 24599
rect 12265 24565 12299 24599
rect 14335 24565 14369 24599
rect 15117 24565 15151 24599
rect 11897 24361 11931 24395
rect 14289 24361 14323 24395
rect 15485 24361 15519 24395
rect 17785 24361 17819 24395
rect 24777 24361 24811 24395
rect 12541 24293 12575 24327
rect 12633 24293 12667 24327
rect 6596 24225 6630 24259
rect 7608 24225 7642 24259
rect 8652 24225 8686 24259
rect 10425 24225 10459 24259
rect 14105 24225 14139 24259
rect 15301 24225 15335 24259
rect 15853 24225 15887 24259
rect 16497 24225 16531 24259
rect 17601 24225 17635 24259
rect 23029 24225 23063 24259
rect 24593 24225 24627 24259
rect 10609 24089 10643 24123
rect 13093 24089 13127 24123
rect 16681 24089 16715 24123
rect 6699 24021 6733 24055
rect 7711 24021 7745 24055
rect 8723 24021 8757 24055
rect 10977 24021 11011 24055
rect 12265 24021 12299 24055
rect 23167 24021 23201 24055
rect 5089 23817 5123 23851
rect 7205 23817 7239 23851
rect 8677 23817 8711 23851
rect 10241 23817 10275 23851
rect 10701 23817 10735 23851
rect 16589 23817 16623 23851
rect 18245 23817 18279 23851
rect 21005 23817 21039 23851
rect 24777 23817 24811 23851
rect 25145 23817 25179 23851
rect 7573 23749 7607 23783
rect 13093 23749 13127 23783
rect 13921 23749 13955 23783
rect 15117 23749 15151 23783
rect 22063 23749 22097 23783
rect 22477 23749 22511 23783
rect 9919 23681 9953 23715
rect 12541 23681 12575 23715
rect 14105 23681 14139 23715
rect 14473 23681 14507 23715
rect 23121 23681 23155 23715
rect 1444 23613 1478 23647
rect 1869 23613 1903 23647
rect 4905 23613 4939 23647
rect 5457 23613 5491 23647
rect 7021 23613 7055 23647
rect 8836 23613 8870 23647
rect 9321 23613 9355 23647
rect 9832 23613 9866 23647
rect 10885 23613 10919 23647
rect 11253 23613 11287 23647
rect 15853 23613 15887 23647
rect 16037 23613 16071 23647
rect 18061 23613 18095 23647
rect 20821 23613 20855 23647
rect 21992 23613 22026 23647
rect 24593 23613 24627 23647
rect 1547 23545 1581 23579
rect 6561 23545 6595 23579
rect 11529 23545 11563 23579
rect 12633 23545 12667 23579
rect 13553 23545 13587 23579
rect 14197 23545 14231 23579
rect 15485 23545 15519 23579
rect 3893 23477 3927 23511
rect 6193 23477 6227 23511
rect 8907 23477 8941 23511
rect 11897 23477 11931 23511
rect 12265 23477 12299 23511
rect 15669 23477 15703 23511
rect 17693 23477 17727 23511
rect 18705 23477 18739 23511
rect 21465 23477 21499 23511
rect 24409 23477 24443 23511
rect 5779 23273 5813 23307
rect 9873 23273 9907 23307
rect 12541 23273 12575 23307
rect 14657 23273 14691 23307
rect 4261 23205 4295 23239
rect 11942 23205 11976 23239
rect 13829 23205 13863 23239
rect 15393 23205 15427 23239
rect 15485 23205 15519 23239
rect 4813 23137 4847 23171
rect 5676 23137 5710 23171
rect 6780 23137 6814 23171
rect 8033 23137 8067 23171
rect 8217 23137 8251 23171
rect 10241 23137 10275 23171
rect 10609 23137 10643 23171
rect 13001 23137 13035 23171
rect 17417 23137 17451 23171
rect 17601 23137 17635 23171
rect 18772 23137 18806 23171
rect 4169 23069 4203 23103
rect 8493 23069 8527 23103
rect 8769 23069 8803 23103
rect 10793 23069 10827 23103
rect 11621 23069 11655 23103
rect 13737 23069 13771 23103
rect 15669 23069 15703 23103
rect 17785 23069 17819 23103
rect 6883 23001 6917 23035
rect 14289 23001 14323 23035
rect 2697 22933 2731 22967
rect 7297 22933 7331 22967
rect 7665 22933 7699 22967
rect 11069 22933 11103 22967
rect 15117 22933 15151 22967
rect 18843 22933 18877 22967
rect 19901 22933 19935 22967
rect 1593 22729 1627 22763
rect 3617 22729 3651 22763
rect 3985 22729 4019 22763
rect 4353 22729 4387 22763
rect 5825 22729 5859 22763
rect 11989 22729 12023 22763
rect 15761 22729 15795 22763
rect 17693 22729 17727 22763
rect 18981 22729 19015 22763
rect 21925 22729 21959 22763
rect 24777 22661 24811 22695
rect 2697 22593 2731 22627
rect 6561 22593 6595 22627
rect 6929 22593 6963 22627
rect 8585 22593 8619 22627
rect 10425 22593 10459 22627
rect 10701 22593 10735 22627
rect 13001 22593 13035 22627
rect 14841 22593 14875 22627
rect 19901 22593 19935 22627
rect 20269 22593 20303 22627
rect 1409 22525 1443 22559
rect 10057 22525 10091 22559
rect 13921 22525 13955 22559
rect 14197 22525 14231 22559
rect 16221 22525 16255 22559
rect 16313 22525 16347 22559
rect 16773 22525 16807 22559
rect 18112 22525 18146 22559
rect 21440 22525 21474 22559
rect 24593 22525 24627 22559
rect 25145 22525 25179 22559
rect 2605 22457 2639 22491
rect 3059 22457 3093 22491
rect 4537 22457 4571 22491
rect 4629 22457 4663 22491
rect 5181 22457 5215 22491
rect 6285 22457 6319 22491
rect 7021 22457 7055 22491
rect 7573 22457 7607 22491
rect 8493 22457 8527 22491
rect 8906 22457 8940 22491
rect 10517 22457 10551 22491
rect 13322 22457 13356 22491
rect 14933 22457 14967 22491
rect 15485 22457 15519 22491
rect 18199 22457 18233 22491
rect 19717 22457 19751 22491
rect 19993 22457 20027 22491
rect 1961 22389 1995 22423
rect 5457 22389 5491 22423
rect 7941 22389 7975 22423
rect 9505 22389 9539 22423
rect 11713 22389 11747 22423
rect 12817 22389 12851 22423
rect 14565 22389 14599 22423
rect 16405 22389 16439 22423
rect 17417 22389 17451 22423
rect 18521 22389 18555 22423
rect 21511 22389 21545 22423
rect 2697 22185 2731 22219
rect 4997 22185 5031 22219
rect 6837 22185 6871 22219
rect 9045 22185 9079 22219
rect 11069 22185 11103 22219
rect 12173 22185 12207 22219
rect 14013 22185 14047 22219
rect 15025 22185 15059 22219
rect 19671 22185 19705 22219
rect 4439 22117 4473 22151
rect 6279 22117 6313 22151
rect 8211 22117 8245 22151
rect 9781 22117 9815 22151
rect 9873 22117 9907 22151
rect 11615 22117 11649 22151
rect 13185 22117 13219 22151
rect 17969 22117 18003 22151
rect 21005 22117 21039 22151
rect 21097 22117 21131 22151
rect 2697 22049 2731 22083
rect 2881 22049 2915 22083
rect 3433 22049 3467 22083
rect 5733 22049 5767 22083
rect 8769 22049 8803 22083
rect 15301 22049 15335 22083
rect 15761 22049 15795 22083
rect 16313 22049 16347 22083
rect 17693 22049 17727 22083
rect 19568 22049 19602 22083
rect 4077 21981 4111 22015
rect 5917 21981 5951 22015
rect 7849 21981 7883 22015
rect 10149 21981 10183 22015
rect 11253 21981 11287 22015
rect 12541 21981 12575 22015
rect 13093 21981 13127 22015
rect 15853 21981 15887 22015
rect 21281 21981 21315 22015
rect 13645 21913 13679 21947
rect 2329 21845 2363 21879
rect 3801 21845 3835 21879
rect 7389 21845 7423 21879
rect 10701 21845 10735 21879
rect 12909 21845 12943 21879
rect 18613 21845 18647 21879
rect 19257 21845 19291 21879
rect 2053 21641 2087 21675
rect 4169 21641 4203 21675
rect 8861 21641 8895 21675
rect 12587 21641 12621 21675
rect 13001 21641 13035 21675
rect 17417 21641 17451 21675
rect 20085 21641 20119 21675
rect 22293 21641 22327 21675
rect 22661 21641 22695 21675
rect 14841 21573 14875 21607
rect 20361 21573 20395 21607
rect 3617 21505 3651 21539
rect 5917 21505 5951 21539
rect 6561 21505 6595 21539
rect 7941 21505 7975 21539
rect 9045 21505 9079 21539
rect 9321 21505 9355 21539
rect 11345 21505 11379 21539
rect 11989 21505 12023 21539
rect 14013 21505 14047 21539
rect 15761 21505 15795 21539
rect 18613 21505 18647 21539
rect 19165 21505 19199 21539
rect 21465 21505 21499 21539
rect 2789 21437 2823 21471
rect 2881 21437 2915 21471
rect 3341 21437 3375 21471
rect 5181 21437 5215 21471
rect 5641 21437 5675 21471
rect 7665 21437 7699 21471
rect 7849 21437 7883 21471
rect 8493 21437 8527 21471
rect 10517 21437 10551 21471
rect 10885 21437 10919 21471
rect 11069 21437 11103 21471
rect 12516 21437 12550 21471
rect 15301 21437 15335 21471
rect 18199 21437 18233 21471
rect 20913 21437 20947 21471
rect 21373 21437 21407 21471
rect 21925 21437 21959 21471
rect 4721 21369 4755 21403
rect 7297 21369 7331 21403
rect 9137 21369 9171 21403
rect 10149 21369 10183 21403
rect 13645 21369 13679 21403
rect 13737 21369 13771 21403
rect 15669 21369 15703 21403
rect 16123 21369 16157 21403
rect 17785 21369 17819 21403
rect 19486 21369 19520 21403
rect 1685 21301 1719 21335
rect 2421 21301 2455 21335
rect 4997 21301 5031 21335
rect 6285 21301 6319 21335
rect 11713 21301 11747 21335
rect 13461 21301 13495 21335
rect 16681 21301 16715 21335
rect 18291 21301 18325 21335
rect 19073 21301 19107 21335
rect 20821 21301 20855 21335
rect 2237 21097 2271 21131
rect 7941 21097 7975 21131
rect 9045 21097 9079 21131
rect 9413 21097 9447 21131
rect 14105 21097 14139 21131
rect 15439 21097 15473 21131
rect 15853 21097 15887 21131
rect 21005 21097 21039 21131
rect 24777 21097 24811 21131
rect 1961 21029 1995 21063
rect 5549 21029 5583 21063
rect 6745 21029 6779 21063
rect 7021 21029 7055 21063
rect 7573 21029 7607 21063
rect 9873 21029 9907 21063
rect 13271 21029 13305 21063
rect 16773 21029 16807 21063
rect 18705 21029 18739 21063
rect 1476 20961 1510 20995
rect 2421 20961 2455 20995
rect 2513 20961 2547 20995
rect 2697 20961 2731 20995
rect 4077 20961 4111 20995
rect 4353 20961 4387 20995
rect 4813 20961 4847 20995
rect 5892 20961 5926 20995
rect 8636 20961 8670 20995
rect 11253 20961 11287 20995
rect 11713 20961 11747 20995
rect 13829 20961 13863 20995
rect 15368 20961 15402 20995
rect 21189 20961 21223 20995
rect 21373 20961 21407 20995
rect 22477 20961 22511 20995
rect 22615 20961 22649 20995
rect 24593 20961 24627 20995
rect 2881 20893 2915 20927
rect 3709 20893 3743 20927
rect 6929 20893 6963 20927
rect 8723 20893 8757 20927
rect 9781 20893 9815 20927
rect 10057 20893 10091 20927
rect 11989 20893 12023 20927
rect 12449 20893 12483 20927
rect 12909 20893 12943 20927
rect 16681 20893 16715 20927
rect 16957 20893 16991 20927
rect 18613 20893 18647 20927
rect 18889 20893 18923 20927
rect 4169 20825 4203 20859
rect 5963 20825 5997 20859
rect 1547 20757 1581 20791
rect 5273 20757 5307 20791
rect 6285 20757 6319 20791
rect 16129 20757 16163 20791
rect 20269 20757 20303 20791
rect 1869 20553 1903 20587
rect 3065 20553 3099 20587
rect 3341 20553 3375 20587
rect 3433 20553 3467 20587
rect 4629 20553 4663 20587
rect 7757 20553 7791 20587
rect 8585 20553 8619 20587
rect 9689 20553 9723 20587
rect 9965 20553 9999 20587
rect 10333 20553 10367 20587
rect 15393 20553 15427 20587
rect 17141 20553 17175 20587
rect 17877 20553 17911 20587
rect 18429 20553 18463 20587
rect 19993 20553 20027 20587
rect 24685 20553 24719 20587
rect 2789 20417 2823 20451
rect 11529 20485 11563 20519
rect 19165 20485 19199 20519
rect 5917 20417 5951 20451
rect 6837 20417 6871 20451
rect 10609 20417 10643 20451
rect 10977 20417 11011 20451
rect 12449 20417 12483 20451
rect 14289 20417 14323 20451
rect 14565 20417 14599 20451
rect 16221 20417 16255 20451
rect 16589 20417 16623 20451
rect 18613 20417 18647 20451
rect 19533 20417 19567 20451
rect 20269 20417 20303 20451
rect 21281 20417 21315 20451
rect 21557 20417 21591 20451
rect 2053 20349 2087 20383
rect 2145 20349 2179 20383
rect 2329 20349 2363 20383
rect 3341 20349 3375 20383
rect 3617 20349 3651 20383
rect 3709 20349 3743 20383
rect 3893 20349 3927 20383
rect 4997 20349 5031 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 8309 20349 8343 20383
rect 8769 20349 8803 20383
rect 13369 20349 13403 20383
rect 14013 20349 14047 20383
rect 21741 20349 21775 20383
rect 22201 20349 22235 20383
rect 4353 20281 4387 20315
rect 6653 20281 6687 20315
rect 7199 20281 7233 20315
rect 9131 20281 9165 20315
rect 10701 20281 10735 20315
rect 12770 20281 12804 20315
rect 14381 20281 14415 20315
rect 16313 20281 16347 20315
rect 18705 20281 18739 20315
rect 20361 20281 20395 20315
rect 20913 20281 20947 20315
rect 22753 20281 22787 20315
rect 6285 20213 6319 20247
rect 12265 20213 12299 20247
rect 13645 20213 13679 20247
rect 16037 20213 16071 20247
rect 21833 20213 21867 20247
rect 2053 20009 2087 20043
rect 6193 20009 6227 20043
rect 8861 20009 8895 20043
rect 9413 20009 9447 20043
rect 10793 20009 10827 20043
rect 13093 20009 13127 20043
rect 14059 20009 14093 20043
rect 14381 20009 14415 20043
rect 15117 20009 15151 20043
rect 16405 20009 16439 20043
rect 16773 20009 16807 20043
rect 18613 20009 18647 20043
rect 19441 20009 19475 20043
rect 19993 20009 20027 20043
rect 22569 20009 22603 20043
rect 6698 19941 6732 19975
rect 9873 19941 9907 19975
rect 10425 19941 10459 19975
rect 12494 19941 12528 19975
rect 15847 19941 15881 19975
rect 17417 19941 17451 19975
rect 21097 19941 21131 19975
rect 22017 19941 22051 19975
rect 1409 19873 1443 19907
rect 2421 19873 2455 19907
rect 2697 19873 2731 19907
rect 3157 19873 3191 19907
rect 4077 19873 4111 19907
rect 4353 19873 4387 19907
rect 13988 19873 14022 19907
rect 15485 19873 15519 19907
rect 18981 19873 19015 19907
rect 20269 19873 20303 19907
rect 22477 19873 22511 19907
rect 22937 19873 22971 19907
rect 4169 19805 4203 19839
rect 4813 19805 4847 19839
rect 6377 19805 6411 19839
rect 8217 19805 8251 19839
rect 9781 19805 9815 19839
rect 12173 19805 12207 19839
rect 17325 19805 17359 19839
rect 17601 19805 17635 19839
rect 19073 19805 19107 19839
rect 21005 19805 21039 19839
rect 21281 19805 21315 19839
rect 2513 19737 2547 19771
rect 3617 19737 3651 19771
rect 5549 19737 5583 19771
rect 1547 19669 1581 19703
rect 5181 19669 5215 19703
rect 7297 19669 7331 19703
rect 7573 19669 7607 19703
rect 7941 19669 7975 19703
rect 11253 19669 11287 19703
rect 13369 19669 13403 19703
rect 1777 19465 1811 19499
rect 3249 19465 3283 19499
rect 4997 19465 5031 19499
rect 8401 19465 8435 19499
rect 9781 19465 9815 19499
rect 10057 19465 10091 19499
rect 16681 19465 16715 19499
rect 16911 19465 16945 19499
rect 17601 19465 17635 19499
rect 18291 19465 18325 19499
rect 20269 19465 20303 19499
rect 2329 19397 2363 19431
rect 2881 19397 2915 19431
rect 6469 19397 6503 19431
rect 15945 19397 15979 19431
rect 7113 19329 7147 19363
rect 7389 19329 7423 19363
rect 11805 19329 11839 19363
rect 13185 19329 13219 19363
rect 15025 19329 15059 19363
rect 17233 19329 17267 19363
rect 18613 19329 18647 19363
rect 19349 19329 19383 19363
rect 21189 19329 21223 19363
rect 21465 19329 21499 19363
rect 2513 19261 2547 19295
rect 3433 19261 3467 19295
rect 3525 19261 3559 19295
rect 3709 19261 3743 19295
rect 4445 19261 4479 19295
rect 5457 19261 5491 19295
rect 5641 19261 5675 19295
rect 5917 19261 5951 19295
rect 8585 19261 8619 19295
rect 9045 19261 9079 19295
rect 10793 19261 10827 19295
rect 11253 19261 11287 19295
rect 11529 19261 11563 19295
rect 12541 19261 12575 19295
rect 12909 19261 12943 19295
rect 14080 19261 14114 19295
rect 14841 19261 14875 19295
rect 16840 19261 16874 19295
rect 18220 19261 18254 19295
rect 7205 19193 7239 19227
rect 15387 19193 15421 19227
rect 19670 19193 19704 19227
rect 21281 19193 21315 19227
rect 22845 19193 22879 19227
rect 3893 19125 3927 19159
rect 8033 19125 8067 19159
rect 8677 19125 8711 19159
rect 10701 19125 10735 19159
rect 12173 19125 12207 19159
rect 14151 19125 14185 19159
rect 14473 19125 14507 19159
rect 16313 19125 16347 19159
rect 19257 19125 19291 19159
rect 20545 19125 20579 19159
rect 21005 19125 21039 19159
rect 22109 19125 22143 19159
rect 22477 19125 22511 19159
rect 23673 19125 23707 19159
rect 5825 18921 5859 18955
rect 6377 18921 6411 18955
rect 7757 18921 7791 18955
rect 8401 18921 8435 18955
rect 9413 18921 9447 18955
rect 12817 18921 12851 18955
rect 15485 18921 15519 18955
rect 18981 18921 19015 18955
rect 19993 18921 20027 18955
rect 20637 18921 20671 18955
rect 3893 18853 3927 18887
rect 7113 18853 7147 18887
rect 11615 18853 11649 18887
rect 12541 18853 12575 18887
rect 13185 18853 13219 18887
rect 13737 18853 13771 18887
rect 15853 18853 15887 18887
rect 17417 18853 17451 18887
rect 19394 18853 19428 18887
rect 21097 18853 21131 18887
rect 21925 18853 21959 18887
rect 2421 18785 2455 18819
rect 2513 18785 2547 18819
rect 2697 18785 2731 18819
rect 3709 18785 3743 18819
rect 4169 18785 4203 18819
rect 5641 18785 5675 18819
rect 8620 18785 8654 18819
rect 9781 18785 9815 18819
rect 10149 18785 10183 18819
rect 22477 18785 22511 18819
rect 22937 18785 22971 18819
rect 24108 18785 24142 18819
rect 1409 18717 1443 18751
rect 2881 18717 2915 18751
rect 2329 18649 2363 18683
rect 4077 18717 4111 18751
rect 7021 18717 7055 18751
rect 10425 18717 10459 18751
rect 11253 18717 11287 18751
rect 13093 18717 13127 18751
rect 15117 18717 15151 18751
rect 15761 18717 15795 18751
rect 16221 18717 16255 18751
rect 17325 18717 17359 18751
rect 17601 18717 17635 18751
rect 19073 18717 19107 18751
rect 21005 18717 21039 18751
rect 21373 18717 21407 18751
rect 23029 18717 23063 18751
rect 1961 18581 1995 18615
rect 3433 18581 3467 18615
rect 3709 18581 3743 18615
rect 5181 18581 5215 18615
rect 6745 18581 6779 18615
rect 8033 18581 8067 18615
rect 8723 18581 8757 18615
rect 9045 18581 9079 18615
rect 10793 18581 10827 18615
rect 12173 18581 12207 18615
rect 24179 18581 24213 18615
rect 1685 18377 1719 18411
rect 2605 18377 2639 18411
rect 3249 18377 3283 18411
rect 7849 18377 7883 18411
rect 9413 18377 9447 18411
rect 11621 18377 11655 18411
rect 13461 18377 13495 18411
rect 13921 18377 13955 18411
rect 14933 18377 14967 18411
rect 16313 18377 16347 18411
rect 16773 18377 16807 18411
rect 17693 18377 17727 18411
rect 20177 18377 20211 18411
rect 24593 18377 24627 18411
rect 2053 18309 2087 18343
rect 16037 18309 16071 18343
rect 22477 18309 22511 18343
rect 8493 18241 8527 18275
rect 10057 18241 10091 18275
rect 12530 18241 12564 18275
rect 19257 18241 19291 18275
rect 24225 18241 24259 18275
rect 2237 18173 2271 18207
rect 6837 18173 6871 18207
rect 7297 18173 7331 18207
rect 13185 18173 13219 18207
rect 14064 18173 14098 18207
rect 15117 18173 15151 18207
rect 16916 18173 16950 18207
rect 18280 18173 18314 18207
rect 18705 18173 18739 18207
rect 23708 18173 23742 18207
rect 24720 18173 24754 18207
rect 25145 18173 25179 18207
rect 4077 18105 4111 18139
rect 4169 18105 4203 18139
rect 4721 18105 4755 18139
rect 8309 18105 8343 18139
rect 8585 18105 8619 18139
rect 9137 18105 9171 18139
rect 10149 18105 10183 18139
rect 10701 18105 10735 18139
rect 12265 18105 12299 18139
rect 12633 18105 12667 18139
rect 15438 18105 15472 18139
rect 17003 18105 17037 18139
rect 18383 18105 18417 18139
rect 19619 18105 19653 18139
rect 20453 18105 20487 18139
rect 21189 18105 21223 18139
rect 21281 18105 21315 18139
rect 21833 18105 21867 18139
rect 3801 18037 3835 18071
rect 4997 18037 5031 18071
rect 5365 18037 5399 18071
rect 5549 18037 5583 18071
rect 6101 18037 6135 18071
rect 6561 18037 6595 18071
rect 7113 18037 7147 18071
rect 9781 18037 9815 18071
rect 11345 18037 11379 18071
rect 14151 18037 14185 18071
rect 14473 18037 14507 18071
rect 17417 18037 17451 18071
rect 19165 18037 19199 18071
rect 21005 18037 21039 18071
rect 22201 18037 22235 18071
rect 22845 18037 22879 18071
rect 23811 18037 23845 18071
rect 24823 18037 24857 18071
rect 1547 17833 1581 17867
rect 4997 17833 5031 17867
rect 6009 17833 6043 17867
rect 7481 17833 7515 17867
rect 10701 17833 10735 17867
rect 12173 17833 12207 17867
rect 12725 17833 12759 17867
rect 19073 17833 19107 17867
rect 20637 17833 20671 17867
rect 21097 17833 21131 17867
rect 3433 17765 3467 17799
rect 3801 17765 3835 17799
rect 4439 17765 4473 17799
rect 9873 17765 9907 17799
rect 13001 17765 13035 17799
rect 13461 17765 13495 17799
rect 13634 17765 13668 17799
rect 13746 17765 13780 17799
rect 14289 17765 14323 17799
rect 16037 17765 16071 17799
rect 18889 17765 18923 17799
rect 20085 17765 20119 17799
rect 21649 17765 21683 17799
rect 1476 17697 1510 17731
rect 2697 17697 2731 17731
rect 2881 17697 2915 17731
rect 5825 17697 5859 17731
rect 6561 17697 6595 17731
rect 7113 17697 7147 17731
rect 9413 17697 9447 17731
rect 17417 17697 17451 17731
rect 17877 17697 17911 17731
rect 18981 17697 19015 17731
rect 19533 17697 19567 17731
rect 23064 17697 23098 17731
rect 24041 17697 24075 17731
rect 3157 17629 3191 17663
rect 4077 17629 4111 17663
rect 5641 17629 5675 17663
rect 9781 17629 9815 17663
rect 10425 17629 10459 17663
rect 11805 17629 11839 17663
rect 15945 17629 15979 17663
rect 17969 17629 18003 17663
rect 21557 17629 21591 17663
rect 5273 17561 5307 17595
rect 8309 17561 8343 17595
rect 15577 17561 15611 17595
rect 16497 17561 16531 17595
rect 16865 17561 16899 17595
rect 17325 17561 17359 17595
rect 22109 17561 22143 17595
rect 1869 17493 1903 17527
rect 2237 17493 2271 17527
rect 6837 17493 6871 17527
rect 8033 17493 8067 17527
rect 8769 17493 8803 17527
rect 14565 17493 14599 17527
rect 15025 17493 15059 17527
rect 23167 17493 23201 17527
rect 24179 17493 24213 17527
rect 4353 17289 4387 17323
rect 7941 17289 7975 17323
rect 8585 17289 8619 17323
rect 11529 17289 11563 17323
rect 13645 17289 13679 17323
rect 15945 17289 15979 17323
rect 17417 17289 17451 17323
rect 18337 17289 18371 17323
rect 22523 17289 22557 17323
rect 4997 17221 5031 17255
rect 13093 17221 13127 17255
rect 17785 17221 17819 17255
rect 22293 17221 22327 17255
rect 24501 17221 24535 17255
rect 1685 17153 1719 17187
rect 5273 17153 5307 17187
rect 5917 17153 5951 17187
rect 8861 17153 8895 17187
rect 9137 17153 9171 17187
rect 10425 17153 10459 17187
rect 10701 17153 10735 17187
rect 12541 17153 12575 17187
rect 16589 17153 16623 17187
rect 18889 17153 18923 17187
rect 20177 17153 20211 17187
rect 1961 17085 1995 17119
rect 2329 17085 2363 17119
rect 2605 17085 2639 17119
rect 3433 17085 3467 17119
rect 7021 17085 7055 17119
rect 8217 17085 8251 17119
rect 14473 17085 14507 17119
rect 14749 17085 14783 17119
rect 15025 17085 15059 17119
rect 22420 17085 22454 17119
rect 23740 17085 23774 17119
rect 24133 17085 24167 17119
rect 3341 17017 3375 17051
rect 3795 17017 3829 17051
rect 5365 17017 5399 17051
rect 7342 17017 7376 17051
rect 8953 17017 8987 17051
rect 10517 17017 10551 17051
rect 12265 17017 12299 17051
rect 12633 17017 12667 17051
rect 16221 17017 16255 17051
rect 16313 17017 16347 17051
rect 20913 17017 20947 17051
rect 21005 17017 21039 17051
rect 21557 17017 21591 17051
rect 2973 16949 3007 16983
rect 4721 16949 4755 16983
rect 6285 16949 6319 16983
rect 6653 16949 6687 16983
rect 9781 16949 9815 16983
rect 10149 16949 10183 16983
rect 11897 16949 11931 16983
rect 14013 16949 14047 16983
rect 14841 16949 14875 16983
rect 18797 16949 18831 16983
rect 19257 16949 19291 16983
rect 19809 16949 19843 16983
rect 20637 16949 20671 16983
rect 21833 16949 21867 16983
rect 23029 16949 23063 16983
rect 23811 16949 23845 16983
rect 4445 16745 4479 16779
rect 5365 16745 5399 16779
rect 7757 16745 7791 16779
rect 9413 16745 9447 16779
rect 10701 16745 10735 16779
rect 15025 16745 15059 16779
rect 16405 16745 16439 16779
rect 16681 16745 16715 16779
rect 18061 16745 18095 16779
rect 19257 16745 19291 16779
rect 21925 16745 21959 16779
rect 24133 16745 24167 16779
rect 9781 16677 9815 16711
rect 9873 16677 9907 16711
rect 13829 16677 13863 16711
rect 14381 16677 14415 16711
rect 15847 16677 15881 16711
rect 18699 16677 18733 16711
rect 19625 16677 19659 16711
rect 21097 16677 21131 16711
rect 22569 16677 22603 16711
rect 22661 16677 22695 16711
rect 1476 16609 1510 16643
rect 2697 16609 2731 16643
rect 2973 16609 3007 16643
rect 3157 16609 3191 16643
rect 4077 16609 4111 16643
rect 6009 16609 6043 16643
rect 6377 16609 6411 16643
rect 7665 16609 7699 16643
rect 8033 16609 8067 16643
rect 12081 16609 12115 16643
rect 12633 16609 12667 16643
rect 15485 16609 15519 16643
rect 17233 16609 17267 16643
rect 24225 16609 24259 16643
rect 24501 16609 24535 16643
rect 1961 16541 1995 16575
rect 3893 16541 3927 16575
rect 6653 16541 6687 16575
rect 10425 16541 10459 16575
rect 12725 16541 12759 16575
rect 13737 16541 13771 16575
rect 17785 16541 17819 16575
rect 18337 16541 18371 16575
rect 20994 16541 21028 16575
rect 21649 16541 21683 16575
rect 22845 16541 22879 16575
rect 1547 16473 1581 16507
rect 4997 16473 5031 16507
rect 5641 16473 5675 16507
rect 2329 16405 2363 16439
rect 3433 16405 3467 16439
rect 7113 16405 7147 16439
rect 8677 16405 8711 16439
rect 8953 16405 8987 16439
rect 13369 16405 13403 16439
rect 17371 16405 17405 16439
rect 20729 16405 20763 16439
rect 2145 16201 2179 16235
rect 2605 16201 2639 16235
rect 4169 16201 4203 16235
rect 9781 16201 9815 16235
rect 12081 16201 12115 16235
rect 12633 16201 12667 16235
rect 14749 16201 14783 16235
rect 16129 16201 16163 16235
rect 17233 16201 17267 16235
rect 20545 16201 20579 16235
rect 24823 16201 24857 16235
rect 6009 16133 6043 16167
rect 7757 16133 7791 16167
rect 16497 16133 16531 16167
rect 20821 16133 20855 16167
rect 22477 16133 22511 16167
rect 22845 16133 22879 16167
rect 24501 16133 24535 16167
rect 9137 16065 9171 16099
rect 13185 16065 13219 16099
rect 14289 16065 14323 16099
rect 16727 16065 16761 16099
rect 19625 16065 19659 16099
rect 21465 16065 21499 16099
rect 1409 15997 1443 16031
rect 2881 15997 2915 16031
rect 6837 15997 6871 16031
rect 8125 15997 8159 16031
rect 14841 15997 14875 16031
rect 16640 15997 16674 16031
rect 17785 15997 17819 16031
rect 18337 15997 18371 16031
rect 18521 15997 18555 16031
rect 23724 15997 23758 16031
rect 24133 15997 24167 16031
rect 24720 15997 24754 16031
rect 25145 15997 25179 16031
rect 3433 15929 3467 15963
rect 4629 15929 4663 15963
rect 4721 15929 4755 15963
rect 5273 15929 5307 15963
rect 7158 15929 7192 15963
rect 8677 15929 8711 15963
rect 8769 15929 8803 15963
rect 10241 15929 10275 15963
rect 10333 15929 10367 15963
rect 10885 15929 10919 15963
rect 13369 15929 13403 15963
rect 13461 15929 13495 15963
rect 14013 15929 14047 15963
rect 15203 15929 15237 15963
rect 19946 15929 19980 15963
rect 21557 15929 21591 15963
rect 22109 15929 22143 15963
rect 23811 15929 23845 15963
rect 1593 15861 1627 15895
rect 3709 15861 3743 15895
rect 5641 15861 5675 15895
rect 6653 15861 6687 15895
rect 8401 15861 8435 15895
rect 11161 15861 11195 15895
rect 15761 15861 15795 15895
rect 18153 15861 18187 15895
rect 19165 15861 19199 15895
rect 19533 15861 19567 15895
rect 21281 15861 21315 15895
rect 4261 15657 4295 15691
rect 7113 15657 7147 15691
rect 7665 15657 7699 15691
rect 12817 15657 12851 15691
rect 13369 15657 13403 15691
rect 13737 15657 13771 15691
rect 14335 15657 14369 15691
rect 14933 15657 14967 15691
rect 17233 15657 17267 15691
rect 19625 15657 19659 15691
rect 22017 15657 22051 15691
rect 24133 15657 24167 15691
rect 24777 15657 24811 15691
rect 3157 15589 3191 15623
rect 7941 15589 7975 15623
rect 9505 15589 9539 15623
rect 9873 15589 9907 15623
rect 15761 15589 15795 15623
rect 19067 15589 19101 15623
rect 20729 15589 20763 15623
rect 21097 15589 21131 15623
rect 22569 15589 22603 15623
rect 22661 15589 22695 15623
rect 1476 15521 1510 15555
rect 2421 15521 2455 15555
rect 4077 15521 4111 15555
rect 5181 15521 5215 15555
rect 5733 15521 5767 15555
rect 6285 15521 6319 15555
rect 6653 15521 6687 15555
rect 8620 15521 8654 15555
rect 11253 15521 11287 15555
rect 12449 15521 12483 15555
rect 14264 15521 14298 15555
rect 17233 15521 17267 15555
rect 17693 15521 17727 15555
rect 24593 15521 24627 15555
rect 1961 15453 1995 15487
rect 2789 15453 2823 15487
rect 5917 15453 5951 15487
rect 6745 15453 6779 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 15669 15453 15703 15487
rect 18705 15453 18739 15487
rect 21005 15453 21039 15487
rect 22845 15453 22879 15487
rect 1547 15385 1581 15419
rect 16221 15385 16255 15419
rect 21557 15385 21591 15419
rect 2329 15317 2363 15351
rect 2559 15317 2593 15351
rect 2697 15317 2731 15351
rect 3433 15317 3467 15351
rect 3893 15317 3927 15351
rect 4629 15317 4663 15351
rect 5089 15317 5123 15351
rect 8309 15317 8343 15351
rect 8723 15317 8757 15351
rect 9137 15317 9171 15351
rect 10701 15317 10735 15351
rect 11069 15317 11103 15351
rect 11391 15317 11425 15351
rect 18521 15317 18555 15351
rect 19901 15317 19935 15351
rect 1685 15113 1719 15147
rect 2053 15113 2087 15147
rect 2789 15113 2823 15147
rect 3617 15113 3651 15147
rect 8125 15113 8159 15147
rect 10057 15113 10091 15147
rect 12265 15113 12299 15147
rect 13093 15113 13127 15147
rect 14289 15113 14323 15147
rect 17141 15113 17175 15147
rect 17601 15113 17635 15147
rect 18337 15113 18371 15147
rect 20729 15113 20763 15147
rect 21833 15113 21867 15147
rect 22523 15113 22557 15147
rect 23213 15113 23247 15147
rect 2421 15045 2455 15079
rect 3138 15045 3172 15079
rect 7849 15045 7883 15079
rect 10425 15045 10459 15079
rect 16681 15045 16715 15079
rect 22845 15045 22879 15079
rect 1777 14977 1811 15011
rect 3341 14977 3375 15011
rect 3985 14977 4019 15011
rect 5917 14977 5951 15011
rect 6929 14977 6963 15011
rect 9781 14977 9815 15011
rect 10977 14977 11011 15011
rect 11621 14977 11655 15011
rect 15945 14977 15979 15011
rect 19165 14977 19199 15011
rect 20361 14977 20395 15011
rect 22293 14977 22327 15011
rect 1556 14909 1590 14943
rect 3203 14909 3237 14943
rect 5181 14909 5215 14943
rect 5733 14909 5767 14943
rect 13185 14909 13219 14943
rect 13645 14909 13679 14943
rect 18429 14909 18463 14943
rect 18889 14909 18923 14943
rect 22385 14909 22419 14943
rect 23708 14909 23742 14943
rect 24133 14909 24167 14943
rect 1409 14841 1443 14875
rect 2972 14841 3006 14875
rect 7291 14841 7325 14875
rect 9137 14841 9171 14875
rect 9229 14841 9263 14875
rect 10701 14841 10735 14875
rect 10793 14841 10827 14875
rect 14749 14841 14783 14875
rect 15669 14841 15703 14875
rect 15761 14841 15795 14875
rect 19809 14841 19843 14875
rect 20913 14841 20947 14875
rect 21005 14841 21039 14875
rect 21557 14841 21591 14875
rect 4353 14773 4387 14807
rect 4721 14773 4755 14807
rect 6285 14773 6319 14807
rect 6561 14773 6595 14807
rect 8585 14773 8619 14807
rect 12725 14773 12759 14807
rect 13461 14773 13495 14807
rect 15117 14773 15151 14807
rect 15485 14773 15519 14807
rect 19533 14773 19567 14807
rect 23811 14773 23845 14807
rect 24593 14773 24627 14807
rect 1869 14569 1903 14603
rect 2237 14569 2271 14603
rect 3065 14569 3099 14603
rect 5181 14569 5215 14603
rect 5825 14569 5859 14603
rect 9505 14569 9539 14603
rect 10793 14569 10827 14603
rect 11069 14569 11103 14603
rect 16957 14569 16991 14603
rect 18705 14569 18739 14603
rect 20729 14569 20763 14603
rect 1547 14501 1581 14535
rect 7158 14501 7192 14535
rect 8493 14501 8527 14535
rect 9873 14501 9907 14535
rect 10425 14501 10459 14535
rect 11805 14501 11839 14535
rect 13823 14501 13857 14535
rect 15485 14501 15519 14535
rect 21097 14501 21131 14535
rect 21649 14501 21683 14535
rect 23627 14501 23661 14535
rect 1460 14433 1494 14467
rect 2421 14433 2455 14467
rect 3525 14433 3559 14467
rect 4077 14433 4111 14467
rect 4813 14433 4847 14467
rect 5641 14433 5675 14467
rect 6837 14433 6871 14467
rect 8033 14433 8067 14467
rect 8652 14433 8686 14467
rect 11989 14433 12023 14467
rect 12357 14433 12391 14467
rect 13185 14433 13219 14467
rect 13461 14433 13495 14467
rect 17141 14433 17175 14467
rect 17325 14433 17359 14467
rect 18429 14433 18463 14467
rect 18889 14433 18923 14467
rect 22544 14433 22578 14467
rect 23540 14433 23574 14467
rect 2789 14365 2823 14399
rect 4445 14365 4479 14399
rect 6285 14365 6319 14399
rect 9781 14365 9815 14399
rect 12449 14365 12483 14399
rect 15393 14365 15427 14399
rect 16037 14365 16071 14399
rect 21005 14365 21039 14399
rect 2586 14297 2620 14331
rect 4353 14297 4387 14331
rect 7757 14297 7791 14331
rect 9045 14297 9079 14331
rect 22615 14297 22649 14331
rect 2697 14229 2731 14263
rect 3893 14229 3927 14263
rect 4242 14229 4276 14263
rect 6561 14229 6595 14263
rect 8723 14229 8757 14263
rect 14381 14229 14415 14263
rect 19717 14229 19751 14263
rect 2605 14025 2639 14059
rect 2881 14025 2915 14059
rect 3230 14025 3264 14059
rect 7849 14025 7883 14059
rect 8677 14025 8711 14059
rect 10057 14025 10091 14059
rect 11989 14025 12023 14059
rect 13829 14025 13863 14059
rect 3341 13957 3375 13991
rect 6009 13957 6043 13991
rect 3433 13889 3467 13923
rect 4169 13889 4203 13923
rect 7573 13889 7607 13923
rect 9137 13889 9171 13923
rect 12725 13889 12759 13923
rect 16405 14025 16439 14059
rect 16589 14025 16623 14059
rect 17785 14025 17819 14059
rect 19073 14025 19107 14059
rect 20545 14025 20579 14059
rect 22385 14025 22419 14059
rect 23949 14025 23983 14059
rect 24961 14025 24995 14059
rect 14105 13957 14139 13991
rect 14289 13889 14323 13923
rect 15301 13889 15335 13923
rect 16865 13957 16899 13991
rect 24501 13957 24535 13991
rect 17233 13889 17267 13923
rect 19625 13889 19659 13923
rect 25145 13889 25179 13923
rect 2145 13821 2179 13855
rect 5181 13821 5215 13855
rect 5457 13821 5491 13855
rect 7113 13821 7147 13855
rect 7389 13821 7423 13855
rect 8217 13821 8251 13855
rect 13829 13821 13863 13855
rect 14013 13821 14047 13855
rect 14105 13821 14139 13855
rect 15209 13821 15243 13855
rect 16405 13821 16439 13855
rect 18061 13821 18095 13855
rect 18613 13821 18647 13855
rect 21189 13821 21223 13855
rect 21465 13821 21499 13855
rect 21925 13821 21959 13855
rect 23708 13821 23742 13855
rect 24720 13821 24754 13855
rect 2237 13753 2271 13787
rect 3065 13753 3099 13787
rect 3801 13753 3835 13787
rect 5641 13753 5675 13787
rect 9229 13753 9263 13787
rect 9781 13753 9815 13787
rect 10701 13753 10735 13787
rect 10793 13753 10827 13787
rect 11345 13753 11379 13787
rect 13046 13753 13080 13787
rect 14841 13753 14875 13787
rect 15663 13753 15697 13787
rect 19946 13753 19980 13787
rect 22753 13753 22787 13787
rect 4537 13685 4571 13719
rect 6561 13685 6595 13719
rect 10517 13685 10551 13719
rect 13645 13685 13679 13719
rect 16221 13685 16255 13719
rect 18337 13685 18371 13719
rect 19441 13685 19475 13719
rect 20821 13685 20855 13719
rect 21465 13685 21499 13719
rect 24133 13685 24167 13719
rect 1547 13481 1581 13515
rect 1961 13481 1995 13515
rect 2237 13481 2271 13515
rect 3525 13481 3559 13515
rect 6561 13481 6595 13515
rect 9413 13481 9447 13515
rect 10701 13481 10735 13515
rect 12817 13481 12851 13515
rect 14197 13481 14231 13515
rect 15117 13481 15151 13515
rect 20729 13481 20763 13515
rect 22569 13481 22603 13515
rect 24777 13481 24811 13515
rect 6003 13413 6037 13447
rect 7573 13413 7607 13447
rect 10102 13413 10136 13447
rect 11713 13413 11747 13447
rect 13369 13413 13403 13447
rect 15485 13413 15519 13447
rect 17049 13413 17083 13447
rect 19394 13413 19428 13447
rect 1476 13345 1510 13379
rect 2421 13345 2455 13379
rect 3985 13345 4019 13379
rect 6837 13345 6871 13379
rect 10977 13345 11011 13379
rect 17601 13345 17635 13379
rect 20913 13345 20947 13379
rect 21373 13345 21407 13379
rect 22477 13345 22511 13379
rect 23029 13345 23063 13379
rect 24593 13345 24627 13379
rect 2789 13277 2823 13311
rect 4445 13277 4479 13311
rect 5641 13277 5675 13311
rect 7481 13277 7515 13311
rect 9781 13277 9815 13311
rect 11621 13277 11655 13311
rect 11897 13277 11931 13311
rect 13277 13277 13311 13311
rect 13921 13277 13955 13311
rect 15393 13277 15427 13311
rect 16957 13277 16991 13311
rect 18981 13277 19015 13311
rect 19073 13277 19107 13311
rect 21465 13277 21499 13311
rect 2697 13209 2731 13243
rect 4353 13209 4387 13243
rect 5089 13209 5123 13243
rect 8033 13209 8067 13243
rect 15945 13209 15979 13243
rect 19993 13209 20027 13243
rect 2559 13141 2593 13175
rect 3065 13141 3099 13175
rect 3801 13141 3835 13175
rect 4215 13141 4249 13175
rect 4721 13141 4755 13175
rect 5457 13141 5491 13175
rect 7297 13141 7331 13175
rect 8401 13141 8435 13175
rect 9137 13141 9171 13175
rect 18061 13141 18095 13175
rect 18429 13141 18463 13175
rect 21925 13141 21959 13175
rect 2881 12937 2915 12971
rect 3341 12937 3375 12971
rect 4169 12937 4203 12971
rect 4537 12937 4571 12971
rect 6285 12937 6319 12971
rect 7757 12937 7791 12971
rect 11069 12937 11103 12971
rect 12173 12937 12207 12971
rect 15209 12937 15243 12971
rect 15577 12937 15611 12971
rect 16957 12937 16991 12971
rect 20913 12937 20947 12971
rect 22201 12937 22235 12971
rect 22937 12937 22971 12971
rect 3203 12869 3237 12903
rect 4813 12869 4847 12903
rect 6561 12869 6595 12903
rect 10701 12869 10735 12903
rect 11437 12869 11471 12903
rect 3433 12801 3467 12835
rect 9045 12801 9079 12835
rect 9505 12801 9539 12835
rect 13001 12801 13035 12835
rect 17233 12801 17267 12835
rect 21557 12801 21591 12835
rect 1869 12733 1903 12767
rect 5181 12733 5215 12767
rect 5733 12733 5767 12767
rect 6980 12733 7014 12767
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 14013 12733 14047 12767
rect 14197 12733 14231 12767
rect 14565 12733 14599 12767
rect 14841 12733 14875 12767
rect 15669 12733 15703 12767
rect 18096 12733 18130 12767
rect 18521 12733 18555 12767
rect 19349 12733 19383 12767
rect 3065 12665 3099 12699
rect 3801 12665 3835 12699
rect 5917 12665 5951 12699
rect 7067 12665 7101 12699
rect 8033 12665 8067 12699
rect 8125 12665 8159 12699
rect 8677 12665 8711 12699
rect 10149 12665 10183 12699
rect 10241 12665 10275 12699
rect 18199 12665 18233 12699
rect 19670 12665 19704 12699
rect 20545 12665 20579 12699
rect 21189 12665 21223 12699
rect 21281 12665 21315 12699
rect 1685 12597 1719 12631
rect 2421 12597 2455 12631
rect 7481 12597 7515 12631
rect 9781 12597 9815 12631
rect 11897 12597 11931 12631
rect 13553 12597 13587 12631
rect 16037 12597 16071 12631
rect 16589 12597 16623 12631
rect 19165 12597 19199 12631
rect 20269 12597 20303 12631
rect 22477 12597 22511 12631
rect 23673 12597 23707 12631
rect 24593 12597 24627 12631
rect 4629 12393 4663 12427
rect 7849 12393 7883 12427
rect 8493 12393 8527 12427
rect 9045 12393 9079 12427
rect 13645 12393 13679 12427
rect 15669 12393 15703 12427
rect 19257 12393 19291 12427
rect 19809 12393 19843 12427
rect 21925 12393 21959 12427
rect 1409 12325 1443 12359
rect 4307 12325 4341 12359
rect 5543 12325 5577 12359
rect 7250 12325 7284 12359
rect 9413 12325 9447 12359
rect 10885 12325 10919 12359
rect 11437 12325 11471 12359
rect 12449 12325 12483 12359
rect 16405 12325 16439 12359
rect 16957 12325 16991 12359
rect 21097 12325 21131 12359
rect 2421 12257 2455 12291
rect 4204 12257 4238 12291
rect 8125 12257 8159 12291
rect 9756 12257 9790 12291
rect 14264 12257 14298 12291
rect 17785 12257 17819 12291
rect 20177 12257 20211 12291
rect 22512 12257 22546 12291
rect 23524 12257 23558 12291
rect 2789 12189 2823 12223
rect 3433 12189 3467 12223
rect 5181 12189 5215 12223
rect 6929 12189 6963 12223
rect 10793 12189 10827 12223
rect 12357 12189 12391 12223
rect 12633 12189 12667 12223
rect 13369 12189 13403 12223
rect 16313 12189 16347 12223
rect 18889 12189 18923 12223
rect 20729 12189 20763 12223
rect 21005 12189 21039 12223
rect 23627 12189 23661 12223
rect 2697 12121 2731 12155
rect 3801 12121 3835 12155
rect 4997 12121 5031 12155
rect 10149 12121 10183 12155
rect 18797 12121 18831 12155
rect 21557 12121 21591 12155
rect 1869 12053 1903 12087
rect 2237 12053 2271 12087
rect 2559 12053 2593 12087
rect 3065 12053 3099 12087
rect 6101 12053 6135 12087
rect 6469 12053 6503 12087
rect 6837 12053 6871 12087
rect 9827 12053 9861 12087
rect 10517 12053 10551 12087
rect 14335 12053 14369 12087
rect 16037 12053 16071 12087
rect 17923 12053 17957 12087
rect 22615 12053 22649 12087
rect 1961 11849 1995 11883
rect 2329 11849 2363 11883
rect 4629 11849 4663 11883
rect 6285 11849 6319 11883
rect 8401 11849 8435 11883
rect 9689 11849 9723 11883
rect 10701 11849 10735 11883
rect 10977 11849 11011 11883
rect 11437 11849 11471 11883
rect 12265 11849 12299 11883
rect 12817 11849 12851 11883
rect 15853 11849 15887 11883
rect 19441 11849 19475 11883
rect 20637 11849 20671 11883
rect 22477 11849 22511 11883
rect 23765 11849 23799 11883
rect 24777 11849 24811 11883
rect 2218 11781 2252 11815
rect 3065 11781 3099 11815
rect 13921 11781 13955 11815
rect 17417 11781 17451 11815
rect 17693 11781 17727 11815
rect 2421 11713 2455 11747
rect 3433 11713 3467 11747
rect 4353 11713 4387 11747
rect 11805 11713 11839 11747
rect 13001 11713 13035 11747
rect 15117 11713 15151 11747
rect 16405 11713 16439 11747
rect 16681 11713 16715 11747
rect 2053 11645 2087 11679
rect 3801 11645 3835 11679
rect 4169 11645 4203 11679
rect 5457 11645 5491 11679
rect 5733 11645 5767 11679
rect 5917 11645 5951 11679
rect 6837 11645 6871 11679
rect 8033 11645 8067 11679
rect 8836 11645 8870 11679
rect 9781 11645 9815 11679
rect 18429 11713 18463 11747
rect 19625 11645 19659 11679
rect 20085 11645 20119 11679
rect 21189 11645 21223 11679
rect 21649 11645 21683 11679
rect 2789 11577 2823 11611
rect 7158 11577 7192 11611
rect 9229 11577 9263 11611
rect 10143 11577 10177 11611
rect 13322 11577 13356 11611
rect 14289 11577 14323 11611
rect 14657 11577 14691 11611
rect 14830 11577 14864 11611
rect 14933 11577 14967 11611
rect 16221 11577 16255 11611
rect 16497 11577 16531 11611
rect 17693 11577 17727 11611
rect 18153 11577 18187 11611
rect 18245 11577 18279 11611
rect 24593 11645 24627 11679
rect 25145 11645 25179 11679
rect 5089 11509 5123 11543
rect 6653 11509 6687 11543
rect 7757 11509 7791 11543
rect 8907 11509 8941 11543
rect 17785 11509 17819 11543
rect 19165 11509 19199 11543
rect 19901 11509 19935 11543
rect 21005 11509 21039 11543
rect 21281 11509 21315 11543
rect 23765 11509 23799 11543
rect 23949 11509 23983 11543
rect 3801 11305 3835 11339
rect 5273 11305 5307 11339
rect 8861 11305 8895 11339
rect 12449 11305 12483 11339
rect 13369 11305 13403 11339
rect 13921 11305 13955 11339
rect 14841 11305 14875 11339
rect 16405 11305 16439 11339
rect 16681 11305 16715 11339
rect 18153 11305 18187 11339
rect 18521 11305 18555 11339
rect 20637 11305 20671 11339
rect 3111 11237 3145 11271
rect 6009 11237 6043 11271
rect 6110 11237 6144 11271
rect 7297 11237 7331 11271
rect 7665 11237 7699 11271
rect 9873 11237 9907 11271
rect 10149 11237 10183 11271
rect 10241 11237 10275 11271
rect 10793 11237 10827 11271
rect 15393 11237 15427 11271
rect 15485 11237 15519 11271
rect 17049 11237 17083 11271
rect 17601 11237 17635 11271
rect 21097 11237 21131 11271
rect 1501 11169 1535 11203
rect 3008 11169 3042 11203
rect 4353 11169 4387 11203
rect 4629 11169 4663 11203
rect 11989 11169 12023 11203
rect 12127 11169 12161 11203
rect 18429 11169 18463 11203
rect 18889 11169 18923 11203
rect 22512 11169 22546 11203
rect 2145 11101 2179 11135
rect 2789 11101 2823 11135
rect 4721 11101 4755 11135
rect 7573 11101 7607 11135
rect 7849 11101 7883 11135
rect 9229 11101 9263 11135
rect 13001 11101 13035 11135
rect 16957 11101 16991 11135
rect 19625 11101 19659 11135
rect 21005 11101 21039 11135
rect 21649 11101 21683 11135
rect 23489 11101 23523 11135
rect 2421 11033 2455 11067
rect 6561 11033 6595 11067
rect 15945 11033 15979 11067
rect 3433 10965 3467 10999
rect 5549 10965 5583 10999
rect 6929 10965 6963 10999
rect 8493 10965 8527 10999
rect 12909 10965 12943 10999
rect 14289 10965 14323 10999
rect 22615 10965 22649 10999
rect 1501 10761 1535 10795
rect 4261 10761 4295 10795
rect 5089 10761 5123 10795
rect 8217 10761 8251 10795
rect 11345 10761 11379 10795
rect 12679 10761 12713 10795
rect 16313 10761 16347 10795
rect 19257 10761 19291 10795
rect 20729 10761 20763 10795
rect 21097 10761 21131 10795
rect 9505 10693 9539 10727
rect 13369 10693 13403 10727
rect 14749 10693 14783 10727
rect 15945 10693 15979 10727
rect 17095 10693 17129 10727
rect 24777 10693 24811 10727
rect 4629 10625 4663 10659
rect 9137 10625 9171 10659
rect 10977 10625 11011 10659
rect 13645 10625 13679 10659
rect 14289 10625 14323 10659
rect 15209 10625 15243 10659
rect 16773 10625 16807 10659
rect 18061 10625 18095 10659
rect 19809 10625 19843 10659
rect 21649 10625 21683 10659
rect 22017 10625 22051 10659
rect 1685 10557 1719 10591
rect 1961 10557 1995 10591
rect 5181 10557 5215 10591
rect 5733 10557 5767 10591
rect 8401 10557 8435 10591
rect 8953 10557 8987 10591
rect 12608 10557 12642 10591
rect 13001 10557 13035 10591
rect 16992 10557 17026 10591
rect 17417 10557 17451 10591
rect 18981 10557 19015 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 3065 10489 3099 10523
rect 3157 10489 3191 10523
rect 3709 10489 3743 10523
rect 5917 10489 5951 10523
rect 6929 10489 6963 10523
rect 7021 10489 7055 10523
rect 7573 10489 7607 10523
rect 7941 10489 7975 10523
rect 10057 10489 10091 10523
rect 10149 10489 10183 10523
rect 10701 10489 10735 10523
rect 12081 10489 12115 10523
rect 13737 10489 13771 10523
rect 15393 10489 15427 10523
rect 15485 10489 15519 10523
rect 18382 10489 18416 10523
rect 20130 10489 20164 10523
rect 21741 10489 21775 10523
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 9873 10421 9907 10455
rect 17785 10421 17819 10455
rect 19625 10421 19659 10455
rect 21465 10421 21499 10455
rect 22569 10421 22603 10455
rect 2237 10217 2271 10251
rect 4261 10217 4295 10251
rect 5641 10217 5675 10251
rect 7481 10217 7515 10251
rect 7849 10217 7883 10251
rect 13001 10217 13035 10251
rect 13921 10217 13955 10251
rect 15393 10217 15427 10251
rect 16773 10217 16807 10251
rect 17233 10217 17267 10251
rect 19993 10217 20027 10251
rect 20637 10217 20671 10251
rect 21925 10217 21959 10251
rect 3433 10149 3467 10183
rect 3801 10149 3835 10183
rect 5083 10149 5117 10183
rect 6653 10149 6687 10183
rect 9965 10149 9999 10183
rect 11529 10149 11563 10183
rect 19073 10149 19107 10183
rect 21097 10149 21131 10183
rect 1476 10081 1510 10115
rect 2513 10081 2547 10115
rect 2973 10081 3007 10115
rect 5917 10081 5951 10115
rect 8033 10081 8067 10115
rect 8493 10081 8527 10115
rect 12909 10081 12943 10115
rect 13369 10081 13403 10115
rect 15301 10081 15335 10115
rect 15853 10081 15887 10115
rect 17325 10081 17359 10115
rect 17785 10081 17819 10115
rect 18521 10081 18555 10115
rect 22512 10081 22546 10115
rect 3157 10013 3191 10047
rect 4721 10013 4755 10047
rect 6561 10013 6595 10047
rect 8769 10013 8803 10047
rect 9873 10013 9907 10047
rect 10149 10013 10183 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 18061 10013 18095 10047
rect 18981 10013 19015 10047
rect 19625 10013 19659 10047
rect 21005 10013 21039 10047
rect 21281 10013 21315 10047
rect 1547 9945 1581 9979
rect 7113 9945 7147 9979
rect 9045 9945 9079 9979
rect 1869 9877 1903 9911
rect 6377 9877 6411 9911
rect 9505 9877 9539 9911
rect 10885 9877 10919 9911
rect 15025 9877 15059 9911
rect 16497 9877 16531 9911
rect 22615 9877 22649 9911
rect 2053 9673 2087 9707
rect 2421 9673 2455 9707
rect 5825 9673 5859 9707
rect 6469 9673 6503 9707
rect 8033 9673 8067 9707
rect 9873 9673 9907 9707
rect 10149 9673 10183 9707
rect 11713 9673 11747 9707
rect 12265 9673 12299 9707
rect 15761 9673 15795 9707
rect 16129 9673 16163 9707
rect 17417 9673 17451 9707
rect 19257 9673 19291 9707
rect 21005 9673 21039 9707
rect 22477 9673 22511 9707
rect 1639 9605 1673 9639
rect 5181 9605 5215 9639
rect 10517 9605 10551 9639
rect 11345 9605 11379 9639
rect 20453 9605 20487 9639
rect 22845 9605 22879 9639
rect 23811 9605 23845 9639
rect 4261 9537 4295 9571
rect 7021 9537 7055 9571
rect 8953 9537 8987 9571
rect 13921 9537 13955 9571
rect 18061 9537 18095 9571
rect 19901 9537 19935 9571
rect 24133 9537 24167 9571
rect 1409 9469 1443 9503
rect 2513 9469 2547 9503
rect 8861 9469 8895 9503
rect 18981 9469 19015 9503
rect 23740 9469 23774 9503
rect 2875 9401 2909 9435
rect 3801 9401 3835 9435
rect 4077 9401 4111 9435
rect 4169 9401 4203 9435
rect 4582 9401 4616 9435
rect 5457 9401 5491 9435
rect 7113 9401 7147 9435
rect 7665 9401 7699 9435
rect 9315 9401 9349 9435
rect 10793 9401 10827 9435
rect 10885 9401 10919 9435
rect 13277 9401 13311 9435
rect 13369 9401 13403 9435
rect 14841 9401 14875 9435
rect 14933 9401 14967 9435
rect 15485 9401 15519 9435
rect 16497 9401 16531 9435
rect 16589 9401 16623 9435
rect 17141 9401 17175 9435
rect 18382 9401 18416 9435
rect 19993 9401 20027 9435
rect 21465 9401 21499 9435
rect 21557 9401 21591 9435
rect 22109 9401 22143 9435
rect 3433 9333 3467 9367
rect 8493 9333 8527 9367
rect 12909 9333 12943 9367
rect 14197 9333 14231 9367
rect 14565 9333 14599 9367
rect 17785 9333 17819 9367
rect 19717 9333 19751 9367
rect 2513 9129 2547 9163
rect 5917 9129 5951 9163
rect 7021 9129 7055 9163
rect 7297 9129 7331 9163
rect 9045 9129 9079 9163
rect 10057 9129 10091 9163
rect 10609 9129 10643 9163
rect 11575 9129 11609 9163
rect 11897 9129 11931 9163
rect 13829 9129 13863 9163
rect 18245 9129 18279 9163
rect 19809 9129 19843 9163
rect 20269 9129 20303 9163
rect 20729 9129 20763 9163
rect 21925 9129 21959 9163
rect 4445 9061 4479 9095
rect 4721 9061 4755 9095
rect 6422 9061 6456 9095
rect 9413 9061 9447 9095
rect 13230 9061 13264 9095
rect 15485 9061 15519 9095
rect 17049 9061 17083 9095
rect 21097 9061 21131 9095
rect 1476 8993 1510 9027
rect 2697 8993 2731 9027
rect 2881 8993 2915 9027
rect 3433 8993 3467 9027
rect 6101 8993 6135 9027
rect 8033 8993 8067 9027
rect 8585 8993 8619 9027
rect 11437 8993 11471 9027
rect 18429 8993 18463 9027
rect 18889 8993 18923 9027
rect 22512 8993 22546 9027
rect 23524 8993 23558 9027
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 5273 8925 5307 8959
rect 8769 8925 8803 8959
rect 9689 8925 9723 8959
rect 12909 8925 12943 8959
rect 15393 8925 15427 8959
rect 16957 8925 16991 8959
rect 17233 8925 17267 8959
rect 17877 8925 17911 8959
rect 19165 8925 19199 8959
rect 19441 8925 19475 8959
rect 21005 8925 21039 8959
rect 22615 8925 22649 8959
rect 1547 8857 1581 8891
rect 15945 8857 15979 8891
rect 21557 8857 21591 8891
rect 1961 8789 1995 8823
rect 2329 8789 2363 8823
rect 5549 8789 5583 8823
rect 7757 8789 7791 8823
rect 10885 8789 10919 8823
rect 12817 8789 12851 8823
rect 14841 8789 14875 8823
rect 16497 8789 16531 8823
rect 23627 8789 23661 8823
rect 2237 8585 2271 8619
rect 2881 8585 2915 8619
rect 5825 8585 5859 8619
rect 8033 8585 8067 8619
rect 9781 8585 9815 8619
rect 11069 8585 11103 8619
rect 14289 8585 14323 8619
rect 16129 8585 16163 8619
rect 16497 8585 16531 8619
rect 17785 8585 17819 8619
rect 18429 8585 18463 8619
rect 19901 8585 19935 8619
rect 20269 8585 20303 8619
rect 21741 8585 21775 8619
rect 23121 8585 23155 8619
rect 23857 8585 23891 8619
rect 1869 8517 1903 8551
rect 2605 8517 2639 8551
rect 1961 8449 1995 8483
rect 1740 8381 1774 8415
rect 1593 8313 1627 8347
rect 7573 8517 7607 8551
rect 10701 8517 10735 8551
rect 12909 8517 12943 8551
rect 14657 8517 14691 8551
rect 16819 8517 16853 8551
rect 3249 8449 3283 8483
rect 3709 8449 3743 8483
rect 4905 8449 4939 8483
rect 7021 8449 7055 8483
rect 13369 8449 13403 8483
rect 15025 8449 15059 8483
rect 15209 8449 15243 8483
rect 18981 8449 19015 8483
rect 20821 8449 20855 8483
rect 8493 8381 8527 8415
rect 8953 8381 8987 8415
rect 16716 8381 16750 8415
rect 22328 8381 22362 8415
rect 22753 8381 22787 8415
rect 3341 8313 3375 8347
rect 5267 8313 5301 8347
rect 6653 8313 6687 8347
rect 7113 8313 7147 8347
rect 9229 8313 9263 8347
rect 10149 8313 10183 8347
rect 10241 8313 10275 8347
rect 13690 8313 13724 8347
rect 15301 8313 15335 8347
rect 15853 8313 15887 8347
rect 18797 8313 18831 8347
rect 19302 8313 19336 8347
rect 20913 8313 20947 8347
rect 21465 8313 21499 8347
rect 2881 8245 2915 8279
rect 2973 8245 3007 8279
rect 4261 8245 4295 8279
rect 4813 8245 4847 8279
rect 6101 8245 6135 8279
rect 8309 8245 8343 8279
rect 11529 8245 11563 8279
rect 17141 8245 17175 8279
rect 20637 8245 20671 8279
rect 22109 8245 22143 8279
rect 22431 8245 22465 8279
rect 1961 8041 1995 8075
rect 3801 8041 3835 8075
rect 4445 8041 4479 8075
rect 6101 8041 6135 8075
rect 8263 8041 8297 8075
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 12081 8041 12115 8075
rect 13001 8041 13035 8075
rect 13645 8041 13679 8075
rect 15117 8041 15151 8075
rect 15485 8041 15519 8075
rect 15899 8041 15933 8075
rect 16681 8041 16715 8075
rect 17693 8041 17727 8075
rect 5175 7973 5209 8007
rect 6745 7973 6779 8007
rect 17094 7973 17128 8007
rect 21097 7973 21131 8007
rect 21649 7973 21683 8007
rect 2697 7905 2731 7939
rect 2881 7905 2915 7939
rect 3433 7905 3467 7939
rect 5733 7905 5767 7939
rect 8192 7905 8226 7939
rect 10241 7905 10275 7939
rect 11989 7905 12023 7939
rect 12449 7905 12483 7939
rect 13553 7905 13587 7939
rect 14105 7905 14139 7939
rect 15828 7905 15862 7939
rect 18521 7905 18555 7939
rect 18981 7905 19015 7939
rect 3157 7837 3191 7871
rect 4813 7837 4847 7871
rect 6653 7837 6687 7871
rect 6929 7837 6963 7871
rect 13369 7837 13403 7871
rect 16773 7837 16807 7871
rect 19257 7837 19291 7871
rect 21005 7837 21039 7871
rect 1685 7701 1719 7735
rect 7941 7701 7975 7735
rect 11161 7701 11195 7735
rect 3433 7497 3467 7531
rect 3893 7497 3927 7531
rect 5733 7497 5767 7531
rect 6653 7497 6687 7531
rect 9413 7497 9447 7531
rect 9735 7497 9769 7531
rect 10057 7497 10091 7531
rect 14013 7497 14047 7531
rect 14427 7497 14461 7531
rect 15209 7497 15243 7531
rect 17003 7497 17037 7531
rect 17325 7497 17359 7531
rect 18981 7497 19015 7531
rect 19257 7497 19291 7531
rect 20361 7497 20395 7531
rect 22385 7497 22419 7531
rect 2789 7429 2823 7463
rect 6975 7429 7009 7463
rect 10425 7429 10459 7463
rect 11253 7429 11287 7463
rect 13093 7429 13127 7463
rect 13645 7429 13679 7463
rect 15945 7429 15979 7463
rect 22109 7429 22143 7463
rect 2053 7361 2087 7395
rect 2973 7361 3007 7395
rect 4905 7361 4939 7395
rect 7389 7361 7423 7395
rect 10701 7361 10735 7395
rect 11713 7361 11747 7395
rect 12541 7361 12575 7395
rect 18061 7361 18095 7395
rect 19441 7361 19475 7395
rect 21005 7361 21039 7395
rect 1501 7293 1535 7327
rect 1685 7293 1719 7327
rect 2329 7293 2363 7327
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 4813 7293 4847 7327
rect 6904 7293 6938 7327
rect 9664 7293 9698 7327
rect 14356 7293 14390 7327
rect 14749 7293 14783 7327
rect 16900 7293 16934 7327
rect 17693 7293 17727 7327
rect 21189 7293 21223 7327
rect 7941 7225 7975 7259
rect 8033 7225 8067 7259
rect 8585 7225 8619 7259
rect 10793 7225 10827 7259
rect 12633 7225 12667 7259
rect 15393 7225 15427 7259
rect 15485 7225 15519 7259
rect 19762 7225 19796 7259
rect 21510 7225 21544 7259
rect 5365 7157 5399 7191
rect 6193 7157 6227 7191
rect 7757 7157 7791 7191
rect 8953 7157 8987 7191
rect 11989 7157 12023 7191
rect 16313 7157 16347 7191
rect 16773 7157 16807 7191
rect 18521 7157 18555 7191
rect 20637 7157 20671 7191
rect 1685 6953 1719 6987
rect 2513 6953 2547 6987
rect 5871 6953 5905 6987
rect 8217 6953 8251 6987
rect 10609 6953 10643 6987
rect 10885 6953 10919 6987
rect 16957 6953 16991 6987
rect 19533 6953 19567 6987
rect 20729 6953 20763 6987
rect 1409 6885 1443 6919
rect 7659 6885 7693 6919
rect 10010 6885 10044 6919
rect 11621 6885 11655 6919
rect 12449 6885 12483 6919
rect 13553 6885 13587 6919
rect 13829 6885 13863 6919
rect 15485 6885 15519 6919
rect 16037 6885 16071 6919
rect 21097 6885 21131 6919
rect 1593 6817 1627 6851
rect 3040 6817 3074 6851
rect 4261 6817 4295 6851
rect 4629 6817 4663 6851
rect 5800 6817 5834 6851
rect 6929 6817 6963 6851
rect 9689 6817 9723 6851
rect 17141 6817 17175 6851
rect 17417 6817 17451 6851
rect 18613 6817 18647 6851
rect 18981 6817 19015 6851
rect 19257 6817 19291 6851
rect 21649 6817 21683 6851
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 7297 6749 7331 6783
rect 11529 6749 11563 6783
rect 13737 6749 13771 6783
rect 15393 6749 15427 6783
rect 21005 6749 21039 6783
rect 3111 6681 3145 6715
rect 8769 6681 8803 6715
rect 12081 6681 12115 6715
rect 14289 6681 14323 6715
rect 11253 6613 11287 6647
rect 12817 6613 12851 6647
rect 15117 6613 15151 6647
rect 19993 6613 20027 6647
rect 2697 6409 2731 6443
rect 3801 6409 3835 6443
rect 8585 6409 8619 6443
rect 9781 6409 9815 6443
rect 10425 6409 10459 6443
rect 11621 6409 11655 6443
rect 13921 6409 13955 6443
rect 14197 6409 14231 6443
rect 17417 6409 17451 6443
rect 19625 6409 19659 6443
rect 21005 6409 21039 6443
rect 21373 6409 21407 6443
rect 5733 6341 5767 6375
rect 11161 6341 11195 6375
rect 16865 6341 16899 6375
rect 17693 6341 17727 6375
rect 17785 6341 17819 6375
rect 18981 6341 19015 6375
rect 4353 6273 4387 6307
rect 7389 6273 7423 6307
rect 8861 6273 8895 6307
rect 9505 6273 9539 6307
rect 16957 6273 16991 6307
rect 2973 6205 3007 6239
rect 3249 6205 3283 6239
rect 6653 6205 6687 6239
rect 7113 6205 7147 6239
rect 7297 6205 7331 6239
rect 13001 6205 13035 6239
rect 14749 6205 14783 6239
rect 19901 6273 19935 6307
rect 20545 6273 20579 6307
rect 18061 6205 18095 6239
rect 19257 6205 19291 6239
rect 3525 6137 3559 6171
rect 4674 6137 4708 6171
rect 8953 6137 8987 6171
rect 10609 6137 10643 6171
rect 10701 6137 10735 6171
rect 12817 6137 12851 6171
rect 13322 6137 13356 6171
rect 14565 6137 14599 6171
rect 15070 6137 15104 6171
rect 17693 6137 17727 6171
rect 18382 6137 18416 6171
rect 19993 6137 20027 6171
rect 1593 6069 1627 6103
rect 1961 6069 1995 6103
rect 4169 6069 4203 6103
rect 5273 6069 5307 6103
rect 7849 6069 7883 6103
rect 11989 6069 12023 6103
rect 15669 6069 15703 6103
rect 15945 6069 15979 6103
rect 16405 6069 16439 6103
rect 2789 5865 2823 5899
rect 3801 5865 3835 5899
rect 4261 5865 4295 5899
rect 7389 5865 7423 5899
rect 9873 5865 9907 5899
rect 12219 5865 12253 5899
rect 18153 5865 18187 5899
rect 18521 5865 18555 5899
rect 19809 5865 19843 5899
rect 4858 5797 4892 5831
rect 6469 5797 6503 5831
rect 8217 5797 8251 5831
rect 10701 5797 10735 5831
rect 13782 5797 13816 5831
rect 15485 5797 15519 5831
rect 17049 5797 17083 5831
rect 12081 5729 12115 5763
rect 18429 5729 18463 5763
rect 18981 5729 19015 5763
rect 23556 5729 23590 5763
rect 4537 5661 4571 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 10609 5661 10643 5695
rect 13461 5661 13495 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 16957 5661 16991 5695
rect 17233 5661 17267 5695
rect 11161 5593 11195 5627
rect 5457 5525 5491 5559
rect 10333 5525 10367 5559
rect 12633 5525 12667 5559
rect 13001 5525 13035 5559
rect 14381 5525 14415 5559
rect 14749 5525 14783 5559
rect 23627 5525 23661 5559
rect 4261 5321 4295 5355
rect 6377 5321 6411 5355
rect 7849 5321 7883 5355
rect 9689 5321 9723 5355
rect 10701 5321 10735 5355
rect 10977 5321 11011 5355
rect 11437 5321 11471 5355
rect 12173 5321 12207 5355
rect 13461 5321 13495 5355
rect 13829 5321 13863 5355
rect 15209 5321 15243 5355
rect 16865 5321 16899 5355
rect 18429 5321 18463 5355
rect 23857 5321 23891 5355
rect 5733 5253 5767 5287
rect 4997 5185 5031 5219
rect 5181 5185 5215 5219
rect 6837 5185 6871 5219
rect 13001 5185 13035 5219
rect 15853 5185 15887 5219
rect 16129 5185 16163 5219
rect 17325 5185 17359 5219
rect 18843 5185 18877 5219
rect 7941 5117 7975 5151
rect 9321 5117 9355 5151
rect 9781 5117 9815 5151
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 14013 5117 14047 5151
rect 14933 5117 14967 5151
rect 15577 5117 15611 5151
rect 18756 5117 18790 5151
rect 24593 5117 24627 5151
rect 25145 5117 25179 5151
rect 5273 5049 5307 5083
rect 8263 5049 8297 5083
rect 10143 5049 10177 5083
rect 14334 5049 14368 5083
rect 15945 5049 15979 5083
rect 4537 4981 4571 5015
rect 7481 4981 7515 5015
rect 8861 4981 8895 5015
rect 19165 4981 19199 5015
rect 24777 4981 24811 5015
rect 5181 4777 5215 4811
rect 8125 4777 8159 4811
rect 8401 4777 8435 4811
rect 8769 4777 8803 4811
rect 12219 4777 12253 4811
rect 13001 4777 13035 4811
rect 14105 4777 14139 4811
rect 15117 4777 15151 4811
rect 16313 4777 16347 4811
rect 17003 4777 17037 4811
rect 18521 4777 18555 4811
rect 7567 4709 7601 4743
rect 9873 4709 9907 4743
rect 10425 4709 10459 4743
rect 12541 4709 12575 4743
rect 13829 4709 13863 4743
rect 15485 4709 15519 4743
rect 4696 4641 4730 4675
rect 5917 4641 5951 4675
rect 6101 4641 6135 4675
rect 12148 4641 12182 4675
rect 13369 4641 13403 4675
rect 13553 4641 13587 4675
rect 16865 4641 16899 4675
rect 6377 4573 6411 4607
rect 7205 4573 7239 4607
rect 9781 4573 9815 4607
rect 15393 4573 15427 4607
rect 15669 4573 15703 4607
rect 4767 4505 4801 4539
rect 6653 4505 6687 4539
rect 6101 4233 6135 4267
rect 9137 4233 9171 4267
rect 9321 4233 9355 4267
rect 10701 4233 10735 4267
rect 11253 4233 11287 4267
rect 12173 4233 12207 4267
rect 12265 4233 12299 4267
rect 12909 4233 12943 4267
rect 14381 4233 14415 4267
rect 14703 4233 14737 4267
rect 15715 4233 15749 4267
rect 16727 4233 16761 4267
rect 4721 4165 4755 4199
rect 5733 4165 5767 4199
rect 7757 4165 7791 4199
rect 8769 4165 8803 4199
rect 6996 4029 7030 4063
rect 7389 4029 7423 4063
rect 9597 4029 9631 4063
rect 9781 4029 9815 4063
rect 10149 4029 10183 4063
rect 11380 4029 11414 4063
rect 7205 3961 7239 3995
rect 8217 3961 8251 3995
rect 8309 3961 8343 3995
rect 9321 3961 9355 3995
rect 15393 4165 15427 4199
rect 13737 4097 13771 4131
rect 16129 4097 16163 4131
rect 13001 4029 13035 4063
rect 13461 4029 13495 4063
rect 14600 4029 14634 4063
rect 15025 4029 15059 4063
rect 15644 4029 15678 4063
rect 16656 4029 16690 4063
rect 17509 4029 17543 4063
rect 12265 3961 12299 3995
rect 14105 3961 14139 3995
rect 9965 3893 9999 3927
rect 11483 3893 11517 3927
rect 17049 3893 17083 3927
rect 7205 3689 7239 3723
rect 7481 3689 7515 3723
rect 8769 3689 8803 3723
rect 10379 3689 10413 3723
rect 13185 3689 13219 3723
rect 15485 3689 15519 3723
rect 19901 3689 19935 3723
rect 8401 3621 8435 3655
rect 9873 3621 9907 3655
rect 13001 3621 13035 3655
rect 7665 3553 7699 3587
rect 7849 3553 7883 3587
rect 11253 3553 11287 3587
rect 13369 3553 13403 3587
rect 13553 3553 13587 3587
rect 19717 3553 19751 3587
rect 10149 3349 10183 3383
rect 11437 3349 11471 3383
rect 6561 3145 6595 3179
rect 7251 3145 7285 3179
rect 10563 3145 10597 3179
rect 12587 3145 12621 3179
rect 13369 3145 13403 3179
rect 13921 3145 13955 3179
rect 14289 3145 14323 3179
rect 19349 3145 19383 3179
rect 19717 3145 19751 3179
rect 11345 3077 11379 3111
rect 13599 3077 13633 3111
rect 20085 3077 20119 3111
rect 24777 3077 24811 3111
rect 7941 3009 7975 3043
rect 10333 3009 10367 3043
rect 13093 3009 13127 3043
rect 7148 2941 7182 2975
rect 7573 2941 7607 2975
rect 8217 2941 8251 2975
rect 8861 2941 8895 2975
rect 10492 2941 10526 2975
rect 10977 2941 11011 2975
rect 12357 2941 12391 2975
rect 12909 2941 12943 2975
rect 13528 2941 13562 2975
rect 18956 2941 18990 2975
rect 19901 2941 19935 2975
rect 24593 2941 24627 2975
rect 25145 2941 25179 2975
rect 20453 2873 20487 2907
rect 8401 2805 8435 2839
rect 13093 2805 13127 2839
rect 19027 2805 19061 2839
rect 4399 2601 4433 2635
rect 7573 2601 7607 2635
rect 10379 2601 10413 2635
rect 12771 2601 12805 2635
rect 25237 2601 25271 2635
rect 4328 2465 4362 2499
rect 6929 2465 6963 2499
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 10276 2465 10310 2499
rect 10701 2465 10735 2499
rect 12700 2465 12734 2499
rect 13093 2465 13127 2499
rect 15945 2465 15979 2499
rect 16497 2465 16531 2499
rect 19165 2465 19199 2499
rect 19717 2465 19751 2499
rect 21373 2465 21407 2499
rect 21925 2465 21959 2499
rect 24593 2465 24627 2499
rect 8769 2329 8803 2363
rect 19349 2329 19383 2363
rect 24777 2329 24811 2363
rect 4721 2261 4755 2295
rect 7113 2261 7147 2295
rect 16129 2261 16163 2295
rect 21557 2261 21591 2295
<< metal1 >>
rect 4430 27072 4436 27124
rect 4488 27112 4494 27124
rect 5442 27112 5448 27124
rect 4488 27084 5448 27112
rect 4488 27072 4494 27084
rect 5442 27072 5448 27084
rect 5500 27072 5506 27124
rect 18966 26868 18972 26920
rect 19024 26908 19030 26920
rect 23382 26908 23388 26920
rect 19024 26880 23388 26908
rect 19024 26868 19030 26880
rect 23382 26868 23388 26880
rect 23440 26868 23446 26920
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 10112 25347 10170 25353
rect 10112 25313 10124 25347
rect 10158 25344 10170 25347
rect 10594 25344 10600 25356
rect 10158 25316 10600 25344
rect 10158 25313 10170 25316
rect 10112 25307 10170 25313
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 11057 25347 11115 25353
rect 11057 25313 11069 25347
rect 11103 25344 11115 25347
rect 11146 25344 11152 25356
rect 11103 25316 11152 25344
rect 11103 25313 11115 25316
rect 11057 25307 11115 25313
rect 11146 25304 11152 25316
rect 11204 25304 11210 25356
rect 13424 25347 13482 25353
rect 13424 25313 13436 25347
rect 13470 25344 13482 25347
rect 13998 25344 14004 25356
rect 13470 25316 14004 25344
rect 13470 25313 13482 25316
rect 13424 25307 13482 25313
rect 13998 25304 14004 25316
rect 14056 25304 14062 25356
rect 14436 25347 14494 25353
rect 14436 25313 14448 25347
rect 14482 25344 14494 25347
rect 14734 25344 14740 25356
rect 14482 25316 14740 25344
rect 14482 25313 14494 25316
rect 14436 25307 14494 25313
rect 14734 25304 14740 25316
rect 14792 25304 14798 25356
rect 10042 25100 10048 25152
rect 10100 25140 10106 25152
rect 10183 25143 10241 25149
rect 10183 25140 10195 25143
rect 10100 25112 10195 25140
rect 10100 25100 10106 25112
rect 10183 25109 10195 25112
rect 10229 25109 10241 25143
rect 10183 25103 10241 25109
rect 10778 25100 10784 25152
rect 10836 25140 10842 25152
rect 11195 25143 11253 25149
rect 11195 25140 11207 25143
rect 10836 25112 11207 25140
rect 10836 25100 10842 25112
rect 11195 25109 11207 25112
rect 11241 25109 11253 25143
rect 12802 25140 12808 25152
rect 12763 25112 12808 25140
rect 11195 25103 11253 25109
rect 12802 25100 12808 25112
rect 12860 25100 12866 25152
rect 13495 25143 13553 25149
rect 13495 25109 13507 25143
rect 13541 25140 13553 25143
rect 14090 25140 14096 25152
rect 13541 25112 14096 25140
rect 13541 25109 13553 25112
rect 13495 25103 13553 25109
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14507 25143 14565 25149
rect 14507 25109 14519 25143
rect 14553 25140 14565 25143
rect 14826 25140 14832 25152
rect 14553 25112 14832 25140
rect 14553 25109 14565 25112
rect 14507 25103 14565 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 15381 24939 15439 24945
rect 15381 24905 15393 24939
rect 15427 24936 15439 24939
rect 16390 24936 16396 24948
rect 15427 24908 16396 24936
rect 15427 24905 15439 24908
rect 15381 24899 15439 24905
rect 16390 24896 16396 24908
rect 16448 24896 16454 24948
rect 10594 24868 10600 24880
rect 10507 24840 10600 24868
rect 10594 24828 10600 24840
rect 10652 24868 10658 24880
rect 11790 24868 11796 24880
rect 10652 24840 11796 24868
rect 10652 24828 10658 24840
rect 11790 24828 11796 24840
rect 11848 24828 11854 24880
rect 14829 24871 14887 24877
rect 14829 24868 14841 24871
rect 14200 24840 14841 24868
rect 11241 24803 11299 24809
rect 11241 24769 11253 24803
rect 11287 24800 11299 24803
rect 11330 24800 11336 24812
rect 11287 24772 11336 24800
rect 11287 24769 11299 24772
rect 11241 24763 11299 24769
rect 11330 24760 11336 24772
rect 11388 24800 11394 24812
rect 12713 24803 12771 24809
rect 11388 24772 11744 24800
rect 11388 24760 11394 24772
rect 11716 24744 11744 24772
rect 12713 24769 12725 24803
rect 12759 24800 12771 24803
rect 12802 24800 12808 24812
rect 12759 24772 12808 24800
rect 12759 24769 12771 24772
rect 12713 24763 12771 24769
rect 12802 24760 12808 24772
rect 12860 24760 12866 24812
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8700 24735 8758 24741
rect 8700 24732 8712 24735
rect 8352 24704 8712 24732
rect 8352 24692 8358 24704
rect 8700 24701 8712 24704
rect 8746 24732 8758 24735
rect 9125 24735 9183 24741
rect 9125 24732 9137 24735
rect 8746 24704 9137 24732
rect 8746 24701 8758 24704
rect 8700 24695 8758 24701
rect 9125 24701 9137 24704
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 9744 24735 9802 24741
rect 9744 24701 9756 24735
rect 9790 24732 9802 24735
rect 10226 24732 10232 24744
rect 9790 24704 10232 24732
rect 9790 24701 9802 24704
rect 9744 24695 9802 24701
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 11698 24692 11704 24744
rect 11756 24732 11762 24744
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 11756 24704 11805 24732
rect 11756 24692 11762 24704
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 13725 24735 13783 24741
rect 13725 24701 13737 24735
rect 13771 24732 13783 24735
rect 13998 24732 14004 24744
rect 13771 24704 14004 24732
rect 13771 24701 13783 24704
rect 13725 24695 13783 24701
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 14200 24741 14228 24840
rect 14829 24837 14841 24840
rect 14875 24837 14887 24871
rect 14829 24831 14887 24837
rect 14200 24735 14278 24741
rect 14200 24704 14232 24735
rect 14220 24701 14232 24704
rect 14266 24701 14278 24735
rect 14220 24695 14278 24701
rect 14550 24692 14556 24744
rect 14608 24732 14614 24744
rect 15197 24735 15255 24741
rect 15197 24732 15209 24735
rect 14608 24704 15209 24732
rect 14608 24692 14614 24704
rect 15197 24701 15209 24704
rect 15243 24732 15255 24735
rect 15749 24735 15807 24741
rect 15749 24732 15761 24735
rect 15243 24704 15761 24732
rect 15243 24701 15255 24704
rect 15197 24695 15255 24701
rect 15749 24701 15761 24704
rect 15795 24701 15807 24735
rect 15749 24695 15807 24701
rect 11146 24664 11152 24676
rect 11059 24636 11152 24664
rect 11146 24624 11152 24636
rect 11204 24664 11210 24676
rect 12158 24664 12164 24676
rect 11204 24636 12164 24664
rect 11204 24624 11210 24636
rect 12158 24624 12164 24636
rect 12216 24624 12222 24676
rect 12805 24667 12863 24673
rect 12805 24633 12817 24667
rect 12851 24633 12863 24667
rect 12805 24627 12863 24633
rect 13357 24667 13415 24673
rect 13357 24633 13369 24667
rect 13403 24664 13415 24667
rect 14458 24664 14464 24676
rect 13403 24636 14464 24664
rect 13403 24633 13415 24636
rect 13357 24627 13415 24633
rect 8803 24599 8861 24605
rect 8803 24565 8815 24599
rect 8849 24596 8861 24599
rect 9030 24596 9036 24608
rect 8849 24568 9036 24596
rect 8849 24565 8861 24568
rect 8803 24559 8861 24565
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9815 24599 9873 24605
rect 9815 24596 9827 24599
rect 9364 24568 9827 24596
rect 9364 24556 9370 24568
rect 9815 24565 9827 24568
rect 9861 24565 9873 24599
rect 9815 24559 9873 24565
rect 11471 24599 11529 24605
rect 11471 24565 11483 24599
rect 11517 24596 11529 24599
rect 11698 24596 11704 24608
rect 11517 24568 11704 24596
rect 11517 24565 11529 24568
rect 11471 24559 11529 24565
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 12253 24599 12311 24605
rect 12253 24565 12265 24599
rect 12299 24596 12311 24599
rect 12618 24596 12624 24608
rect 12299 24568 12624 24596
rect 12299 24565 12311 24568
rect 12253 24559 12311 24565
rect 12618 24556 12624 24568
rect 12676 24596 12682 24608
rect 12820 24596 12848 24627
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 14645 24667 14703 24673
rect 14645 24633 14657 24667
rect 14691 24664 14703 24667
rect 14829 24667 14887 24673
rect 14829 24664 14841 24667
rect 14691 24636 14841 24664
rect 14691 24633 14703 24636
rect 14645 24627 14703 24633
rect 14829 24633 14841 24636
rect 14875 24664 14887 24667
rect 15838 24664 15844 24676
rect 14875 24636 15844 24664
rect 14875 24633 14887 24636
rect 14829 24627 14887 24633
rect 15838 24624 15844 24636
rect 15896 24624 15902 24676
rect 12676 24568 12848 24596
rect 12676 24556 12682 24568
rect 13722 24556 13728 24608
rect 13780 24596 13786 24608
rect 14323 24599 14381 24605
rect 14323 24596 14335 24599
rect 13780 24568 14335 24596
rect 13780 24556 13786 24568
rect 14323 24565 14335 24568
rect 14369 24565 14381 24599
rect 14323 24559 14381 24565
rect 14734 24556 14740 24608
rect 14792 24596 14798 24608
rect 15105 24599 15163 24605
rect 15105 24596 15117 24599
rect 14792 24568 15117 24596
rect 14792 24556 14798 24568
rect 15105 24565 15117 24568
rect 15151 24596 15163 24599
rect 15930 24596 15936 24608
rect 15151 24568 15936 24596
rect 15151 24565 15163 24568
rect 15105 24559 15163 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 11698 24352 11704 24404
rect 11756 24392 11762 24404
rect 11885 24395 11943 24401
rect 11885 24392 11897 24395
rect 11756 24364 11897 24392
rect 11756 24352 11762 24364
rect 11885 24361 11897 24364
rect 11931 24361 11943 24395
rect 11885 24355 11943 24361
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 15378 24392 15384 24404
rect 14323 24364 15384 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 4706 24284 4712 24336
rect 4764 24324 4770 24336
rect 6730 24324 6736 24336
rect 4764 24296 6736 24324
rect 4764 24284 4770 24296
rect 6730 24284 6736 24296
rect 6788 24324 6794 24336
rect 11900 24324 11928 24355
rect 15378 24352 15384 24364
rect 15436 24352 15442 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 17402 24392 17408 24404
rect 15519 24364 17408 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 17773 24395 17831 24401
rect 17773 24361 17785 24395
rect 17819 24392 17831 24395
rect 19426 24392 19432 24404
rect 17819 24364 19432 24392
rect 17819 24361 17831 24364
rect 17773 24355 17831 24361
rect 19426 24352 19432 24364
rect 19484 24352 19490 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 27706 24392 27712 24404
rect 24811 24364 27712 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 27706 24352 27712 24364
rect 27764 24352 27770 24404
rect 12529 24327 12587 24333
rect 12529 24324 12541 24327
rect 6788 24296 7639 24324
rect 11900 24296 12541 24324
rect 6788 24284 6794 24296
rect 7611 24268 7639 24296
rect 12529 24293 12541 24296
rect 12575 24293 12587 24327
rect 12529 24287 12587 24293
rect 12618 24284 12624 24336
rect 12676 24324 12682 24336
rect 12676 24296 12721 24324
rect 12676 24284 12682 24296
rect 13446 24284 13452 24336
rect 13504 24324 13510 24336
rect 13906 24324 13912 24336
rect 13504 24296 13912 24324
rect 13504 24284 13510 24296
rect 13906 24284 13912 24296
rect 13964 24324 13970 24336
rect 13964 24296 16528 24324
rect 13964 24284 13970 24296
rect 6178 24216 6184 24268
rect 6236 24256 6242 24268
rect 6584 24259 6642 24265
rect 6584 24256 6596 24259
rect 6236 24228 6596 24256
rect 6236 24216 6242 24228
rect 6584 24225 6596 24228
rect 6630 24225 6642 24259
rect 7558 24256 7564 24268
rect 7616 24265 7639 24268
rect 7616 24259 7654 24265
rect 7506 24228 7564 24256
rect 6584 24219 6642 24225
rect 7558 24216 7564 24228
rect 7642 24225 7654 24259
rect 7616 24219 7654 24225
rect 8640 24259 8698 24265
rect 8640 24225 8652 24259
rect 8686 24256 8698 24259
rect 9398 24256 9404 24268
rect 8686 24228 9404 24256
rect 8686 24225 8698 24228
rect 8640 24219 8698 24225
rect 7616 24216 7622 24219
rect 9398 24216 9404 24228
rect 9456 24216 9462 24268
rect 10410 24256 10416 24268
rect 10371 24228 10416 24256
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 13998 24216 14004 24268
rect 14056 24256 14062 24268
rect 14093 24259 14151 24265
rect 14093 24256 14105 24259
rect 14056 24228 14105 24256
rect 14056 24216 14062 24228
rect 14093 24225 14105 24228
rect 14139 24225 14151 24259
rect 14093 24219 14151 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15562 24256 15568 24268
rect 15335 24228 15568 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15562 24216 15568 24228
rect 15620 24256 15626 24268
rect 16500 24265 16528 24296
rect 15841 24259 15899 24265
rect 15841 24256 15853 24259
rect 15620 24228 15853 24256
rect 15620 24216 15626 24228
rect 15841 24225 15853 24228
rect 15887 24225 15899 24259
rect 15841 24219 15899 24225
rect 16485 24259 16543 24265
rect 16485 24225 16497 24259
rect 16531 24256 16543 24259
rect 16574 24256 16580 24268
rect 16531 24228 16580 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16574 24216 16580 24228
rect 16632 24216 16638 24268
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 17678 24256 17684 24268
rect 17635 24228 17684 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 23017 24259 23075 24265
rect 23017 24225 23029 24259
rect 23063 24256 23075 24259
rect 23106 24256 23112 24268
rect 23063 24228 23112 24256
rect 23063 24225 23075 24228
rect 23017 24219 23075 24225
rect 23106 24216 23112 24228
rect 23164 24216 23170 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25130 24256 25136 24268
rect 24627 24228 25136 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 27614 24188 27620 24200
rect 23446 24160 27620 24188
rect 106 24080 112 24132
rect 164 24120 170 24132
rect 10597 24123 10655 24129
rect 10597 24120 10609 24123
rect 164 24092 10609 24120
rect 164 24080 170 24092
rect 10597 24089 10609 24092
rect 10643 24089 10655 24123
rect 13078 24120 13084 24132
rect 13039 24092 13084 24120
rect 10597 24083 10655 24089
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 16669 24123 16727 24129
rect 16669 24089 16681 24123
rect 16715 24120 16727 24123
rect 23446 24120 23474 24160
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 16715 24092 23474 24120
rect 16715 24089 16727 24092
rect 16669 24083 16727 24089
rect 6687 24055 6745 24061
rect 6687 24021 6699 24055
rect 6733 24052 6745 24055
rect 6914 24052 6920 24064
rect 6733 24024 6920 24052
rect 6733 24021 6745 24024
rect 6687 24015 6745 24021
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 7699 24055 7757 24061
rect 7699 24021 7711 24055
rect 7745 24052 7757 24055
rect 7834 24052 7840 24064
rect 7745 24024 7840 24052
rect 7745 24021 7757 24024
rect 7699 24015 7757 24021
rect 7834 24012 7840 24024
rect 7892 24012 7898 24064
rect 8711 24055 8769 24061
rect 8711 24021 8723 24055
rect 8757 24052 8769 24055
rect 9214 24052 9220 24064
rect 8757 24024 9220 24052
rect 8757 24021 8769 24024
rect 8711 24015 8769 24021
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 10870 24012 10876 24064
rect 10928 24052 10934 24064
rect 10965 24055 11023 24061
rect 10965 24052 10977 24055
rect 10928 24024 10977 24052
rect 10928 24012 10934 24024
rect 10965 24021 10977 24024
rect 11011 24021 11023 24055
rect 12250 24052 12256 24064
rect 12211 24024 12256 24052
rect 10965 24015 11023 24021
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 21910 24012 21916 24064
rect 21968 24052 21974 24064
rect 23155 24055 23213 24061
rect 23155 24052 23167 24055
rect 21968 24024 23167 24052
rect 21968 24012 21974 24024
rect 23155 24021 23167 24024
rect 23201 24021 23213 24055
rect 23155 24015 23213 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 5077 23851 5135 23857
rect 5077 23817 5089 23851
rect 5123 23848 5135 23851
rect 6454 23848 6460 23860
rect 5123 23820 6460 23848
rect 5123 23817 5135 23820
rect 5077 23811 5135 23817
rect 6454 23808 6460 23820
rect 6512 23808 6518 23860
rect 7193 23851 7251 23857
rect 7193 23817 7205 23851
rect 7239 23848 7251 23851
rect 8386 23848 8392 23860
rect 7239 23820 8392 23848
rect 7239 23817 7251 23820
rect 7193 23811 7251 23817
rect 8386 23808 8392 23820
rect 8444 23808 8450 23860
rect 8665 23851 8723 23857
rect 8665 23817 8677 23851
rect 8711 23848 8723 23851
rect 9398 23848 9404 23860
rect 8711 23820 9404 23848
rect 8711 23817 8723 23820
rect 8665 23811 8723 23817
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10229 23851 10287 23857
rect 10229 23848 10241 23851
rect 10192 23820 10241 23848
rect 10192 23808 10198 23820
rect 10229 23817 10241 23820
rect 10275 23817 10287 23851
rect 10229 23811 10287 23817
rect 10410 23808 10416 23860
rect 10468 23848 10474 23860
rect 10689 23851 10747 23857
rect 10689 23848 10701 23851
rect 10468 23820 10701 23848
rect 10468 23808 10474 23820
rect 10689 23817 10701 23820
rect 10735 23848 10747 23851
rect 12342 23848 12348 23860
rect 10735 23820 12348 23848
rect 10735 23817 10747 23820
rect 10689 23811 10747 23817
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 16574 23848 16580 23860
rect 16535 23820 16580 23848
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 18230 23848 18236 23860
rect 18191 23820 18236 23848
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 20993 23851 21051 23857
rect 20993 23817 21005 23851
rect 21039 23848 21051 23851
rect 22370 23848 22376 23860
rect 21039 23820 22376 23848
rect 21039 23817 21051 23820
rect 20993 23811 21051 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 24946 23848 24952 23860
rect 24811 23820 24952 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 7558 23780 7564 23792
rect 7519 23752 7564 23780
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 13078 23780 13084 23792
rect 13039 23752 13084 23780
rect 13078 23740 13084 23752
rect 13136 23740 13142 23792
rect 13909 23783 13967 23789
rect 13909 23749 13921 23783
rect 13955 23780 13967 23783
rect 13998 23780 14004 23792
rect 13955 23752 14004 23780
rect 13955 23749 13967 23752
rect 13909 23743 13967 23749
rect 13998 23740 14004 23752
rect 14056 23780 14062 23792
rect 14642 23780 14648 23792
rect 14056 23752 14648 23780
rect 14056 23740 14062 23752
rect 14642 23740 14648 23752
rect 14700 23740 14706 23792
rect 15105 23783 15163 23789
rect 15105 23749 15117 23783
rect 15151 23780 15163 23783
rect 15378 23780 15384 23792
rect 15151 23752 15384 23780
rect 15151 23749 15163 23752
rect 15105 23743 15163 23749
rect 15378 23740 15384 23752
rect 15436 23780 15442 23792
rect 15436 23752 16068 23780
rect 15436 23740 15442 23752
rect 9907 23715 9965 23721
rect 9907 23681 9919 23715
rect 9953 23712 9965 23715
rect 12250 23712 12256 23724
rect 9953 23684 12256 23712
rect 9953 23681 9965 23684
rect 9907 23675 9965 23681
rect 12250 23672 12256 23684
rect 12308 23712 12314 23724
rect 12529 23715 12587 23721
rect 12529 23712 12541 23715
rect 12308 23684 12541 23712
rect 12308 23672 12314 23684
rect 12529 23681 12541 23684
rect 12575 23681 12587 23715
rect 14090 23712 14096 23724
rect 14051 23684 14096 23712
rect 12529 23675 12587 23681
rect 14090 23672 14096 23684
rect 14148 23672 14154 23724
rect 14458 23712 14464 23724
rect 14419 23684 14464 23712
rect 14458 23672 14464 23684
rect 14516 23672 14522 23724
rect 1118 23604 1124 23656
rect 1176 23644 1182 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 1176 23616 1444 23644
rect 1176 23604 1182 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 1857 23647 1915 23653
rect 1857 23644 1869 23647
rect 1478 23616 1869 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 1857 23613 1869 23616
rect 1903 23613 1915 23647
rect 1857 23607 1915 23613
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23644 4951 23647
rect 5445 23647 5503 23653
rect 5445 23644 5457 23647
rect 4939 23616 5457 23644
rect 4939 23613 4951 23616
rect 4893 23607 4951 23613
rect 5445 23613 5457 23616
rect 5491 23644 5503 23647
rect 5534 23644 5540 23656
rect 5491 23616 5540 23644
rect 5491 23613 5503 23616
rect 5445 23607 5503 23613
rect 5534 23604 5540 23616
rect 5592 23604 5598 23656
rect 7009 23647 7067 23653
rect 7009 23613 7021 23647
rect 7055 23613 7067 23647
rect 7009 23607 7067 23613
rect 8824 23647 8882 23653
rect 8824 23613 8836 23647
rect 8870 23644 8882 23647
rect 9309 23647 9367 23653
rect 9309 23644 9321 23647
rect 8870 23616 9321 23644
rect 8870 23613 8882 23616
rect 8824 23607 8882 23613
rect 9309 23613 9321 23616
rect 9355 23644 9367 23647
rect 9820 23647 9878 23653
rect 9820 23644 9832 23647
rect 9355 23616 9832 23644
rect 9355 23613 9367 23616
rect 9309 23607 9367 23613
rect 9820 23613 9832 23616
rect 9866 23644 9878 23647
rect 10134 23644 10140 23656
rect 9866 23616 10140 23644
rect 9866 23613 9878 23616
rect 9820 23607 9878 23613
rect 1535 23579 1593 23585
rect 1535 23545 1547 23579
rect 1581 23576 1593 23579
rect 3786 23576 3792 23588
rect 1581 23548 3792 23576
rect 1581 23545 1593 23548
rect 1535 23539 1593 23545
rect 3786 23536 3792 23548
rect 3844 23536 3850 23588
rect 5350 23536 5356 23588
rect 5408 23576 5414 23588
rect 6549 23579 6607 23585
rect 6549 23576 6561 23579
rect 5408 23548 6561 23576
rect 5408 23536 5414 23548
rect 6549 23545 6561 23548
rect 6595 23576 6607 23579
rect 7024 23576 7052 23607
rect 10134 23604 10140 23616
rect 10192 23604 10198 23656
rect 10870 23644 10876 23656
rect 10831 23616 10876 23644
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 10962 23604 10968 23656
rect 11020 23644 11026 23656
rect 16040 23653 16068 23752
rect 19518 23740 19524 23792
rect 19576 23780 19582 23792
rect 22051 23783 22109 23789
rect 22051 23780 22063 23783
rect 19576 23752 22063 23780
rect 19576 23740 19582 23752
rect 22051 23749 22063 23752
rect 22097 23749 22109 23783
rect 22051 23743 22109 23749
rect 22465 23783 22523 23789
rect 22465 23749 22477 23783
rect 22511 23780 22523 23783
rect 27430 23780 27436 23792
rect 22511 23752 27436 23780
rect 22511 23749 22523 23752
rect 22465 23743 22523 23749
rect 11241 23647 11299 23653
rect 11241 23644 11253 23647
rect 11020 23616 11253 23644
rect 11020 23604 11026 23616
rect 11241 23613 11253 23616
rect 11287 23613 11299 23647
rect 11241 23607 11299 23613
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23613 15899 23647
rect 15841 23607 15899 23613
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23613 16083 23647
rect 16025 23607 16083 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 20809 23647 20867 23653
rect 18095 23616 18736 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 6595 23548 7052 23576
rect 10888 23576 10916 23604
rect 11146 23576 11152 23588
rect 10888 23548 11152 23576
rect 6595 23545 6607 23548
rect 6549 23539 6607 23545
rect 11146 23536 11152 23548
rect 11204 23536 11210 23588
rect 11514 23576 11520 23588
rect 11475 23548 11520 23576
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 12621 23579 12679 23585
rect 12621 23545 12633 23579
rect 12667 23545 12679 23579
rect 13538 23576 13544 23588
rect 13451 23548 13544 23576
rect 12621 23539 12679 23545
rect 3881 23511 3939 23517
rect 3881 23477 3893 23511
rect 3927 23508 3939 23511
rect 4338 23508 4344 23520
rect 3927 23480 4344 23508
rect 3927 23477 3939 23480
rect 3881 23471 3939 23477
rect 4338 23468 4344 23480
rect 4396 23468 4402 23520
rect 4890 23468 4896 23520
rect 4948 23508 4954 23520
rect 6178 23508 6184 23520
rect 4948 23480 6184 23508
rect 4948 23468 4954 23480
rect 6178 23468 6184 23480
rect 6236 23468 6242 23520
rect 8895 23511 8953 23517
rect 8895 23477 8907 23511
rect 8941 23508 8953 23511
rect 9122 23508 9128 23520
rect 8941 23480 9128 23508
rect 8941 23477 8953 23480
rect 8895 23471 8953 23477
rect 9122 23468 9128 23480
rect 9180 23468 9186 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12066 23508 12072 23520
rect 11931 23480 12072 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 12250 23508 12256 23520
rect 12163 23480 12256 23508
rect 12250 23468 12256 23480
rect 12308 23508 12314 23520
rect 12636 23508 12664 23539
rect 13538 23536 13544 23548
rect 13596 23576 13602 23588
rect 14185 23579 14243 23585
rect 13596 23548 14044 23576
rect 13596 23536 13602 23548
rect 13170 23508 13176 23520
rect 12308 23480 13176 23508
rect 12308 23468 12314 23480
rect 13170 23468 13176 23480
rect 13228 23468 13234 23520
rect 14016 23508 14044 23548
rect 14185 23545 14197 23579
rect 14231 23545 14243 23579
rect 14185 23539 14243 23545
rect 14200 23508 14228 23539
rect 14274 23536 14280 23588
rect 14332 23576 14338 23588
rect 15473 23579 15531 23585
rect 15473 23576 15485 23579
rect 14332 23548 15485 23576
rect 14332 23536 14338 23548
rect 15473 23545 15485 23548
rect 15519 23576 15531 23579
rect 15856 23576 15884 23607
rect 17494 23576 17500 23588
rect 15519 23548 17500 23576
rect 15519 23545 15531 23548
rect 15473 23539 15531 23545
rect 17494 23536 17500 23548
rect 17552 23536 17558 23588
rect 15654 23508 15660 23520
rect 14016 23480 14228 23508
rect 15615 23480 15660 23508
rect 15654 23468 15660 23480
rect 15712 23468 15718 23520
rect 17678 23508 17684 23520
rect 17639 23480 17684 23508
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18708 23517 18736 23616
rect 20809 23613 20821 23647
rect 20855 23644 20867 23647
rect 21980 23647 22038 23653
rect 20855 23616 21496 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 18693 23511 18751 23517
rect 18693 23477 18705 23511
rect 18739 23508 18751 23511
rect 19058 23508 19064 23520
rect 18739 23480 19064 23508
rect 18739 23477 18751 23480
rect 18693 23471 18751 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 21468 23517 21496 23616
rect 21980 23613 21992 23647
rect 22026 23644 22038 23647
rect 22480 23644 22508 23743
rect 27430 23740 27436 23752
rect 27488 23740 27494 23792
rect 23106 23712 23112 23724
rect 23019 23684 23112 23712
rect 23106 23672 23112 23684
rect 23164 23712 23170 23724
rect 25038 23712 25044 23724
rect 23164 23684 25044 23712
rect 23164 23672 23170 23684
rect 25038 23672 25044 23684
rect 25096 23672 25102 23724
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22026 23616 22508 23644
rect 24412 23616 24593 23644
rect 22026 23613 22038 23616
rect 21980 23607 22038 23613
rect 21453 23511 21511 23517
rect 21453 23477 21465 23511
rect 21499 23508 21511 23511
rect 22922 23508 22928 23520
rect 21499 23480 22928 23508
rect 21499 23477 21511 23480
rect 21453 23471 21511 23477
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23842 23468 23848 23520
rect 23900 23508 23906 23520
rect 24412 23517 24440 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 23900 23480 24409 23508
rect 23900 23468 23906 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 5767 23307 5825 23313
rect 5767 23304 5779 23307
rect 5592 23276 5779 23304
rect 5592 23264 5598 23276
rect 5767 23273 5779 23276
rect 5813 23273 5825 23307
rect 5767 23267 5825 23273
rect 9122 23264 9128 23316
rect 9180 23304 9186 23316
rect 9861 23307 9919 23313
rect 9861 23304 9873 23307
rect 9180 23276 9873 23304
rect 9180 23264 9186 23276
rect 9861 23273 9873 23276
rect 9907 23304 9919 23307
rect 10134 23304 10140 23316
rect 9907 23276 10140 23304
rect 9907 23273 9919 23276
rect 9861 23267 9919 23273
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 12066 23264 12072 23316
rect 12124 23304 12130 23316
rect 12529 23307 12587 23313
rect 12529 23304 12541 23307
rect 12124 23276 12541 23304
rect 12124 23264 12130 23276
rect 12529 23273 12541 23276
rect 12575 23304 12587 23307
rect 12618 23304 12624 23316
rect 12575 23276 12624 23304
rect 12575 23273 12587 23276
rect 12529 23267 12587 23273
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13228 23276 14044 23304
rect 13228 23264 13234 23276
rect 4246 23236 4252 23248
rect 4207 23208 4252 23236
rect 4246 23196 4252 23208
rect 4304 23196 4310 23248
rect 11698 23196 11704 23248
rect 11756 23236 11762 23248
rect 11930 23239 11988 23245
rect 11930 23236 11942 23239
rect 11756 23208 11942 23236
rect 11756 23196 11762 23208
rect 11930 23205 11942 23208
rect 11976 23205 11988 23239
rect 11930 23199 11988 23205
rect 13538 23196 13544 23248
rect 13596 23236 13602 23248
rect 13817 23239 13875 23245
rect 13817 23236 13829 23239
rect 13596 23208 13829 23236
rect 13596 23196 13602 23208
rect 13817 23205 13829 23208
rect 13863 23205 13875 23239
rect 14016 23236 14044 23276
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14148 23276 14657 23304
rect 14148 23264 14154 23276
rect 14645 23273 14657 23276
rect 14691 23273 14703 23307
rect 14645 23267 14703 23273
rect 14752 23276 15516 23304
rect 14752 23236 14780 23276
rect 14016 23208 14780 23236
rect 13817 23199 13875 23205
rect 14826 23196 14832 23248
rect 14884 23236 14890 23248
rect 15488 23245 15516 23276
rect 15930 23264 15936 23316
rect 15988 23304 15994 23316
rect 17218 23304 17224 23316
rect 15988 23276 17224 23304
rect 15988 23264 15994 23276
rect 17218 23264 17224 23276
rect 17276 23304 17282 23316
rect 21450 23304 21456 23316
rect 17276 23276 21456 23304
rect 17276 23264 17282 23276
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 15381 23239 15439 23245
rect 15381 23236 15393 23239
rect 14884 23208 15393 23236
rect 14884 23196 14890 23208
rect 15381 23205 15393 23208
rect 15427 23205 15439 23239
rect 15381 23199 15439 23205
rect 15473 23239 15531 23245
rect 15473 23205 15485 23239
rect 15519 23236 15531 23239
rect 15746 23236 15752 23248
rect 15519 23208 15752 23236
rect 15519 23205 15531 23208
rect 15473 23199 15531 23205
rect 15746 23196 15752 23208
rect 15804 23196 15810 23248
rect 4801 23171 4859 23177
rect 4801 23137 4813 23171
rect 4847 23168 4859 23171
rect 5166 23168 5172 23180
rect 4847 23140 5172 23168
rect 4847 23137 4859 23140
rect 4801 23131 4859 23137
rect 5166 23128 5172 23140
rect 5224 23168 5230 23180
rect 5664 23171 5722 23177
rect 5664 23168 5676 23171
rect 5224 23140 5676 23168
rect 5224 23128 5230 23140
rect 5664 23137 5676 23140
rect 5710 23137 5722 23171
rect 5664 23131 5722 23137
rect 6638 23128 6644 23180
rect 6696 23168 6702 23180
rect 6768 23171 6826 23177
rect 6768 23168 6780 23171
rect 6696 23140 6780 23168
rect 6696 23128 6702 23140
rect 6768 23137 6780 23140
rect 6814 23137 6826 23171
rect 8018 23168 8024 23180
rect 7979 23140 8024 23168
rect 6768 23131 6826 23137
rect 8018 23128 8024 23140
rect 8076 23128 8082 23180
rect 8202 23168 8208 23180
rect 8163 23140 8208 23168
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 10226 23168 10232 23180
rect 10187 23140 10232 23168
rect 10226 23128 10232 23140
rect 10284 23128 10290 23180
rect 10597 23171 10655 23177
rect 10597 23137 10609 23171
rect 10643 23168 10655 23171
rect 11054 23168 11060 23180
rect 10643 23140 11060 23168
rect 10643 23137 10655 23140
rect 10597 23131 10655 23137
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 11514 23128 11520 23180
rect 11572 23168 11578 23180
rect 12986 23168 12992 23180
rect 11572 23140 12992 23168
rect 11572 23128 11578 23140
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 17402 23168 17408 23180
rect 17363 23140 17408 23168
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 17494 23128 17500 23180
rect 17552 23168 17558 23180
rect 17589 23171 17647 23177
rect 17589 23168 17601 23171
rect 17552 23140 17601 23168
rect 17552 23128 17558 23140
rect 17589 23137 17601 23140
rect 17635 23137 17647 23171
rect 17589 23131 17647 23137
rect 18760 23171 18818 23177
rect 18760 23137 18772 23171
rect 18806 23168 18818 23171
rect 18966 23168 18972 23180
rect 18806 23140 18972 23168
rect 18806 23137 18818 23140
rect 18760 23131 18818 23137
rect 18966 23128 18972 23140
rect 19024 23128 19030 23180
rect 3786 23060 3792 23112
rect 3844 23100 3850 23112
rect 4157 23103 4215 23109
rect 4157 23100 4169 23103
rect 3844 23072 4169 23100
rect 3844 23060 3850 23072
rect 4157 23069 4169 23072
rect 4203 23100 4215 23103
rect 4522 23100 4528 23112
rect 4203 23072 4528 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4522 23060 4528 23072
rect 4580 23060 4586 23112
rect 8481 23103 8539 23109
rect 8481 23069 8493 23103
rect 8527 23100 8539 23103
rect 8570 23100 8576 23112
rect 8527 23072 8576 23100
rect 8527 23069 8539 23072
rect 8481 23063 8539 23069
rect 8570 23060 8576 23072
rect 8628 23100 8634 23112
rect 8757 23103 8815 23109
rect 8757 23100 8769 23103
rect 8628 23072 8769 23100
rect 8628 23060 8634 23072
rect 8757 23069 8769 23072
rect 8803 23069 8815 23103
rect 8757 23063 8815 23069
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23100 10839 23103
rect 11609 23103 11667 23109
rect 11609 23100 11621 23103
rect 10827 23072 11621 23100
rect 10827 23069 10839 23072
rect 10781 23063 10839 23069
rect 11609 23069 11621 23072
rect 11655 23100 11667 23103
rect 11974 23100 11980 23112
rect 11655 23072 11980 23100
rect 11655 23069 11667 23072
rect 11609 23063 11667 23069
rect 11974 23060 11980 23072
rect 12032 23060 12038 23112
rect 13722 23100 13728 23112
rect 13683 23072 13728 23100
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 14458 23060 14464 23112
rect 14516 23100 14522 23112
rect 15470 23100 15476 23112
rect 14516 23072 15476 23100
rect 14516 23060 14522 23072
rect 15470 23060 15476 23072
rect 15528 23100 15534 23112
rect 15657 23103 15715 23109
rect 15657 23100 15669 23103
rect 15528 23072 15669 23100
rect 15528 23060 15534 23072
rect 15657 23069 15669 23072
rect 15703 23069 15715 23103
rect 17770 23100 17776 23112
rect 17731 23072 17776 23100
rect 15657 23063 15715 23069
rect 17770 23060 17776 23072
rect 17828 23060 17834 23112
rect 6871 23035 6929 23041
rect 6871 23001 6883 23035
rect 6917 23032 6929 23035
rect 9950 23032 9956 23044
rect 6917 23004 9956 23032
rect 6917 23001 6929 23004
rect 6871 22995 6929 23001
rect 9950 22992 9956 23004
rect 10008 22992 10014 23044
rect 14277 23035 14335 23041
rect 14277 23001 14289 23035
rect 14323 23001 14335 23035
rect 14277 22995 14335 23001
rect 2682 22964 2688 22976
rect 2643 22936 2688 22964
rect 2682 22924 2688 22936
rect 2740 22924 2746 22976
rect 7285 22967 7343 22973
rect 7285 22933 7297 22967
rect 7331 22964 7343 22967
rect 7374 22964 7380 22976
rect 7331 22936 7380 22964
rect 7331 22933 7343 22936
rect 7285 22927 7343 22933
rect 7374 22924 7380 22936
rect 7432 22924 7438 22976
rect 7653 22967 7711 22973
rect 7653 22933 7665 22967
rect 7699 22964 7711 22967
rect 7742 22964 7748 22976
rect 7699 22936 7748 22964
rect 7699 22933 7711 22936
rect 7653 22927 7711 22933
rect 7742 22924 7748 22936
rect 7800 22964 7806 22976
rect 8202 22964 8208 22976
rect 7800 22936 8208 22964
rect 7800 22924 7806 22936
rect 8202 22924 8208 22936
rect 8260 22924 8266 22976
rect 11054 22964 11060 22976
rect 11015 22936 11060 22964
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 13998 22964 14004 22976
rect 13136 22936 14004 22964
rect 13136 22924 13142 22936
rect 13998 22924 14004 22936
rect 14056 22964 14062 22976
rect 14292 22964 14320 22995
rect 14550 22992 14556 23044
rect 14608 23032 14614 23044
rect 20346 23032 20352 23044
rect 14608 23004 20352 23032
rect 14608 22992 14614 23004
rect 20346 22992 20352 23004
rect 20404 22992 20410 23044
rect 14056 22936 14320 22964
rect 15105 22967 15163 22973
rect 14056 22924 14062 22936
rect 15105 22933 15117 22967
rect 15151 22964 15163 22967
rect 15286 22964 15292 22976
rect 15151 22936 15292 22964
rect 15151 22933 15163 22936
rect 15105 22927 15163 22933
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 16758 22924 16764 22976
rect 16816 22964 16822 22976
rect 18831 22967 18889 22973
rect 18831 22964 18843 22967
rect 16816 22936 18843 22964
rect 16816 22924 16822 22936
rect 18831 22933 18843 22936
rect 18877 22933 18889 22967
rect 19886 22964 19892 22976
rect 19847 22936 19892 22964
rect 18831 22927 18889 22933
rect 19886 22924 19892 22936
rect 19944 22924 19950 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 3973 22763 4031 22769
rect 3973 22760 3985 22763
rect 3651 22732 3985 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 3973 22729 3985 22732
rect 4019 22760 4031 22763
rect 4246 22760 4252 22772
rect 4019 22732 4252 22760
rect 4019 22729 4031 22732
rect 3973 22723 4031 22729
rect 4246 22720 4252 22732
rect 4304 22720 4310 22772
rect 4338 22720 4344 22772
rect 4396 22760 4402 22772
rect 4396 22732 4441 22760
rect 4396 22720 4402 22732
rect 4522 22720 4528 22772
rect 4580 22760 4586 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 4580 22732 5825 22760
rect 4580 22720 4586 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 11974 22760 11980 22772
rect 11935 22732 11980 22760
rect 5813 22723 5871 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 13538 22720 13544 22772
rect 13596 22760 13602 22772
rect 15746 22760 15752 22772
rect 13596 22732 13814 22760
rect 15707 22732 15752 22760
rect 13596 22720 13602 22732
rect 106 22652 112 22704
rect 164 22692 170 22704
rect 164 22664 3049 22692
rect 164 22652 170 22664
rect 2682 22624 2688 22636
rect 2643 22596 2688 22624
rect 2682 22584 2688 22596
rect 2740 22584 2746 22636
rect 3021 22624 3049 22664
rect 6178 22624 6184 22636
rect 3021 22596 6184 22624
rect 6178 22584 6184 22596
rect 6236 22624 6242 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 6236 22596 6561 22624
rect 6236 22584 6242 22596
rect 6549 22593 6561 22596
rect 6595 22624 6607 22627
rect 6638 22624 6644 22636
rect 6595 22596 6644 22624
rect 6595 22593 6607 22596
rect 6549 22587 6607 22593
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7374 22624 7380 22636
rect 6963 22596 7380 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 8570 22624 8576 22636
rect 8531 22596 8576 22624
rect 8570 22584 8576 22596
rect 8628 22584 8634 22636
rect 10134 22584 10140 22636
rect 10192 22624 10198 22636
rect 10413 22627 10471 22633
rect 10413 22624 10425 22627
rect 10192 22596 10425 22624
rect 10192 22584 10198 22596
rect 10413 22593 10425 22596
rect 10459 22593 10471 22627
rect 10686 22624 10692 22636
rect 10647 22596 10692 22624
rect 10413 22587 10471 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 12986 22624 12992 22636
rect 12947 22596 12992 22624
rect 12986 22584 12992 22596
rect 13044 22584 13050 22636
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 10045 22559 10103 22565
rect 10045 22556 10057 22559
rect 1443 22528 1532 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 1504 22432 1532 22528
rect 8036 22528 10057 22556
rect 2593 22491 2651 22497
rect 2593 22457 2605 22491
rect 2639 22488 2651 22491
rect 3047 22491 3105 22497
rect 3047 22488 3059 22491
rect 2639 22460 3059 22488
rect 2639 22457 2651 22460
rect 2593 22451 2651 22457
rect 3047 22457 3059 22460
rect 3093 22488 3105 22491
rect 4154 22488 4160 22500
rect 3093 22460 4160 22488
rect 3093 22457 3105 22460
rect 3047 22451 3105 22457
rect 4154 22448 4160 22460
rect 4212 22448 4218 22500
rect 4338 22448 4344 22500
rect 4396 22488 4402 22500
rect 4525 22491 4583 22497
rect 4525 22488 4537 22491
rect 4396 22460 4537 22488
rect 4396 22448 4402 22460
rect 4525 22457 4537 22460
rect 4571 22457 4583 22491
rect 4525 22451 4583 22457
rect 4617 22491 4675 22497
rect 4617 22457 4629 22491
rect 4663 22457 4675 22491
rect 5166 22488 5172 22500
rect 5127 22460 5172 22488
rect 4617 22451 4675 22457
rect 1486 22380 1492 22432
rect 1544 22420 1550 22432
rect 1949 22423 2007 22429
rect 1949 22420 1961 22423
rect 1544 22392 1961 22420
rect 1544 22380 1550 22392
rect 1949 22389 1961 22392
rect 1995 22389 2007 22423
rect 4632 22420 4660 22451
rect 5166 22448 5172 22460
rect 5224 22448 5230 22500
rect 6273 22491 6331 22497
rect 6273 22457 6285 22491
rect 6319 22488 6331 22491
rect 7009 22491 7067 22497
rect 6319 22460 6729 22488
rect 6319 22457 6331 22460
rect 6273 22451 6331 22457
rect 4982 22420 4988 22432
rect 4632 22392 4988 22420
rect 1949 22383 2007 22389
rect 4982 22380 4988 22392
rect 5040 22420 5046 22432
rect 5445 22423 5503 22429
rect 5445 22420 5457 22423
rect 5040 22392 5457 22420
rect 5040 22380 5046 22392
rect 5445 22389 5457 22392
rect 5491 22389 5503 22423
rect 6701 22420 6729 22460
rect 7009 22457 7021 22491
rect 7055 22457 7067 22491
rect 7558 22488 7564 22500
rect 7519 22460 7564 22488
rect 7009 22451 7067 22457
rect 6822 22420 6828 22432
rect 6701 22392 6828 22420
rect 5445 22383 5503 22389
rect 6822 22380 6828 22392
rect 6880 22420 6886 22432
rect 7024 22420 7052 22451
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8036 22432 8064 22528
rect 10045 22525 10057 22528
rect 10091 22556 10103 22559
rect 10226 22556 10232 22568
rect 10091 22528 10232 22556
rect 10091 22525 10103 22528
rect 10045 22519 10103 22525
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 13786 22556 13814 22732
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 17494 22720 17500 22772
rect 17552 22760 17558 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 17552 22732 17693 22760
rect 17552 22720 17558 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 18966 22760 18972 22772
rect 18927 22732 18972 22760
rect 17681 22723 17739 22729
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 21913 22763 21971 22769
rect 21913 22729 21925 22763
rect 21959 22760 21971 22763
rect 26418 22760 26424 22772
rect 21959 22732 26424 22760
rect 21959 22729 21971 22732
rect 21913 22723 21971 22729
rect 14829 22627 14887 22633
rect 14829 22593 14841 22627
rect 14875 22624 14887 22627
rect 15286 22624 15292 22636
rect 14875 22596 15292 22624
rect 14875 22593 14887 22596
rect 14829 22587 14887 22593
rect 15286 22584 15292 22596
rect 15344 22584 15350 22636
rect 19426 22624 19432 22636
rect 16316 22596 19432 22624
rect 16316 22565 16344 22596
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 19886 22624 19892 22636
rect 19847 22596 19892 22624
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 20254 22624 20260 22636
rect 20215 22596 20260 22624
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 13786 22528 13921 22556
rect 13909 22525 13921 22528
rect 13955 22556 13967 22559
rect 14185 22559 14243 22565
rect 14185 22556 14197 22559
rect 13955 22528 14197 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 14185 22525 14197 22528
rect 14231 22525 14243 22559
rect 14185 22519 14243 22525
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 16301 22559 16359 22565
rect 16301 22556 16313 22559
rect 16255 22528 16313 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 16301 22525 16313 22528
rect 16347 22525 16359 22559
rect 16301 22519 16359 22525
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16724 22528 16773 22556
rect 16724 22516 16730 22528
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 18100 22559 18158 22565
rect 18100 22525 18112 22559
rect 18146 22556 18158 22559
rect 21428 22559 21486 22565
rect 18146 22528 18368 22556
rect 18146 22525 18158 22528
rect 18100 22519 18158 22525
rect 8481 22491 8539 22497
rect 8481 22457 8493 22491
rect 8527 22488 8539 22491
rect 8754 22488 8760 22500
rect 8527 22460 8760 22488
rect 8527 22457 8539 22460
rect 8481 22451 8539 22457
rect 8754 22448 8760 22460
rect 8812 22488 8818 22500
rect 8894 22491 8952 22497
rect 8894 22488 8906 22491
rect 8812 22460 8906 22488
rect 8812 22448 8818 22460
rect 8894 22457 8906 22460
rect 8940 22457 8952 22491
rect 10505 22491 10563 22497
rect 10505 22488 10517 22491
rect 8894 22451 8952 22457
rect 9784 22460 10517 22488
rect 9784 22432 9812 22460
rect 10505 22457 10517 22460
rect 10551 22488 10563 22491
rect 10870 22488 10876 22500
rect 10551 22460 10876 22488
rect 10551 22457 10563 22460
rect 10505 22451 10563 22457
rect 10870 22448 10876 22460
rect 10928 22448 10934 22500
rect 13310 22491 13368 22497
rect 13310 22488 13322 22491
rect 12820 22460 13322 22488
rect 6880 22392 7052 22420
rect 7929 22423 7987 22429
rect 6880 22380 6886 22392
rect 7929 22389 7941 22423
rect 7975 22420 7987 22423
rect 8018 22420 8024 22432
rect 7975 22392 8024 22420
rect 7975 22389 7987 22392
rect 7929 22383 7987 22389
rect 8018 22380 8024 22392
rect 8076 22380 8082 22432
rect 9493 22423 9551 22429
rect 9493 22389 9505 22423
rect 9539 22420 9551 22423
rect 9766 22420 9772 22432
rect 9539 22392 9772 22420
rect 9539 22389 9551 22392
rect 9493 22383 9551 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 11698 22420 11704 22432
rect 11659 22392 11704 22420
rect 11698 22380 11704 22392
rect 11756 22420 11762 22432
rect 12820 22429 12848 22460
rect 13310 22457 13322 22460
rect 13356 22457 13368 22491
rect 14921 22491 14979 22497
rect 14921 22488 14933 22491
rect 13310 22451 13368 22457
rect 14568 22460 14933 22488
rect 12805 22423 12863 22429
rect 12805 22420 12817 22423
rect 11756 22392 12817 22420
rect 11756 22380 11762 22392
rect 12805 22389 12817 22392
rect 12851 22389 12863 22423
rect 12805 22383 12863 22389
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 14568 22429 14596 22460
rect 14921 22457 14933 22460
rect 14967 22457 14979 22491
rect 15470 22488 15476 22500
rect 15431 22460 15476 22488
rect 14921 22451 14979 22457
rect 15470 22448 15476 22460
rect 15528 22448 15534 22500
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 18187 22491 18245 22497
rect 18187 22488 18199 22491
rect 16908 22460 18199 22488
rect 16908 22448 16914 22460
rect 18187 22457 18199 22460
rect 18233 22457 18245 22491
rect 18187 22451 18245 22457
rect 18340 22432 18368 22528
rect 21428 22525 21440 22559
rect 21474 22556 21486 22559
rect 21928 22556 21956 22723
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 24762 22692 24768 22704
rect 24723 22664 24768 22692
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 21474 22528 21956 22556
rect 21474 22525 21486 22528
rect 21428 22519 21486 22525
rect 22002 22516 22008 22568
rect 22060 22556 22066 22568
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 22060 22528 24593 22556
rect 22060 22516 22066 22528
rect 24581 22525 24593 22528
rect 24627 22556 24639 22559
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24627 22528 25145 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 19705 22491 19763 22497
rect 19705 22457 19717 22491
rect 19751 22488 19763 22491
rect 19981 22491 20039 22497
rect 19981 22488 19993 22491
rect 19751 22460 19993 22488
rect 19751 22457 19763 22460
rect 19705 22451 19763 22457
rect 19981 22457 19993 22460
rect 20027 22488 20039 22491
rect 20070 22488 20076 22500
rect 20027 22460 20076 22488
rect 20027 22457 20039 22460
rect 19981 22451 20039 22457
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 14553 22423 14611 22429
rect 14553 22420 14565 22423
rect 13872 22392 14565 22420
rect 13872 22380 13878 22392
rect 14553 22389 14565 22392
rect 14599 22389 14611 22423
rect 14553 22383 14611 22389
rect 16206 22380 16212 22432
rect 16264 22420 16270 22432
rect 16393 22423 16451 22429
rect 16393 22420 16405 22423
rect 16264 22392 16405 22420
rect 16264 22380 16270 22392
rect 16393 22389 16405 22392
rect 16439 22389 16451 22423
rect 16393 22383 16451 22389
rect 17405 22423 17463 22429
rect 17405 22389 17417 22423
rect 17451 22420 17463 22423
rect 17494 22420 17500 22432
rect 17451 22392 17500 22420
rect 17451 22389 17463 22392
rect 17405 22383 17463 22389
rect 17494 22380 17500 22392
rect 17552 22380 17558 22432
rect 18322 22380 18328 22432
rect 18380 22420 18386 22432
rect 18509 22423 18567 22429
rect 18509 22420 18521 22423
rect 18380 22392 18521 22420
rect 18380 22380 18386 22392
rect 18509 22389 18521 22392
rect 18555 22389 18567 22423
rect 18509 22383 18567 22389
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21499 22423 21557 22429
rect 21499 22420 21511 22423
rect 21048 22392 21511 22420
rect 21048 22380 21054 22392
rect 21499 22389 21511 22392
rect 21545 22420 21557 22423
rect 22646 22420 22652 22432
rect 21545 22392 22652 22420
rect 21545 22389 21557 22392
rect 21499 22383 21557 22389
rect 22646 22380 22652 22392
rect 22704 22380 22710 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2682 22216 2688 22228
rect 2643 22188 2688 22216
rect 2682 22176 2688 22188
rect 2740 22176 2746 22228
rect 4982 22216 4988 22228
rect 4943 22188 4988 22216
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 6822 22216 6828 22228
rect 6783 22188 6828 22216
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 9030 22216 9036 22228
rect 8991 22188 9036 22216
rect 9030 22176 9036 22188
rect 9088 22176 9094 22228
rect 9140 22188 9904 22216
rect 4154 22108 4160 22160
rect 4212 22148 4218 22160
rect 4427 22151 4485 22157
rect 4427 22148 4439 22151
rect 4212 22120 4439 22148
rect 4212 22108 4218 22120
rect 4427 22117 4439 22120
rect 4473 22148 4485 22151
rect 6267 22151 6325 22157
rect 6267 22148 6279 22151
rect 4473 22120 6279 22148
rect 4473 22117 4485 22120
rect 4427 22111 4485 22117
rect 6267 22117 6279 22120
rect 6313 22148 6325 22151
rect 6454 22148 6460 22160
rect 6313 22120 6460 22148
rect 6313 22117 6325 22120
rect 6267 22111 6325 22117
rect 6454 22108 6460 22120
rect 6512 22108 6518 22160
rect 8199 22151 8257 22157
rect 8199 22117 8211 22151
rect 8245 22148 8257 22151
rect 8662 22148 8668 22160
rect 8245 22120 8668 22148
rect 8245 22117 8257 22120
rect 8199 22111 8257 22117
rect 8662 22108 8668 22120
rect 8720 22108 8726 22160
rect 2682 22080 2688 22092
rect 2643 22052 2688 22080
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 2866 22080 2872 22092
rect 2827 22052 2872 22080
rect 2866 22040 2872 22052
rect 2924 22080 2930 22092
rect 3421 22083 3479 22089
rect 3421 22080 3433 22083
rect 2924 22052 3433 22080
rect 2924 22040 2930 22052
rect 3421 22049 3433 22052
rect 3467 22049 3479 22083
rect 3421 22043 3479 22049
rect 5166 22040 5172 22092
rect 5224 22080 5230 22092
rect 5721 22083 5779 22089
rect 5721 22080 5733 22083
rect 5224 22052 5733 22080
rect 5224 22040 5230 22052
rect 5721 22049 5733 22052
rect 5767 22080 5779 22083
rect 7558 22080 7564 22092
rect 5767 22052 7564 22080
rect 5767 22049 5779 22052
rect 5721 22043 5779 22049
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22080 8815 22083
rect 8846 22080 8852 22092
rect 8803 22052 8852 22080
rect 8803 22049 8815 22052
rect 8757 22043 8815 22049
rect 8846 22040 8852 22052
rect 8904 22080 8910 22092
rect 9140 22080 9168 22188
rect 9214 22108 9220 22160
rect 9272 22148 9278 22160
rect 9876 22157 9904 22188
rect 10870 22176 10876 22228
rect 10928 22216 10934 22228
rect 11057 22219 11115 22225
rect 11057 22216 11069 22219
rect 10928 22188 11069 22216
rect 10928 22176 10934 22188
rect 11057 22185 11069 22188
rect 11103 22185 11115 22219
rect 11057 22179 11115 22185
rect 12161 22219 12219 22225
rect 12161 22185 12173 22219
rect 12207 22216 12219 22219
rect 12250 22216 12256 22228
rect 12207 22188 12256 22216
rect 12207 22185 12219 22188
rect 12161 22179 12219 22185
rect 12250 22176 12256 22188
rect 12308 22176 12314 22228
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 14001 22219 14059 22225
rect 14001 22216 14013 22219
rect 13780 22188 14013 22216
rect 13780 22176 13786 22188
rect 14001 22185 14013 22188
rect 14047 22185 14059 22219
rect 14001 22179 14059 22185
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 15013 22219 15071 22225
rect 15013 22216 15025 22219
rect 14884 22188 15025 22216
rect 14884 22176 14890 22188
rect 15013 22185 15025 22188
rect 15059 22185 15071 22219
rect 15013 22179 15071 22185
rect 15838 22176 15844 22228
rect 15896 22216 15902 22228
rect 19659 22219 19717 22225
rect 15896 22188 19517 22216
rect 15896 22176 15902 22188
rect 9769 22151 9827 22157
rect 9769 22148 9781 22151
rect 9272 22120 9781 22148
rect 9272 22108 9278 22120
rect 9769 22117 9781 22120
rect 9815 22117 9827 22151
rect 9769 22111 9827 22117
rect 9861 22151 9919 22157
rect 9861 22117 9873 22151
rect 9907 22117 9919 22151
rect 9861 22111 9919 22117
rect 11603 22151 11661 22157
rect 11603 22117 11615 22151
rect 11649 22148 11661 22151
rect 11698 22148 11704 22160
rect 11649 22120 11704 22148
rect 11649 22117 11661 22120
rect 11603 22111 11661 22117
rect 11698 22108 11704 22120
rect 11756 22108 11762 22160
rect 13078 22108 13084 22160
rect 13136 22148 13142 22160
rect 13173 22151 13231 22157
rect 13173 22148 13185 22151
rect 13136 22120 13185 22148
rect 13136 22108 13142 22120
rect 13173 22117 13185 22120
rect 13219 22117 13231 22151
rect 15930 22148 15936 22160
rect 13173 22111 13231 22117
rect 15304 22120 15936 22148
rect 15304 22089 15332 22120
rect 15930 22108 15936 22120
rect 15988 22108 15994 22160
rect 17954 22148 17960 22160
rect 17915 22120 17960 22148
rect 17954 22108 17960 22120
rect 18012 22108 18018 22160
rect 8904 22052 9168 22080
rect 15289 22083 15347 22089
rect 8904 22040 8910 22052
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 15436 22052 15761 22080
rect 15436 22040 15442 22052
rect 15749 22049 15761 22052
rect 15795 22080 15807 22083
rect 16301 22083 16359 22089
rect 16301 22080 16313 22083
rect 15795 22052 16313 22080
rect 15795 22049 15807 22052
rect 15749 22043 15807 22049
rect 16301 22049 16313 22052
rect 16347 22080 16359 22083
rect 16666 22080 16672 22092
rect 16347 22052 16672 22080
rect 16347 22049 16359 22052
rect 16301 22043 16359 22049
rect 16666 22040 16672 22052
rect 16724 22040 16730 22092
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22080 17739 22083
rect 17770 22080 17776 22092
rect 17727 22052 17776 22080
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 17770 22040 17776 22052
rect 17828 22040 17834 22092
rect 19489 22080 19517 22188
rect 19659 22185 19671 22219
rect 19705 22216 19717 22219
rect 19978 22216 19984 22228
rect 19705 22188 19984 22216
rect 19705 22185 19717 22188
rect 19659 22179 19717 22185
rect 19978 22176 19984 22188
rect 20036 22176 20042 22228
rect 22002 22216 22008 22228
rect 20364 22188 22008 22216
rect 20364 22092 20392 22188
rect 22002 22176 22008 22188
rect 22060 22176 22066 22228
rect 20990 22148 20996 22160
rect 20951 22120 20996 22148
rect 20990 22108 20996 22120
rect 21048 22108 21054 22160
rect 21085 22151 21143 22157
rect 21085 22117 21097 22151
rect 21131 22148 21143 22151
rect 22278 22148 22284 22160
rect 21131 22120 22284 22148
rect 21131 22117 21143 22120
rect 21085 22111 21143 22117
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 19556 22083 19614 22089
rect 19556 22080 19568 22083
rect 19489 22052 19568 22080
rect 19556 22049 19568 22052
rect 19602 22080 19614 22083
rect 20346 22080 20352 22092
rect 19602 22052 20352 22080
rect 19602 22049 19614 22052
rect 19556 22043 19614 22049
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 3804 21984 4077 22012
rect 2317 21879 2375 21885
rect 2317 21845 2329 21879
rect 2363 21876 2375 21879
rect 2498 21876 2504 21888
rect 2363 21848 2504 21876
rect 2363 21845 2375 21848
rect 2317 21839 2375 21845
rect 2498 21836 2504 21848
rect 2556 21836 2562 21888
rect 3602 21836 3608 21888
rect 3660 21876 3666 21888
rect 3804 21885 3832 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 5905 22015 5963 22021
rect 5905 21981 5917 22015
rect 5951 22012 5963 22015
rect 5994 22012 6000 22024
rect 5951 21984 6000 22012
rect 5951 21981 5963 21984
rect 5905 21975 5963 21981
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 7926 22012 7932 22024
rect 7883 21984 7932 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 7926 21972 7932 21984
rect 7984 21972 7990 22024
rect 10134 22012 10140 22024
rect 10095 21984 10140 22012
rect 10134 21972 10140 21984
rect 10192 22012 10198 22024
rect 10686 22012 10692 22024
rect 10192 21984 10692 22012
rect 10192 21972 10198 21984
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 11238 22012 11244 22024
rect 11199 21984 11244 22012
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 13081 22015 13139 22021
rect 13081 22012 13093 22015
rect 12575 21984 13093 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 13081 21981 13093 21984
rect 13127 22012 13139 22015
rect 15470 22012 15476 22024
rect 13127 21984 15476 22012
rect 13127 21981 13139 21984
rect 13081 21975 13139 21981
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 15838 22012 15844 22024
rect 15799 21984 15844 22012
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 21269 22015 21327 22021
rect 21269 22012 21281 22015
rect 21232 21984 21281 22012
rect 21232 21972 21238 21984
rect 21269 21981 21281 21984
rect 21315 21981 21327 22015
rect 21269 21975 21327 21981
rect 10870 21904 10876 21956
rect 10928 21944 10934 21956
rect 11974 21944 11980 21956
rect 10928 21916 11980 21944
rect 10928 21904 10934 21916
rect 11974 21904 11980 21916
rect 12032 21944 12038 21956
rect 13633 21947 13691 21953
rect 12032 21916 13308 21944
rect 12032 21904 12038 21916
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 3660 21848 3801 21876
rect 3660 21836 3666 21848
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 5534 21836 5540 21888
rect 5592 21876 5598 21888
rect 7377 21879 7435 21885
rect 7377 21876 7389 21879
rect 5592 21848 7389 21876
rect 5592 21836 5598 21848
rect 7377 21845 7389 21848
rect 7423 21876 7435 21879
rect 7742 21876 7748 21888
rect 7423 21848 7748 21876
rect 7423 21845 7435 21848
rect 7377 21839 7435 21845
rect 7742 21836 7748 21848
rect 7800 21836 7806 21888
rect 10686 21876 10692 21888
rect 10647 21848 10692 21876
rect 10686 21836 10692 21848
rect 10744 21876 10750 21888
rect 11054 21876 11060 21888
rect 10744 21848 11060 21876
rect 10744 21836 10750 21848
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 12897 21879 12955 21885
rect 12897 21845 12909 21879
rect 12943 21876 12955 21879
rect 13078 21876 13084 21888
rect 12943 21848 13084 21876
rect 12943 21845 12955 21848
rect 12897 21839 12955 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13280 21876 13308 21916
rect 13633 21913 13645 21947
rect 13679 21944 13691 21947
rect 14458 21944 14464 21956
rect 13679 21916 14464 21944
rect 13679 21913 13691 21916
rect 13633 21907 13691 21913
rect 14458 21904 14464 21916
rect 14516 21904 14522 21956
rect 14274 21876 14280 21888
rect 13280 21848 14280 21876
rect 14274 21836 14280 21848
rect 14332 21836 14338 21888
rect 18598 21876 18604 21888
rect 18559 21848 18604 21876
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19242 21876 19248 21888
rect 19203 21848 19248 21876
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2041 21675 2099 21681
rect 2041 21641 2053 21675
rect 2087 21672 2099 21675
rect 2866 21672 2872 21684
rect 2087 21644 2872 21672
rect 2087 21641 2099 21644
rect 2041 21635 2099 21641
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 8846 21672 8852 21684
rect 4212 21644 4257 21672
rect 8807 21644 8852 21672
rect 4212 21632 4218 21644
rect 8846 21632 8852 21644
rect 8904 21632 8910 21684
rect 12575 21675 12633 21681
rect 12575 21641 12587 21675
rect 12621 21672 12633 21675
rect 12710 21672 12716 21684
rect 12621 21644 12716 21672
rect 12621 21641 12633 21644
rect 12575 21635 12633 21641
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 12989 21675 13047 21681
rect 12989 21641 13001 21675
rect 13035 21672 13047 21675
rect 17405 21675 17463 21681
rect 13035 21644 17356 21672
rect 13035 21641 13047 21644
rect 12989 21635 13047 21641
rect 2884 21536 2912 21632
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 7708 21576 9352 21604
rect 7708 21564 7714 21576
rect 3602 21536 3608 21548
rect 2884 21508 3372 21536
rect 3563 21508 3608 21536
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 2866 21468 2872 21480
rect 2823 21440 2872 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 2866 21428 2872 21440
rect 2924 21428 2930 21480
rect 3344 21477 3372 21508
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21536 5963 21539
rect 5994 21536 6000 21548
rect 5951 21508 6000 21536
rect 5951 21505 5963 21508
rect 5905 21499 5963 21505
rect 5994 21496 6000 21508
rect 6052 21536 6058 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6052 21508 6561 21536
rect 6052 21496 6058 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 7926 21536 7932 21548
rect 7887 21508 7932 21536
rect 6549 21499 6607 21505
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 9030 21536 9036 21548
rect 8991 21508 9036 21536
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9324 21545 9352 21576
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 11238 21496 11244 21548
rect 11296 21536 11302 21548
rect 11333 21539 11391 21545
rect 11333 21536 11345 21539
rect 11296 21508 11345 21536
rect 11296 21496 11302 21508
rect 11333 21505 11345 21508
rect 11379 21536 11391 21539
rect 11977 21539 12035 21545
rect 11977 21536 11989 21539
rect 11379 21508 11989 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 11977 21505 11989 21508
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 3329 21471 3387 21477
rect 3329 21437 3341 21471
rect 3375 21437 3387 21471
rect 3329 21431 3387 21437
rect 3344 21400 3372 21431
rect 4982 21428 4988 21480
rect 5040 21468 5046 21480
rect 5169 21471 5227 21477
rect 5169 21468 5181 21471
rect 5040 21440 5181 21468
rect 5040 21428 5046 21440
rect 5169 21437 5181 21440
rect 5215 21437 5227 21471
rect 5169 21431 5227 21437
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 7653 21471 7711 21477
rect 7653 21437 7665 21471
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 4709 21403 4767 21409
rect 4709 21400 4721 21403
rect 3344 21372 4721 21400
rect 4709 21369 4721 21372
rect 4755 21400 4767 21403
rect 5534 21400 5540 21412
rect 4755 21372 5540 21400
rect 4755 21369 4767 21372
rect 4709 21363 4767 21369
rect 5534 21360 5540 21372
rect 5592 21400 5598 21412
rect 5644 21400 5672 21431
rect 5592 21372 5672 21400
rect 5592 21360 5598 21372
rect 5718 21360 5724 21412
rect 5776 21400 5782 21412
rect 7285 21403 7343 21409
rect 7285 21400 7297 21403
rect 5776 21372 7297 21400
rect 5776 21360 5782 21372
rect 7285 21369 7297 21372
rect 7331 21400 7343 21403
rect 7668 21400 7696 21431
rect 7742 21428 7748 21480
rect 7800 21468 7806 21480
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7800 21440 7849 21468
rect 7800 21428 7806 21440
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 7837 21431 7895 21437
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21468 8539 21471
rect 8754 21468 8760 21480
rect 8527 21440 8760 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 10060 21440 10517 21468
rect 7331 21372 8524 21400
rect 7331 21369 7343 21372
rect 7285 21363 7343 21369
rect 1673 21335 1731 21341
rect 1673 21301 1685 21335
rect 1719 21332 1731 21335
rect 2222 21332 2228 21344
rect 1719 21304 2228 21332
rect 1719 21301 1731 21304
rect 1673 21295 1731 21301
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 2409 21335 2467 21341
rect 2409 21301 2421 21335
rect 2455 21332 2467 21335
rect 2682 21332 2688 21344
rect 2455 21304 2688 21332
rect 2455 21301 2467 21304
rect 2409 21295 2467 21301
rect 2682 21292 2688 21304
rect 2740 21292 2746 21344
rect 4982 21332 4988 21344
rect 4943 21304 4988 21332
rect 4982 21292 4988 21304
rect 5040 21292 5046 21344
rect 6273 21335 6331 21341
rect 6273 21301 6285 21335
rect 6319 21332 6331 21335
rect 6454 21332 6460 21344
rect 6319 21304 6460 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 6454 21292 6460 21304
rect 6512 21292 6518 21344
rect 8496 21332 8524 21372
rect 8846 21360 8852 21412
rect 8904 21400 8910 21412
rect 9125 21403 9183 21409
rect 9125 21400 9137 21403
rect 8904 21372 9137 21400
rect 8904 21360 8910 21372
rect 9125 21369 9137 21372
rect 9171 21369 9183 21403
rect 9125 21363 9183 21369
rect 10060 21332 10088 21440
rect 10505 21437 10517 21440
rect 10551 21468 10563 21471
rect 10870 21468 10876 21480
rect 10551 21440 10876 21468
rect 10551 21437 10563 21440
rect 10505 21431 10563 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 12504 21471 12562 21477
rect 12504 21437 12516 21471
rect 12550 21468 12562 21471
rect 13004 21468 13032 21635
rect 13538 21564 13544 21616
rect 13596 21604 13602 21616
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 13596 21576 14841 21604
rect 13596 21564 13602 21576
rect 14829 21573 14841 21576
rect 14875 21604 14887 21607
rect 15378 21604 15384 21616
rect 14875 21576 15384 21604
rect 14875 21573 14887 21576
rect 14829 21567 14887 21573
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 17328 21604 17356 21644
rect 17405 21641 17417 21675
rect 17451 21672 17463 21675
rect 17770 21672 17776 21684
rect 17451 21644 17776 21672
rect 17451 21641 17463 21644
rect 17405 21635 17463 21641
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 20070 21672 20076 21684
rect 19983 21644 20076 21672
rect 20070 21632 20076 21644
rect 20128 21672 20134 21684
rect 22278 21672 22284 21684
rect 20128 21644 22284 21672
rect 20128 21632 20134 21644
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 22646 21672 22652 21684
rect 22607 21644 22652 21672
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 19058 21604 19064 21616
rect 17328 21576 19064 21604
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 20346 21604 20352 21616
rect 20307 21576 20352 21604
rect 20346 21564 20352 21576
rect 20404 21564 20410 21616
rect 13998 21536 14004 21548
rect 13959 21508 14004 21536
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 15749 21539 15807 21545
rect 15749 21505 15761 21539
rect 15795 21536 15807 21539
rect 15838 21536 15844 21548
rect 15795 21508 15844 21536
rect 15795 21505 15807 21508
rect 15749 21499 15807 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16482 21496 16488 21548
rect 16540 21536 16546 21548
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 16540 21508 18613 21536
rect 16540 21496 16546 21508
rect 12550 21440 13032 21468
rect 12550 21437 12562 21440
rect 12504 21431 12562 21437
rect 10137 21403 10195 21409
rect 10137 21369 10149 21403
rect 10183 21400 10195 21403
rect 10686 21400 10692 21412
rect 10183 21372 10692 21400
rect 10183 21369 10195 21372
rect 10137 21363 10195 21369
rect 10686 21360 10692 21372
rect 10744 21400 10750 21412
rect 11072 21400 11100 21431
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 15252 21440 15301 21468
rect 15252 21428 15258 21440
rect 15289 21437 15301 21440
rect 15335 21468 15347 21471
rect 15930 21468 15936 21480
rect 15335 21440 15936 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 15930 21428 15936 21440
rect 15988 21468 15994 21480
rect 17034 21468 17040 21480
rect 15988 21440 17040 21468
rect 15988 21428 15994 21440
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 18202 21477 18230 21508
rect 18601 21505 18613 21508
rect 18647 21536 18659 21539
rect 18690 21536 18696 21548
rect 18647 21508 18696 21536
rect 18647 21505 18659 21508
rect 18601 21499 18659 21505
rect 18690 21496 18696 21508
rect 18748 21496 18754 21548
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 19242 21536 19248 21548
rect 19199 21508 19248 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 19242 21496 19248 21508
rect 19300 21536 19306 21548
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 19300 21508 21465 21536
rect 19300 21496 19306 21508
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 18187 21471 18245 21477
rect 18187 21468 18199 21471
rect 18165 21440 18199 21468
rect 18187 21437 18199 21440
rect 18233 21437 18245 21471
rect 18187 21431 18245 21437
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21437 20959 21471
rect 21358 21468 21364 21480
rect 21271 21440 21364 21468
rect 20901 21431 20959 21437
rect 11238 21400 11244 21412
rect 10744 21372 11244 21400
rect 10744 21360 10750 21372
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 13630 21400 13636 21412
rect 13591 21372 13636 21400
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 13725 21403 13783 21409
rect 13725 21369 13737 21403
rect 13771 21400 13783 21403
rect 13814 21400 13820 21412
rect 13771 21372 13820 21400
rect 13771 21369 13783 21372
rect 13725 21363 13783 21369
rect 11698 21332 11704 21344
rect 8496 21304 10088 21332
rect 11611 21304 11704 21332
rect 11698 21292 11704 21304
rect 11756 21332 11762 21344
rect 12250 21332 12256 21344
rect 11756 21304 12256 21332
rect 11756 21292 11762 21304
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 13449 21335 13507 21341
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 13740 21332 13768 21363
rect 13814 21360 13820 21372
rect 13872 21360 13878 21412
rect 15657 21403 15715 21409
rect 15657 21369 15669 21403
rect 15703 21400 15715 21403
rect 16111 21403 16169 21409
rect 16111 21400 16123 21403
rect 15703 21372 16123 21400
rect 15703 21369 15715 21372
rect 15657 21363 15715 21369
rect 16111 21369 16123 21372
rect 16157 21400 16169 21403
rect 17773 21403 17831 21409
rect 17773 21400 17785 21403
rect 16157 21372 17785 21400
rect 16157 21369 16169 21372
rect 16111 21363 16169 21369
rect 17773 21369 17785 21372
rect 17819 21400 17831 21403
rect 17954 21400 17960 21412
rect 17819 21372 17960 21400
rect 17819 21369 17831 21372
rect 17773 21363 17831 21369
rect 17954 21360 17960 21372
rect 18012 21400 18018 21412
rect 19474 21403 19532 21409
rect 18012 21372 19104 21400
rect 18012 21360 18018 21372
rect 16666 21332 16672 21344
rect 13495 21304 13768 21332
rect 16627 21304 16672 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 16666 21292 16672 21304
rect 16724 21292 16730 21344
rect 18279 21335 18337 21341
rect 18279 21301 18291 21335
rect 18325 21332 18337 21335
rect 18414 21332 18420 21344
rect 18325 21304 18420 21332
rect 18325 21301 18337 21304
rect 18279 21295 18337 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 19076 21341 19104 21372
rect 19474 21369 19486 21403
rect 19520 21369 19532 21403
rect 19474 21363 19532 21369
rect 19061 21335 19119 21341
rect 19061 21301 19073 21335
rect 19107 21332 19119 21335
rect 19334 21332 19340 21344
rect 19107 21304 19340 21332
rect 19107 21301 19119 21304
rect 19061 21295 19119 21301
rect 19334 21292 19340 21304
rect 19392 21332 19398 21344
rect 19489 21332 19517 21363
rect 19392 21304 19517 21332
rect 20809 21335 20867 21341
rect 19392 21292 19398 21304
rect 20809 21301 20821 21335
rect 20855 21332 20867 21335
rect 20916 21332 20944 21431
rect 21358 21428 21364 21440
rect 21416 21468 21422 21480
rect 21913 21471 21971 21477
rect 21913 21468 21925 21471
rect 21416 21440 21925 21468
rect 21416 21428 21422 21440
rect 21913 21437 21925 21440
rect 21959 21437 21971 21471
rect 21913 21431 21971 21437
rect 21266 21332 21272 21344
rect 20855 21304 21272 21332
rect 20855 21301 20867 21304
rect 20809 21295 20867 21301
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2222 21128 2228 21140
rect 2183 21100 2228 21128
rect 2222 21088 2228 21100
rect 2280 21128 2286 21140
rect 7926 21128 7932 21140
rect 2280 21100 2728 21128
rect 7887 21100 7932 21128
rect 2280 21088 2286 21100
rect 1946 21060 1952 21072
rect 1479 21032 1952 21060
rect 1479 21001 1507 21032
rect 1946 21020 1952 21032
rect 2004 21020 2010 21072
rect 1464 20995 1522 21001
rect 1464 20961 1476 20995
rect 1510 20961 1522 20995
rect 2406 20992 2412 21004
rect 2367 20964 2412 20992
rect 1464 20955 1522 20961
rect 2406 20952 2412 20964
rect 2464 20952 2470 21004
rect 2498 20952 2504 21004
rect 2556 20992 2562 21004
rect 2700 21001 2728 21100
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 9033 21131 9091 21137
rect 9033 21128 9045 21131
rect 8904 21100 9045 21128
rect 8904 21088 8910 21100
rect 9033 21097 9045 21100
rect 9079 21097 9091 21131
rect 9033 21091 9091 21097
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 9272 21100 9413 21128
rect 9272 21088 9278 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 11330 21128 11336 21140
rect 9401 21091 9459 21097
rect 9600 21100 11336 21128
rect 5537 21063 5595 21069
rect 5537 21060 5549 21063
rect 4172 21032 5549 21060
rect 2685 20995 2743 21001
rect 2556 20964 2601 20992
rect 2556 20952 2562 20964
rect 2685 20961 2697 20995
rect 2731 20961 2743 20995
rect 4062 20992 4068 21004
rect 3975 20964 4068 20992
rect 2685 20955 2743 20961
rect 4062 20952 4068 20964
rect 4120 20992 4126 21004
rect 4172 20992 4200 21032
rect 5537 21029 5549 21032
rect 5583 21029 5595 21063
rect 5537 21023 5595 21029
rect 6733 21063 6791 21069
rect 6733 21029 6745 21063
rect 6779 21060 6791 21063
rect 7006 21060 7012 21072
rect 6779 21032 7012 21060
rect 6779 21029 6791 21032
rect 6733 21023 6791 21029
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 7558 21060 7564 21072
rect 7519 21032 7564 21060
rect 7558 21020 7564 21032
rect 7616 21020 7622 21072
rect 4120 20964 4200 20992
rect 4341 20995 4399 21001
rect 4120 20952 4126 20964
rect 4341 20961 4353 20995
rect 4387 20961 4399 20995
rect 4341 20955 4399 20961
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 5718 20992 5724 21004
rect 4847 20964 5724 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 3697 20927 3755 20933
rect 3697 20893 3709 20927
rect 3743 20924 3755 20927
rect 3878 20924 3884 20936
rect 3743 20896 3884 20924
rect 3743 20893 3755 20896
rect 3697 20887 3755 20893
rect 2682 20816 2688 20868
rect 2740 20856 2746 20868
rect 2884 20856 2912 20887
rect 3878 20884 3884 20896
rect 3936 20924 3942 20936
rect 4356 20924 4384 20955
rect 5718 20952 5724 20964
rect 5776 20952 5782 21004
rect 5880 20995 5938 21001
rect 5880 20961 5892 20995
rect 5926 20992 5938 20995
rect 5994 20992 6000 21004
rect 5926 20964 6000 20992
rect 5926 20961 5938 20964
rect 5880 20955 5938 20961
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 8570 20992 8576 21004
rect 8534 20964 8576 20992
rect 8570 20952 8576 20964
rect 8628 21001 8634 21004
rect 8628 20995 8682 21001
rect 8628 20961 8636 20995
rect 8670 20992 8682 20995
rect 9600 20992 9628 21100
rect 11330 21088 11336 21100
rect 11388 21128 11394 21140
rect 11388 21100 13584 21128
rect 11388 21088 11394 21100
rect 9858 21060 9864 21072
rect 9819 21032 9864 21060
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 13259 21063 13317 21069
rect 13259 21029 13271 21063
rect 13305 21060 13317 21063
rect 13446 21060 13452 21072
rect 13305 21032 13452 21060
rect 13305 21029 13317 21032
rect 13259 21023 13317 21029
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 13556 21060 13584 21100
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 13688 21100 14105 21128
rect 13688 21088 13694 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14093 21091 14151 21097
rect 15286 21088 15292 21140
rect 15344 21128 15350 21140
rect 15427 21131 15485 21137
rect 15427 21128 15439 21131
rect 15344 21100 15439 21128
rect 15344 21088 15350 21100
rect 15427 21097 15439 21100
rect 15473 21097 15485 21131
rect 15838 21128 15844 21140
rect 15799 21100 15844 21128
rect 15427 21091 15485 21097
rect 15838 21088 15844 21100
rect 15896 21088 15902 21140
rect 20070 21088 20076 21140
rect 20128 21128 20134 21140
rect 20993 21131 21051 21137
rect 20993 21128 21005 21131
rect 20128 21100 21005 21128
rect 20128 21088 20134 21100
rect 20993 21097 21005 21100
rect 21039 21097 21051 21131
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 20993 21091 21051 21097
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 16482 21060 16488 21072
rect 13556 21032 16488 21060
rect 16482 21020 16488 21032
rect 16540 21020 16546 21072
rect 16666 21020 16672 21072
rect 16724 21060 16730 21072
rect 16761 21063 16819 21069
rect 16761 21060 16773 21063
rect 16724 21032 16773 21060
rect 16724 21020 16730 21032
rect 16761 21029 16773 21032
rect 16807 21060 16819 21063
rect 17126 21060 17132 21072
rect 16807 21032 17132 21060
rect 16807 21029 16819 21032
rect 16761 21023 16819 21029
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 18693 21063 18751 21069
rect 18693 21060 18705 21063
rect 18656 21032 18705 21060
rect 18656 21020 18662 21032
rect 18693 21029 18705 21032
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 8670 20964 9628 20992
rect 8670 20961 8682 20964
rect 8628 20955 8682 20961
rect 8628 20952 8634 20955
rect 11146 20952 11152 21004
rect 11204 20992 11210 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 11204 20964 11253 20992
rect 11204 20952 11210 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 11701 20995 11759 21001
rect 11701 20992 11713 20995
rect 11388 20964 11713 20992
rect 11388 20952 11394 20964
rect 11701 20961 11713 20964
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 15378 21001 15384 21004
rect 15356 20995 15384 21001
rect 15356 20992 15368 20995
rect 13872 20964 13917 20992
rect 15291 20964 15368 20992
rect 13872 20952 13878 20964
rect 15356 20961 15368 20964
rect 15436 20992 15442 21004
rect 15746 20992 15752 21004
rect 15436 20964 15752 20992
rect 15356 20955 15384 20961
rect 15378 20952 15384 20955
rect 15436 20952 15442 20964
rect 15746 20952 15752 20964
rect 15804 20952 15810 21004
rect 21177 20995 21235 21001
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 21266 20992 21272 21004
rect 21223 20964 21272 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 21361 20995 21419 21001
rect 21361 20961 21373 20995
rect 21407 20961 21419 20995
rect 22462 20992 22468 21004
rect 22423 20964 22468 20992
rect 21361 20955 21419 20961
rect 3936 20896 4384 20924
rect 6917 20927 6975 20933
rect 3936 20884 3942 20896
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 7650 20924 7656 20936
rect 6963 20896 7656 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 8711 20927 8769 20933
rect 8711 20893 8723 20927
rect 8757 20924 8769 20927
rect 9398 20924 9404 20936
rect 8757 20896 9404 20924
rect 8757 20893 8769 20896
rect 8711 20887 8769 20893
rect 9398 20884 9404 20896
rect 9456 20924 9462 20936
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 9456 20896 9781 20924
rect 9456 20884 9462 20896
rect 9769 20893 9781 20896
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20924 10103 20927
rect 10134 20924 10140 20936
rect 10091 20896 10140 20924
rect 10091 20893 10103 20896
rect 10045 20887 10103 20893
rect 2740 20828 2912 20856
rect 2740 20816 2746 20828
rect 4154 20816 4160 20868
rect 4212 20856 4218 20868
rect 5951 20859 6009 20865
rect 4212 20828 4257 20856
rect 4212 20816 4218 20828
rect 5951 20825 5963 20859
rect 5997 20856 6009 20859
rect 9214 20856 9220 20868
rect 5997 20828 9220 20856
rect 5997 20825 6009 20828
rect 5951 20819 6009 20825
rect 9214 20816 9220 20828
rect 9272 20816 9278 20868
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 2130 20788 2136 20800
rect 1581 20760 2136 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 2130 20748 2136 20760
rect 2188 20748 2194 20800
rect 5261 20791 5319 20797
rect 5261 20757 5273 20791
rect 5307 20788 5319 20791
rect 5534 20788 5540 20800
rect 5307 20760 5540 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 6270 20788 6276 20800
rect 6231 20760 6276 20788
rect 6270 20748 6276 20760
rect 6328 20748 6334 20800
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 10060 20788 10088 20887
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 11977 20927 12035 20933
rect 11977 20893 11989 20927
rect 12023 20924 12035 20927
rect 12434 20924 12440 20936
rect 12023 20896 12440 20924
rect 12023 20893 12035 20896
rect 11977 20887 12035 20893
rect 12434 20884 12440 20896
rect 12492 20884 12498 20936
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20924 12955 20927
rect 13170 20924 13176 20936
rect 12943 20896 13176 20924
rect 12943 20893 12955 20896
rect 12897 20887 12955 20893
rect 13170 20884 13176 20896
rect 13228 20884 13234 20936
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20924 16727 20927
rect 16758 20924 16764 20936
rect 16715 20896 16764 20924
rect 16715 20893 16727 20896
rect 16669 20887 16727 20893
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20893 17003 20927
rect 16945 20887 17003 20893
rect 16574 20816 16580 20868
rect 16632 20856 16638 20868
rect 16960 20856 16988 20887
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 18601 20927 18659 20933
rect 18601 20924 18613 20927
rect 17920 20896 18613 20924
rect 17920 20884 17926 20896
rect 18601 20893 18613 20896
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 18877 20927 18935 20933
rect 18877 20924 18889 20927
rect 18840 20896 18889 20924
rect 18840 20884 18846 20896
rect 18877 20893 18889 20896
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 21376 20924 21404 20955
rect 22462 20952 22468 20964
rect 22520 20952 22526 21004
rect 22603 20995 22661 21001
rect 22603 20961 22615 20995
rect 22649 20992 22661 20995
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 22649 20964 24593 20992
rect 22649 20961 22661 20964
rect 22603 20955 22661 20961
rect 24581 20961 24593 20964
rect 24627 20992 24639 20995
rect 24670 20992 24676 21004
rect 24627 20964 24676 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 21450 20924 21456 20936
rect 19484 20896 21456 20924
rect 19484 20884 19490 20896
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 16632 20828 16988 20856
rect 16632 20816 16638 20828
rect 17034 20816 17040 20868
rect 17092 20856 17098 20868
rect 22738 20856 22744 20868
rect 17092 20828 22744 20856
rect 17092 20816 17098 20828
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 16114 20788 16120 20800
rect 7432 20760 10088 20788
rect 16075 20760 16120 20788
rect 7432 20748 7438 20760
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 20257 20791 20315 20797
rect 20257 20757 20269 20791
rect 20303 20788 20315 20791
rect 20346 20788 20352 20800
rect 20303 20760 20352 20788
rect 20303 20757 20315 20760
rect 20257 20751 20315 20757
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 474 20544 480 20596
rect 532 20584 538 20596
rect 1857 20587 1915 20593
rect 1857 20584 1869 20587
rect 532 20556 1869 20584
rect 532 20544 538 20556
rect 1857 20553 1869 20556
rect 1903 20584 1915 20587
rect 2406 20584 2412 20596
rect 1903 20556 2412 20584
rect 1903 20553 1915 20556
rect 1857 20547 1915 20553
rect 1762 20340 1768 20392
rect 1820 20380 1826 20392
rect 1872 20380 1900 20547
rect 2406 20544 2412 20556
rect 2464 20584 2470 20596
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 2464 20556 3065 20584
rect 2464 20544 2470 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 3329 20587 3387 20593
rect 3329 20584 3341 20587
rect 3099 20556 3341 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3329 20553 3341 20556
rect 3375 20584 3387 20587
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3375 20556 3433 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 4154 20544 4160 20596
rect 4212 20584 4218 20596
rect 4617 20587 4675 20593
rect 4617 20584 4629 20587
rect 4212 20556 4629 20584
rect 4212 20544 4218 20556
rect 4617 20553 4629 20556
rect 4663 20553 4675 20587
rect 4617 20547 4675 20553
rect 7006 20544 7012 20596
rect 7064 20584 7070 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7064 20556 7757 20584
rect 7064 20544 7070 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 8570 20584 8576 20596
rect 8531 20556 8576 20584
rect 7745 20547 7803 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 9677 20587 9735 20593
rect 9677 20553 9689 20587
rect 9723 20584 9735 20587
rect 9858 20584 9864 20596
rect 9723 20556 9864 20584
rect 9723 20553 9735 20556
rect 9677 20547 9735 20553
rect 9858 20544 9864 20556
rect 9916 20584 9922 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 9916 20556 9965 20584
rect 9916 20544 9922 20556
rect 9953 20553 9965 20556
rect 9999 20584 10011 20587
rect 10321 20587 10379 20593
rect 10321 20584 10333 20587
rect 9999 20556 10333 20584
rect 9999 20553 10011 20556
rect 9953 20547 10011 20553
rect 10321 20553 10333 20556
rect 10367 20553 10379 20587
rect 15378 20584 15384 20596
rect 15339 20556 15384 20584
rect 10321 20547 10379 20553
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 5905 20451 5963 20457
rect 2823 20420 5212 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 5184 20392 5212 20420
rect 5905 20417 5917 20451
rect 5951 20448 5963 20451
rect 6270 20448 6276 20460
rect 5951 20420 6276 20448
rect 5951 20417 5963 20420
rect 5905 20411 5963 20417
rect 6270 20408 6276 20420
rect 6328 20448 6334 20460
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 6328 20420 6837 20448
rect 6328 20408 6334 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 6825 20411 6883 20417
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1820 20352 2053 20380
rect 1820 20340 1826 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20349 2191 20383
rect 2133 20343 2191 20349
rect 1394 20272 1400 20324
rect 1452 20312 1458 20324
rect 1946 20312 1952 20324
rect 1452 20284 1952 20312
rect 1452 20272 1458 20284
rect 1946 20272 1952 20284
rect 2004 20312 2010 20324
rect 2148 20312 2176 20343
rect 2222 20340 2228 20392
rect 2280 20380 2286 20392
rect 2317 20383 2375 20389
rect 2317 20380 2329 20383
rect 2280 20352 2329 20380
rect 2280 20340 2286 20352
rect 2317 20349 2329 20352
rect 2363 20349 2375 20383
rect 2317 20343 2375 20349
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20380 3387 20383
rect 3605 20383 3663 20389
rect 3605 20380 3617 20383
rect 3375 20352 3617 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 3605 20349 3617 20352
rect 3651 20349 3663 20383
rect 3605 20343 3663 20349
rect 3694 20340 3700 20392
rect 3752 20380 3758 20392
rect 3878 20380 3884 20392
rect 3752 20352 3797 20380
rect 3839 20352 3884 20380
rect 3752 20340 3758 20352
rect 3878 20340 3884 20352
rect 3936 20380 3942 20392
rect 4985 20383 5043 20389
rect 4985 20380 4997 20383
rect 3936 20352 4997 20380
rect 3936 20340 3942 20352
rect 4985 20349 4997 20352
rect 5031 20349 5043 20383
rect 5166 20380 5172 20392
rect 5127 20352 5172 20380
rect 4985 20343 5043 20349
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5592 20352 5641 20380
rect 5592 20340 5598 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 8297 20383 8355 20389
rect 8297 20349 8309 20383
rect 8343 20380 8355 20383
rect 8662 20380 8668 20392
rect 8343 20352 8668 20380
rect 8343 20349 8355 20352
rect 8297 20343 8355 20349
rect 8662 20340 8668 20352
rect 8720 20380 8726 20392
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 8720 20352 8769 20380
rect 8720 20340 8726 20352
rect 8757 20349 8769 20352
rect 8803 20349 8815 20383
rect 8757 20343 8815 20349
rect 2004 20284 2176 20312
rect 3712 20312 3740 20340
rect 4154 20312 4160 20324
rect 3712 20284 4160 20312
rect 2004 20272 2010 20284
rect 4154 20272 4160 20284
rect 4212 20272 4218 20324
rect 4246 20272 4252 20324
rect 4304 20312 4310 20324
rect 4341 20315 4399 20321
rect 4341 20312 4353 20315
rect 4304 20284 4353 20312
rect 4304 20272 4310 20284
rect 4341 20281 4353 20284
rect 4387 20281 4399 20315
rect 4341 20275 4399 20281
rect 6454 20272 6460 20324
rect 6512 20312 6518 20324
rect 6641 20315 6699 20321
rect 6641 20312 6653 20315
rect 6512 20284 6653 20312
rect 6512 20272 6518 20284
rect 6641 20281 6653 20284
rect 6687 20312 6699 20315
rect 7187 20315 7245 20321
rect 7187 20312 7199 20315
rect 6687 20284 7199 20312
rect 6687 20281 6699 20284
rect 6641 20275 6699 20281
rect 7187 20281 7199 20284
rect 7233 20312 7245 20315
rect 8846 20312 8852 20324
rect 7233 20284 8852 20312
rect 7233 20281 7245 20284
rect 7187 20275 7245 20281
rect 8846 20272 8852 20284
rect 8904 20312 8910 20324
rect 9119 20315 9177 20321
rect 9119 20312 9131 20315
rect 8904 20284 9131 20312
rect 8904 20272 8910 20284
rect 9119 20281 9131 20284
rect 9165 20312 9177 20315
rect 10336 20312 10364 20547
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 17862 20584 17868 20596
rect 17823 20556 17868 20584
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 18417 20587 18475 20593
rect 18417 20553 18429 20587
rect 18463 20584 18475 20587
rect 18598 20584 18604 20596
rect 18463 20556 18604 20584
rect 18463 20553 18475 20556
rect 18417 20547 18475 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19981 20587 20039 20593
rect 19981 20584 19993 20587
rect 19484 20556 19993 20584
rect 19484 20544 19490 20556
rect 19981 20553 19993 20556
rect 20027 20553 20039 20587
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 19981 20547 20039 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 10778 20516 10784 20528
rect 10612 20488 10784 20516
rect 10612 20457 10640 20488
rect 10778 20476 10784 20488
rect 10836 20476 10842 20528
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 11517 20519 11575 20525
rect 11517 20516 11529 20519
rect 11204 20488 11529 20516
rect 11204 20476 11210 20488
rect 11517 20485 11529 20488
rect 11563 20516 11575 20519
rect 13262 20516 13268 20528
rect 11563 20488 13268 20516
rect 11563 20485 11575 20488
rect 11517 20479 11575 20485
rect 13262 20476 13268 20488
rect 13320 20476 13326 20528
rect 13998 20476 14004 20528
rect 14056 20516 14062 20528
rect 14056 20488 14320 20516
rect 14056 20476 14062 20488
rect 10597 20451 10655 20457
rect 10597 20417 10609 20451
rect 10643 20417 10655 20451
rect 10962 20448 10968 20460
rect 10923 20420 10968 20448
rect 10597 20411 10655 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 12434 20448 12440 20460
rect 12395 20420 12440 20448
rect 12434 20408 12440 20420
rect 12492 20408 12498 20460
rect 14292 20457 14320 20488
rect 16114 20476 16120 20528
rect 16172 20516 16178 20528
rect 17586 20516 17592 20528
rect 16172 20488 17592 20516
rect 16172 20476 16178 20488
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20448 14335 20451
rect 14366 20448 14372 20460
rect 14323 20420 14372 20448
rect 14323 20417 14335 20420
rect 14277 20411 14335 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 16224 20457 16252 20488
rect 17586 20476 17592 20488
rect 17644 20476 17650 20528
rect 18506 20476 18512 20528
rect 18564 20516 18570 20528
rect 19153 20519 19211 20525
rect 19153 20516 19165 20519
rect 18564 20488 19165 20516
rect 18564 20476 18570 20488
rect 19153 20485 19165 20488
rect 19199 20516 19211 20519
rect 19199 20488 20300 20516
rect 19199 20485 19211 20488
rect 19153 20479 19211 20485
rect 20272 20460 20300 20488
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 14516 20420 14565 20448
rect 14516 20408 14522 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20417 16267 20451
rect 16574 20448 16580 20460
rect 16535 20420 16580 20448
rect 16209 20411 16267 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 18601 20451 18659 20457
rect 18601 20448 18613 20451
rect 18472 20420 18613 20448
rect 18472 20408 18478 20420
rect 18601 20417 18613 20420
rect 18647 20448 18659 20451
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 18647 20420 19533 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 20254 20448 20260 20460
rect 20167 20420 20260 20448
rect 19521 20411 19579 20417
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 21266 20448 21272 20460
rect 21179 20420 21272 20448
rect 21266 20408 21272 20420
rect 21324 20448 21330 20460
rect 21545 20451 21603 20457
rect 21545 20448 21557 20451
rect 21324 20420 21557 20448
rect 21324 20408 21330 20420
rect 21545 20417 21557 20420
rect 21591 20448 21603 20451
rect 22830 20448 22836 20460
rect 21591 20420 22836 20448
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 21744 20389 21772 20420
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 13357 20383 13415 20389
rect 13357 20349 13369 20383
rect 13403 20380 13415 20383
rect 14001 20383 14059 20389
rect 14001 20380 14013 20383
rect 13403 20352 14013 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 14001 20349 14013 20352
rect 14047 20349 14059 20383
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21707 20352 21741 20380
rect 14001 20343 14059 20349
rect 21729 20349 21741 20352
rect 21775 20349 21787 20383
rect 21729 20343 21787 20349
rect 10689 20315 10747 20321
rect 10689 20312 10701 20315
rect 9165 20284 10272 20312
rect 10336 20284 10701 20312
rect 9165 20281 9177 20284
rect 9119 20275 9177 20281
rect 2406 20204 2412 20256
rect 2464 20244 2470 20256
rect 4062 20244 4068 20256
rect 2464 20216 4068 20244
rect 2464 20204 2470 20216
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 6270 20244 6276 20256
rect 6052 20216 6276 20244
rect 6052 20204 6058 20216
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 10244 20244 10272 20284
rect 10689 20281 10701 20284
rect 10735 20281 10747 20315
rect 12758 20315 12816 20321
rect 12758 20312 12770 20315
rect 10689 20275 10747 20281
rect 12268 20284 12770 20312
rect 12268 20256 12296 20284
rect 12758 20281 12770 20284
rect 12804 20281 12816 20315
rect 12758 20275 12816 20281
rect 12250 20244 12256 20256
rect 10244 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13504 20216 13645 20244
rect 13504 20204 13510 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 14016 20244 14044 20343
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 22189 20383 22247 20389
rect 22189 20380 22201 20383
rect 22060 20352 22201 20380
rect 22060 20340 22066 20352
rect 22189 20349 22201 20352
rect 22235 20349 22247 20383
rect 22189 20343 22247 20349
rect 14369 20315 14427 20321
rect 14369 20281 14381 20315
rect 14415 20281 14427 20315
rect 14369 20275 14427 20281
rect 16301 20315 16359 20321
rect 16301 20281 16313 20315
rect 16347 20281 16359 20315
rect 16301 20275 16359 20281
rect 14384 20244 14412 20275
rect 14016 20216 14412 20244
rect 16025 20247 16083 20253
rect 13633 20207 13691 20213
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 16316 20244 16344 20275
rect 18690 20272 18696 20324
rect 18748 20312 18754 20324
rect 18748 20284 18793 20312
rect 18748 20272 18754 20284
rect 20346 20272 20352 20324
rect 20404 20312 20410 20324
rect 20901 20315 20959 20321
rect 20404 20284 20449 20312
rect 20404 20272 20410 20284
rect 20901 20281 20913 20315
rect 20947 20312 20959 20315
rect 21266 20312 21272 20324
rect 20947 20284 21272 20312
rect 20947 20281 20959 20284
rect 20901 20275 20959 20281
rect 21266 20272 21272 20284
rect 21324 20312 21330 20324
rect 22462 20312 22468 20324
rect 21324 20284 22468 20312
rect 21324 20272 21330 20284
rect 22462 20272 22468 20284
rect 22520 20312 22526 20324
rect 22741 20315 22799 20321
rect 22741 20312 22753 20315
rect 22520 20284 22753 20312
rect 22520 20272 22526 20284
rect 22741 20281 22753 20284
rect 22787 20281 22799 20315
rect 22741 20275 22799 20281
rect 16390 20244 16396 20256
rect 16071 20216 16396 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 21818 20244 21824 20256
rect 21779 20216 21824 20244
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2041 20043 2099 20049
rect 2041 20040 2053 20043
rect 2004 20012 2053 20040
rect 2004 20000 2010 20012
rect 2041 20009 2053 20012
rect 2087 20009 2099 20043
rect 2041 20003 2099 20009
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1486 19904 1492 19916
rect 1443 19876 1492 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1486 19864 1492 19876
rect 1544 19864 1550 19916
rect 2056 19780 2084 20003
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 2188 20012 6193 20040
rect 2188 20000 2194 20012
rect 6181 20009 6193 20012
rect 6227 20040 6239 20043
rect 7098 20040 7104 20052
rect 6227 20012 7104 20040
rect 6227 20009 6239 20012
rect 6181 20003 6239 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8846 20040 8852 20052
rect 8807 20012 8852 20040
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9398 20040 9404 20052
rect 9359 20012 9404 20040
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 10778 20040 10784 20052
rect 10739 20012 10784 20040
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 13078 20040 13084 20052
rect 13039 20012 13084 20040
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13630 20000 13636 20052
rect 13688 20040 13694 20052
rect 14047 20043 14105 20049
rect 14047 20040 14059 20043
rect 13688 20012 14059 20040
rect 13688 20000 13694 20012
rect 14047 20009 14059 20012
rect 14093 20009 14105 20043
rect 14366 20040 14372 20052
rect 14327 20012 14372 20040
rect 14047 20003 14105 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 15105 20043 15163 20049
rect 15105 20009 15117 20043
rect 15151 20040 15163 20043
rect 15654 20040 15660 20052
rect 15151 20012 15660 20040
rect 15151 20009 15163 20012
rect 15105 20003 15163 20009
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16390 20040 16396 20052
rect 16351 20012 16396 20040
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16758 20040 16764 20052
rect 16719 20012 16764 20040
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 18598 20040 18604 20052
rect 18559 20012 18604 20040
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 19426 20040 19432 20052
rect 19387 20012 19432 20040
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 19981 20043 20039 20049
rect 19981 20009 19993 20043
rect 20027 20040 20039 20043
rect 20346 20040 20352 20052
rect 20027 20012 20352 20040
rect 20027 20009 20039 20012
rect 19981 20003 20039 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 22557 20043 22615 20049
rect 22557 20040 22569 20043
rect 20916 20012 22569 20040
rect 3878 19932 3884 19984
rect 3936 19972 3942 19984
rect 3936 19944 4384 19972
rect 3936 19932 3942 19944
rect 4356 19916 4384 19944
rect 6454 19932 6460 19984
rect 6512 19972 6518 19984
rect 6686 19975 6744 19981
rect 6686 19972 6698 19975
rect 6512 19944 6698 19972
rect 6512 19932 6518 19944
rect 6686 19941 6698 19944
rect 6732 19941 6744 19975
rect 6686 19935 6744 19941
rect 9766 19932 9772 19984
rect 9824 19972 9830 19984
rect 9861 19975 9919 19981
rect 9861 19972 9873 19975
rect 9824 19944 9873 19972
rect 9824 19932 9830 19944
rect 9861 19941 9873 19944
rect 9907 19941 9919 19975
rect 9861 19935 9919 19941
rect 10413 19975 10471 19981
rect 10413 19941 10425 19975
rect 10459 19972 10471 19975
rect 10962 19972 10968 19984
rect 10459 19944 10968 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 2406 19904 2412 19916
rect 2367 19876 2412 19904
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2685 19907 2743 19913
rect 2685 19873 2697 19907
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 3786 19904 3792 19916
rect 3191 19876 3792 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 2222 19796 2228 19848
rect 2280 19836 2286 19848
rect 2700 19836 2728 19867
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 4062 19904 4068 19916
rect 4023 19876 4068 19904
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4338 19904 4344 19916
rect 4299 19876 4344 19904
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 2280 19808 2728 19836
rect 4157 19839 4215 19845
rect 2280 19796 2286 19808
rect 4157 19805 4169 19839
rect 4203 19805 4215 19839
rect 4157 19799 4215 19805
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19836 4859 19839
rect 6086 19836 6092 19848
rect 4847 19808 6092 19836
rect 4847 19805 4859 19808
rect 4801 19799 4859 19805
rect 2038 19768 2044 19780
rect 1951 19740 2044 19768
rect 2038 19728 2044 19740
rect 2096 19768 2102 19780
rect 2501 19771 2559 19777
rect 2501 19768 2513 19771
rect 2096 19740 2513 19768
rect 2096 19728 2102 19740
rect 2501 19737 2513 19740
rect 2547 19768 2559 19771
rect 2774 19768 2780 19780
rect 2547 19740 2780 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2774 19728 2780 19740
rect 2832 19768 2838 19780
rect 3605 19771 3663 19777
rect 3605 19768 3617 19771
rect 2832 19740 3617 19768
rect 2832 19728 2838 19740
rect 3605 19737 3617 19740
rect 3651 19768 3663 19771
rect 3694 19768 3700 19780
rect 3651 19740 3700 19768
rect 3651 19737 3663 19740
rect 3605 19731 3663 19737
rect 3694 19728 3700 19740
rect 3752 19728 3758 19780
rect 4172 19768 4200 19799
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6362 19836 6368 19848
rect 6323 19808 6368 19836
rect 6362 19796 6368 19808
rect 6420 19796 6426 19848
rect 8202 19836 8208 19848
rect 8163 19808 8208 19836
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 10042 19836 10048 19848
rect 9815 19808 10048 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 10042 19796 10048 19808
rect 10100 19796 10106 19848
rect 5537 19771 5595 19777
rect 5537 19768 5549 19771
rect 4172 19740 5549 19768
rect 4172 19712 4200 19740
rect 5537 19737 5549 19740
rect 5583 19737 5595 19771
rect 10428 19768 10456 19935
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 12482 19975 12540 19981
rect 12482 19972 12494 19975
rect 12308 19944 12494 19972
rect 12308 19932 12314 19944
rect 12482 19941 12494 19944
rect 12528 19972 12540 19975
rect 13446 19972 13452 19984
rect 12528 19944 13452 19972
rect 12528 19941 12540 19944
rect 12482 19935 12540 19941
rect 13446 19932 13452 19944
rect 13504 19972 13510 19984
rect 15835 19975 15893 19981
rect 15835 19972 15847 19975
rect 13504 19944 15847 19972
rect 13504 19932 13510 19944
rect 15835 19941 15847 19944
rect 15881 19972 15893 19975
rect 16298 19972 16304 19984
rect 15881 19944 16304 19972
rect 15881 19941 15893 19944
rect 15835 19935 15893 19941
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 17402 19972 17408 19984
rect 17363 19944 17408 19972
rect 17402 19932 17408 19944
rect 17460 19932 17466 19984
rect 20916 19972 20944 20012
rect 22557 20009 22569 20012
rect 22603 20009 22615 20043
rect 22557 20003 22615 20009
rect 21082 19972 21088 19984
rect 19673 19944 20944 19972
rect 21043 19944 21088 19972
rect 13976 19907 14034 19913
rect 13976 19873 13988 19907
rect 14022 19904 14034 19907
rect 14274 19904 14280 19916
rect 14022 19876 14280 19904
rect 14022 19873 14034 19876
rect 13976 19867 14034 19873
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 15470 19904 15476 19916
rect 15383 19876 15476 19904
rect 15470 19864 15476 19876
rect 15528 19904 15534 19916
rect 16206 19904 16212 19916
rect 15528 19876 16212 19904
rect 15528 19864 15534 19876
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19904 19027 19907
rect 19242 19904 19248 19916
rect 19015 19876 19248 19904
rect 19015 19873 19027 19876
rect 18969 19867 19027 19873
rect 19242 19864 19248 19876
rect 19300 19904 19306 19916
rect 19673 19904 19701 19944
rect 21082 19932 21088 19944
rect 21140 19932 21146 19984
rect 22002 19972 22008 19984
rect 21963 19944 22008 19972
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 20254 19904 20260 19916
rect 19300 19876 19701 19904
rect 20215 19876 20260 19904
rect 19300 19864 19306 19876
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 22462 19904 22468 19916
rect 22423 19876 22468 19904
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 22830 19864 22836 19916
rect 22888 19904 22894 19916
rect 22925 19907 22983 19913
rect 22925 19904 22937 19907
rect 22888 19876 22937 19904
rect 22888 19864 22894 19876
rect 22925 19873 22937 19876
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 12158 19836 12164 19848
rect 12119 19808 12164 19836
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 17310 19836 17316 19848
rect 17271 19808 17316 19836
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17586 19836 17592 19848
rect 17547 19808 17592 19836
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19805 19119 19839
rect 20990 19836 20996 19848
rect 20951 19808 20996 19836
rect 19061 19799 19119 19805
rect 5537 19731 5595 19737
rect 7944 19740 10456 19768
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 1946 19700 1952 19712
rect 1581 19672 1952 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 2590 19660 2596 19712
rect 2648 19700 2654 19712
rect 4154 19700 4160 19712
rect 2648 19672 4160 19700
rect 2648 19660 2654 19672
rect 4154 19660 4160 19672
rect 4212 19660 4218 19712
rect 5166 19700 5172 19712
rect 5127 19672 5172 19700
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7285 19703 7343 19709
rect 7285 19700 7297 19703
rect 7248 19672 7297 19700
rect 7248 19660 7254 19672
rect 7285 19669 7297 19672
rect 7331 19700 7343 19703
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 7331 19672 7573 19700
rect 7331 19669 7343 19672
rect 7285 19663 7343 19669
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7561 19663 7619 19669
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 7944 19709 7972 19740
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19076 19768 19104 19799
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21266 19836 21272 19848
rect 21227 19808 21272 19836
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 21818 19768 21824 19780
rect 19024 19740 21824 19768
rect 19024 19728 19030 19740
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7708 19672 7941 19700
rect 7708 19660 7714 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 11238 19700 11244 19712
rect 11199 19672 11244 19700
rect 7929 19663 7987 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 13170 19660 13176 19712
rect 13228 19700 13234 19712
rect 13357 19703 13415 19709
rect 13357 19700 13369 19703
rect 13228 19672 13369 19700
rect 13228 19660 13234 19672
rect 13357 19669 13369 19672
rect 13403 19669 13415 19703
rect 13357 19663 13415 19669
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 21358 19700 21364 19712
rect 18472 19672 21364 19700
rect 18472 19660 18478 19672
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1762 19496 1768 19508
rect 1723 19468 1768 19496
rect 1762 19456 1768 19468
rect 1820 19496 1826 19508
rect 3237 19499 3295 19505
rect 3237 19496 3249 19499
rect 1820 19468 3249 19496
rect 1820 19456 1826 19468
rect 2317 19431 2375 19437
rect 2317 19397 2329 19431
rect 2363 19428 2375 19431
rect 2406 19428 2412 19440
rect 2363 19400 2412 19428
rect 2363 19397 2375 19400
rect 2317 19391 2375 19397
rect 2406 19388 2412 19400
rect 2464 19388 2470 19440
rect 2516 19301 2544 19468
rect 3237 19465 3249 19468
rect 3283 19465 3295 19499
rect 3237 19459 3295 19465
rect 2774 19388 2780 19440
rect 2832 19428 2838 19440
rect 2869 19431 2927 19437
rect 2869 19428 2881 19431
rect 2832 19400 2881 19428
rect 2832 19388 2838 19400
rect 2869 19397 2881 19400
rect 2915 19397 2927 19431
rect 2869 19391 2927 19397
rect 2501 19295 2559 19301
rect 2501 19261 2513 19295
rect 2547 19261 2559 19295
rect 3252 19292 3280 19459
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4246 19496 4252 19508
rect 4028 19468 4252 19496
rect 4028 19456 4034 19468
rect 4246 19456 4252 19468
rect 4304 19496 4310 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 4304 19468 4997 19496
rect 4304 19456 4310 19468
rect 4985 19465 4997 19468
rect 5031 19465 5043 19499
rect 4985 19459 5043 19465
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 6144 19468 8401 19496
rect 6144 19456 6150 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 8389 19459 8447 19465
rect 6454 19428 6460 19440
rect 6415 19400 6460 19428
rect 6454 19388 6460 19400
rect 6512 19388 6518 19440
rect 7098 19360 7104 19372
rect 7059 19332 7104 19360
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 7374 19360 7380 19372
rect 7335 19332 7380 19360
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 8404 19360 8432 19459
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16899 19499 16957 19505
rect 16899 19496 16911 19499
rect 16715 19468 16911 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16899 19465 16911 19468
rect 16945 19496 16957 19499
rect 17310 19496 17316 19508
rect 16945 19468 17316 19496
rect 16945 19465 16957 19468
rect 16899 19459 16957 19465
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 17402 19456 17408 19508
rect 17460 19496 17466 19508
rect 17589 19499 17647 19505
rect 17589 19496 17601 19499
rect 17460 19468 17601 19496
rect 17460 19456 17466 19468
rect 17589 19465 17601 19468
rect 17635 19465 17647 19499
rect 17589 19459 17647 19465
rect 17862 19456 17868 19508
rect 17920 19496 17926 19508
rect 18279 19499 18337 19505
rect 18279 19496 18291 19499
rect 17920 19468 18291 19496
rect 17920 19456 17926 19468
rect 18279 19465 18291 19468
rect 18325 19465 18337 19499
rect 18279 19459 18337 19465
rect 20257 19499 20315 19505
rect 20257 19465 20269 19499
rect 20303 19496 20315 19499
rect 20622 19496 20628 19508
rect 20303 19468 20628 19496
rect 20303 19465 20315 19468
rect 20257 19459 20315 19465
rect 20622 19456 20628 19468
rect 20680 19496 20686 19508
rect 21082 19496 21088 19508
rect 20680 19468 21088 19496
rect 20680 19456 20686 19468
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 14458 19428 14464 19440
rect 8628 19400 14464 19428
rect 8628 19388 8634 19400
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15838 19388 15844 19440
rect 15896 19428 15902 19440
rect 15933 19431 15991 19437
rect 15933 19428 15945 19431
rect 15896 19400 15945 19428
rect 15896 19388 15902 19400
rect 15933 19397 15945 19400
rect 15979 19428 15991 19431
rect 17420 19428 17448 19456
rect 15979 19400 17448 19428
rect 15979 19397 15991 19400
rect 15933 19391 15991 19397
rect 18782 19388 18788 19440
rect 18840 19428 18846 19440
rect 18840 19400 21220 19428
rect 18840 19388 18846 19400
rect 21192 19372 21220 19400
rect 11793 19363 11851 19369
rect 11793 19360 11805 19363
rect 8404 19332 11100 19360
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3252 19264 3433 19292
rect 2501 19255 2559 19261
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3421 19255 3479 19261
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3559 19264 3648 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3620 19224 3648 19264
rect 3694 19252 3700 19304
rect 3752 19292 3758 19304
rect 4338 19292 4344 19304
rect 3752 19264 4344 19292
rect 3752 19252 3758 19264
rect 4338 19252 4344 19264
rect 4396 19292 4402 19304
rect 4433 19295 4491 19301
rect 4433 19292 4445 19295
rect 4396 19264 4445 19292
rect 4396 19252 4402 19264
rect 4433 19261 4445 19264
rect 4479 19261 4491 19295
rect 5442 19292 5448 19304
rect 5403 19264 5448 19292
rect 4433 19255 4491 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 5905 19295 5963 19301
rect 5905 19261 5917 19295
rect 5951 19292 5963 19295
rect 6362 19292 6368 19304
rect 5951 19264 6368 19292
rect 5951 19261 5963 19264
rect 5905 19255 5963 19261
rect 4154 19224 4160 19236
rect 3620 19196 4160 19224
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 5534 19224 5540 19236
rect 5040 19196 5540 19224
rect 5040 19184 5046 19196
rect 5534 19184 5540 19196
rect 5592 19224 5598 19236
rect 5644 19224 5672 19255
rect 6362 19252 6368 19264
rect 6420 19252 6426 19304
rect 8404 19292 8432 19332
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8404 19264 8585 19292
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19261 10839 19295
rect 10781 19255 10839 19261
rect 5592 19196 6500 19224
rect 5592 19184 5598 19196
rect 3881 19159 3939 19165
rect 3881 19125 3893 19159
rect 3927 19156 3939 19159
rect 6270 19156 6276 19168
rect 3927 19128 6276 19156
rect 3927 19125 3939 19128
rect 3881 19119 3939 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6472 19156 6500 19196
rect 7190 19184 7196 19236
rect 7248 19224 7254 19236
rect 9048 19224 9076 19255
rect 7248 19196 7293 19224
rect 8036 19196 9076 19224
rect 7248 19184 7254 19196
rect 8036 19165 8064 19196
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 6472 19128 8033 19156
rect 8021 19125 8033 19128
rect 8067 19125 8079 19159
rect 8662 19156 8668 19168
rect 8623 19128 8668 19156
rect 8021 19119 8079 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 10689 19159 10747 19165
rect 10689 19125 10701 19159
rect 10735 19156 10747 19159
rect 10796 19156 10824 19255
rect 11072 19224 11100 19332
rect 11256 19332 11805 19360
rect 11256 19304 11284 19332
rect 11793 19329 11805 19332
rect 11839 19360 11851 19363
rect 13170 19360 13176 19372
rect 11839 19332 12940 19360
rect 13131 19332 13176 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 11238 19292 11244 19304
rect 11199 19264 11244 19292
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 11517 19295 11575 19301
rect 11517 19261 11529 19295
rect 11563 19292 11575 19295
rect 12158 19292 12164 19304
rect 11563 19264 12164 19292
rect 11563 19261 11575 19264
rect 11517 19255 11575 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12912 19301 12940 19332
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 15013 19363 15071 19369
rect 15013 19329 15025 19363
rect 15059 19360 15071 19363
rect 15654 19360 15660 19372
rect 15059 19332 15660 19360
rect 15059 19329 15071 19332
rect 15013 19323 15071 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 17218 19360 17224 19372
rect 17179 19332 17224 19360
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 18598 19360 18604 19372
rect 18559 19332 18604 19360
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19337 19363 19395 19369
rect 19337 19360 19349 19363
rect 19300 19332 19349 19360
rect 19300 19320 19306 19332
rect 19337 19329 19349 19332
rect 19383 19329 19395 19363
rect 21174 19360 21180 19372
rect 21087 19332 21180 19360
rect 19337 19323 19395 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21453 19363 21511 19369
rect 21453 19360 21465 19363
rect 21324 19332 21465 19360
rect 21324 19320 21330 19332
rect 21453 19329 21465 19332
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 14068 19295 14126 19301
rect 14068 19261 14080 19295
rect 14114 19292 14126 19295
rect 14826 19292 14832 19304
rect 14114 19264 14832 19292
rect 14114 19261 14126 19264
rect 14068 19255 14126 19261
rect 11072 19196 12388 19224
rect 10962 19156 10968 19168
rect 10735 19128 10968 19156
rect 10735 19125 10747 19128
rect 10689 19119 10747 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 12124 19128 12173 19156
rect 12124 19116 12130 19128
rect 12161 19125 12173 19128
rect 12207 19156 12219 19159
rect 12250 19156 12256 19168
rect 12207 19128 12256 19156
rect 12207 19125 12219 19128
rect 12161 19119 12219 19125
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12360 19156 12388 19196
rect 12544 19168 12572 19255
rect 14826 19252 14832 19264
rect 14884 19252 14890 19304
rect 16828 19295 16886 19301
rect 16828 19261 16840 19295
rect 16874 19292 16886 19295
rect 17236 19292 17264 19320
rect 16874 19264 17264 19292
rect 18208 19295 18266 19301
rect 16874 19261 16886 19264
rect 16828 19255 16886 19261
rect 18208 19261 18220 19295
rect 18254 19292 18266 19295
rect 18616 19292 18644 19320
rect 18254 19264 18644 19292
rect 18254 19261 18266 19264
rect 18208 19255 18266 19261
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15375 19227 15433 19233
rect 15375 19224 15387 19227
rect 15160 19196 15387 19224
rect 15160 19184 15166 19196
rect 15375 19193 15387 19196
rect 15421 19224 15433 19227
rect 19658 19227 19716 19233
rect 15421 19196 16344 19224
rect 15421 19193 15433 19196
rect 15375 19187 15433 19193
rect 16316 19168 16344 19196
rect 19658 19193 19670 19227
rect 19704 19193 19716 19227
rect 19658 19187 19716 19193
rect 12526 19156 12532 19168
rect 12360 19128 12532 19156
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 14139 19159 14197 19165
rect 14139 19156 14151 19159
rect 13964 19128 14151 19156
rect 13964 19116 13970 19128
rect 14139 19125 14151 19128
rect 14185 19125 14197 19159
rect 14139 19119 14197 19125
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 14461 19159 14519 19165
rect 14461 19156 14473 19159
rect 14332 19128 14473 19156
rect 14332 19116 14338 19128
rect 14461 19125 14473 19128
rect 14507 19125 14519 19159
rect 16298 19156 16304 19168
rect 16211 19128 16304 19156
rect 14461 19119 14519 19125
rect 16298 19116 16304 19128
rect 16356 19156 16362 19168
rect 19242 19156 19248 19168
rect 16356 19128 19248 19156
rect 16356 19116 16362 19128
rect 19242 19116 19248 19128
rect 19300 19156 19306 19168
rect 19426 19156 19432 19168
rect 19300 19128 19432 19156
rect 19300 19116 19306 19128
rect 19426 19116 19432 19128
rect 19484 19156 19490 19168
rect 19673 19156 19701 19187
rect 21266 19184 21272 19236
rect 21324 19224 21330 19236
rect 21324 19196 21369 19224
rect 21324 19184 21330 19196
rect 22370 19184 22376 19236
rect 22428 19224 22434 19236
rect 22830 19224 22836 19236
rect 22428 19196 22836 19224
rect 22428 19184 22434 19196
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 19484 19128 20545 19156
rect 19484 19116 19490 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 20990 19156 20996 19168
rect 20951 19128 20996 19156
rect 20533 19119 20591 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21284 19156 21312 19184
rect 22097 19159 22155 19165
rect 22097 19156 22109 19159
rect 21284 19128 22109 19156
rect 22097 19125 22109 19128
rect 22143 19125 22155 19159
rect 22462 19156 22468 19168
rect 22423 19128 22468 19156
rect 22097 19119 22155 19125
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 23658 19156 23664 19168
rect 23619 19128 23664 19156
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 106 18912 112 18964
rect 164 18952 170 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 164 18924 5825 18952
rect 164 18912 170 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 6362 18952 6368 18964
rect 6323 18924 6368 18952
rect 5813 18915 5871 18921
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 7745 18955 7803 18961
rect 7745 18952 7757 18955
rect 7708 18924 7757 18952
rect 7708 18912 7714 18924
rect 7745 18921 7757 18924
rect 7791 18921 7803 18955
rect 7745 18915 7803 18921
rect 7926 18912 7932 18964
rect 7984 18952 7990 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 7984 18924 8401 18952
rect 7984 18912 7990 18924
rect 8389 18921 8401 18924
rect 8435 18952 8447 18955
rect 8478 18952 8484 18964
rect 8435 18924 8484 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9214 18912 9220 18964
rect 9272 18952 9278 18964
rect 9401 18955 9459 18961
rect 9401 18952 9413 18955
rect 9272 18924 9413 18952
rect 9272 18912 9278 18924
rect 9401 18921 9413 18924
rect 9447 18952 9459 18955
rect 10042 18952 10048 18964
rect 9447 18924 10048 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12805 18955 12863 18961
rect 12805 18952 12817 18955
rect 12216 18924 12817 18952
rect 12216 18912 12222 18924
rect 12805 18921 12817 18924
rect 12851 18921 12863 18955
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 12805 18915 12863 18921
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 18506 18952 18512 18964
rect 15672 18924 18512 18952
rect 2590 18884 2596 18896
rect 2503 18856 2596 18884
rect 2406 18816 2412 18828
rect 2367 18788 2412 18816
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2516 18825 2544 18856
rect 2590 18844 2596 18856
rect 2648 18884 2654 18896
rect 3881 18887 3939 18893
rect 3881 18884 3893 18887
rect 2648 18856 3893 18884
rect 2648 18844 2654 18856
rect 3881 18853 3893 18856
rect 3927 18884 3939 18887
rect 4246 18884 4252 18896
rect 3927 18856 4252 18884
rect 3927 18853 3939 18856
rect 3881 18847 3939 18853
rect 4246 18844 4252 18856
rect 4304 18844 4310 18896
rect 7101 18887 7159 18893
rect 7101 18853 7113 18887
rect 7147 18884 7159 18887
rect 7190 18884 7196 18896
rect 7147 18856 7196 18884
rect 7147 18853 7159 18856
rect 7101 18847 7159 18853
rect 7190 18844 7196 18856
rect 7248 18884 7254 18896
rect 7834 18884 7840 18896
rect 7248 18856 7840 18884
rect 7248 18844 7254 18856
rect 7834 18844 7840 18856
rect 7892 18844 7898 18896
rect 11603 18887 11661 18893
rect 11603 18853 11615 18887
rect 11649 18884 11661 18887
rect 12066 18884 12072 18896
rect 11649 18856 12072 18884
rect 11649 18853 11661 18856
rect 11603 18847 11661 18853
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 12526 18884 12532 18896
rect 12487 18856 12532 18884
rect 12526 18844 12532 18856
rect 12584 18844 12590 18896
rect 13170 18884 13176 18896
rect 13131 18856 13176 18884
rect 13170 18844 13176 18856
rect 13228 18844 13234 18896
rect 13725 18887 13783 18893
rect 13725 18853 13737 18887
rect 13771 18884 13783 18887
rect 14090 18884 14096 18896
rect 13771 18856 14096 18884
rect 13771 18853 13783 18856
rect 13725 18847 13783 18853
rect 14090 18844 14096 18856
rect 14148 18884 14154 18896
rect 15672 18884 15700 18924
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 18966 18952 18972 18964
rect 18927 18924 18972 18952
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 19981 18955 20039 18961
rect 19981 18921 19993 18955
rect 20027 18952 20039 18955
rect 20622 18952 20628 18964
rect 20027 18924 20392 18952
rect 20583 18924 20628 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 15838 18884 15844 18896
rect 14148 18856 15700 18884
rect 15799 18856 15844 18884
rect 14148 18844 14154 18856
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 17402 18884 17408 18896
rect 17363 18856 17408 18884
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 19382 18887 19440 18893
rect 19382 18884 19394 18887
rect 19300 18856 19394 18884
rect 19300 18844 19306 18856
rect 19382 18853 19394 18856
rect 19428 18853 19440 18887
rect 20364 18884 20392 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 23658 18952 23664 18964
rect 21048 18924 23664 18952
rect 21048 18912 21054 18924
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 21082 18884 21088 18896
rect 20364 18856 21088 18884
rect 19382 18847 19440 18853
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 21174 18844 21180 18896
rect 21232 18884 21238 18896
rect 21913 18887 21971 18893
rect 21913 18884 21925 18887
rect 21232 18856 21925 18884
rect 21232 18844 21238 18856
rect 21913 18853 21925 18856
rect 21959 18853 21971 18887
rect 21913 18847 21971 18853
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18785 2559 18819
rect 2682 18816 2688 18828
rect 2643 18788 2688 18816
rect 2501 18779 2559 18785
rect 2682 18776 2688 18788
rect 2740 18776 2746 18828
rect 3694 18816 3700 18828
rect 3607 18788 3700 18816
rect 3694 18776 3700 18788
rect 3752 18816 3758 18828
rect 4157 18819 4215 18825
rect 4157 18816 4169 18819
rect 3752 18788 4169 18816
rect 3752 18776 3758 18788
rect 4157 18785 4169 18788
rect 4203 18785 4215 18819
rect 4157 18779 4215 18785
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 5629 18819 5687 18825
rect 5629 18816 5641 18819
rect 4948 18788 5641 18816
rect 4948 18776 4954 18788
rect 5629 18785 5641 18788
rect 5675 18816 5687 18819
rect 6086 18816 6092 18828
rect 5675 18788 6092 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 8608 18819 8666 18825
rect 8608 18785 8620 18819
rect 8654 18785 8666 18819
rect 9766 18816 9772 18828
rect 9727 18788 9772 18816
rect 8608 18779 8666 18785
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 3326 18708 3332 18760
rect 3384 18748 3390 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3384 18720 4077 18748
rect 3384 18708 3390 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 5442 18708 5448 18760
rect 5500 18748 5506 18760
rect 7006 18748 7012 18760
rect 5500 18720 5948 18748
rect 6967 18720 7012 18748
rect 5500 18708 5506 18720
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 2317 18683 2375 18689
rect 2317 18680 2329 18683
rect 2280 18652 2329 18680
rect 2280 18640 2286 18652
rect 2317 18649 2329 18652
rect 2363 18680 2375 18683
rect 2682 18680 2688 18692
rect 2363 18652 2688 18680
rect 2363 18649 2375 18652
rect 2317 18643 2375 18649
rect 2682 18640 2688 18652
rect 2740 18680 2746 18692
rect 3344 18680 3372 18708
rect 2740 18652 3372 18680
rect 5920 18680 5948 18720
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 8623 18748 8651 18779
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 10137 18819 10195 18825
rect 10137 18785 10149 18819
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 9398 18748 9404 18760
rect 7524 18720 9404 18748
rect 7524 18708 7530 18720
rect 7944 18692 7972 18720
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 10152 18748 10180 18779
rect 22370 18776 22376 18828
rect 22428 18816 22434 18828
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 22428 18788 22477 18816
rect 22428 18776 22434 18788
rect 22465 18785 22477 18788
rect 22511 18785 22523 18819
rect 22465 18779 22523 18785
rect 22830 18776 22836 18828
rect 22888 18816 22894 18828
rect 22925 18819 22983 18825
rect 22925 18816 22937 18819
rect 22888 18788 22937 18816
rect 22888 18776 22894 18788
rect 22925 18785 22937 18788
rect 22971 18785 22983 18819
rect 22925 18779 22983 18785
rect 24096 18819 24154 18825
rect 24096 18785 24108 18819
rect 24142 18816 24154 18819
rect 24670 18816 24676 18828
rect 24142 18788 24676 18816
rect 24142 18785 24154 18788
rect 24096 18779 24154 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 9548 18720 10180 18748
rect 10413 18751 10471 18757
rect 9548 18708 9554 18720
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10459 18720 11253 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11241 18717 11253 18720
rect 11287 18748 11299 18751
rect 11606 18748 11612 18760
rect 11287 18720 11612 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 13081 18751 13139 18757
rect 13081 18717 13093 18751
rect 13127 18748 13139 18751
rect 13906 18748 13912 18760
rect 13127 18720 13912 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 13906 18708 13912 18720
rect 13964 18708 13970 18760
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 15102 18748 15108 18760
rect 14884 18720 15108 18748
rect 14884 18708 14890 18720
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15749 18751 15807 18757
rect 15749 18717 15761 18751
rect 15795 18717 15807 18751
rect 16206 18748 16212 18760
rect 16167 18720 16212 18748
rect 15749 18711 15807 18717
rect 7650 18680 7656 18692
rect 5920 18652 7656 18680
rect 2740 18640 2746 18652
rect 7650 18640 7656 18652
rect 7708 18640 7714 18692
rect 7926 18640 7932 18692
rect 7984 18640 7990 18692
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 15764 18680 15792 18711
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 17310 18748 17316 18760
rect 17271 18720 17316 18748
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 17586 18748 17592 18760
rect 17547 18720 17592 18748
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 19061 18751 19119 18757
rect 19061 18717 19073 18751
rect 19107 18717 19119 18751
rect 19061 18711 19119 18717
rect 16850 18680 16856 18692
rect 9824 18652 15700 18680
rect 15764 18652 16856 18680
rect 9824 18640 9830 18652
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1544 18584 1961 18612
rect 1544 18572 1550 18584
rect 1949 18581 1961 18584
rect 1995 18612 2007 18615
rect 2130 18612 2136 18624
rect 1995 18584 2136 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2130 18572 2136 18584
rect 2188 18572 2194 18624
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3292 18584 3433 18612
rect 3292 18572 3298 18584
rect 3421 18581 3433 18584
rect 3467 18612 3479 18615
rect 3697 18615 3755 18621
rect 3697 18612 3709 18615
rect 3467 18584 3709 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3697 18581 3709 18584
rect 3743 18581 3755 18615
rect 3697 18575 3755 18581
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 5169 18615 5227 18621
rect 5169 18612 5181 18615
rect 5040 18584 5181 18612
rect 5040 18572 5046 18584
rect 5169 18581 5181 18584
rect 5215 18581 5227 18615
rect 5169 18575 5227 18581
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 5500 18584 6745 18612
rect 5500 18572 5506 18584
rect 6733 18581 6745 18584
rect 6779 18581 6791 18615
rect 6733 18575 6791 18581
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 8021 18615 8079 18621
rect 8021 18612 8033 18615
rect 7064 18584 8033 18612
rect 7064 18572 7070 18584
rect 8021 18581 8033 18584
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 8711 18615 8769 18621
rect 8711 18581 8723 18615
rect 8757 18612 8769 18615
rect 8846 18612 8852 18624
rect 8757 18584 8852 18612
rect 8757 18581 8769 18584
rect 8711 18575 8769 18581
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 9030 18612 9036 18624
rect 8991 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 10781 18615 10839 18621
rect 10781 18612 10793 18615
rect 9640 18584 10793 18612
rect 9640 18572 9646 18584
rect 10781 18581 10793 18584
rect 10827 18612 10839 18615
rect 11238 18612 11244 18624
rect 10827 18584 11244 18612
rect 10827 18581 10839 18584
rect 10781 18575 10839 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 12158 18612 12164 18624
rect 12119 18584 12164 18612
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 15672 18612 15700 18652
rect 16850 18640 16856 18652
rect 16908 18640 16914 18692
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 19076 18680 19104 18711
rect 20622 18708 20628 18760
rect 20680 18748 20686 18760
rect 20993 18751 21051 18757
rect 20993 18748 21005 18751
rect 20680 18720 21005 18748
rect 20680 18708 20686 18720
rect 20993 18717 21005 18720
rect 21039 18717 21051 18751
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 20993 18711 21051 18717
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 23017 18751 23075 18757
rect 23017 18748 23029 18751
rect 21560 18720 23029 18748
rect 21560 18680 21588 18720
rect 23017 18717 23029 18720
rect 23063 18717 23075 18751
rect 23017 18711 23075 18717
rect 18932 18652 21588 18680
rect 18932 18640 18938 18652
rect 17494 18612 17500 18624
rect 15672 18584 17500 18612
rect 17494 18572 17500 18584
rect 17552 18612 17558 18624
rect 18322 18612 18328 18624
rect 17552 18584 18328 18612
rect 17552 18572 17558 18584
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 22554 18572 22560 18624
rect 22612 18612 22618 18624
rect 24167 18615 24225 18621
rect 24167 18612 24179 18615
rect 22612 18584 24179 18612
rect 22612 18572 22618 18584
rect 24167 18581 24179 18584
rect 24213 18581 24225 18615
rect 24167 18575 24225 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1673 18411 1731 18417
rect 1673 18377 1685 18411
rect 1719 18408 1731 18411
rect 2590 18408 2596 18420
rect 1719 18380 2596 18408
rect 1719 18377 1731 18380
rect 1673 18371 1731 18377
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 3237 18411 3295 18417
rect 3237 18377 3249 18411
rect 3283 18408 3295 18411
rect 3326 18408 3332 18420
rect 3283 18380 3332 18408
rect 3283 18377 3295 18380
rect 3237 18371 3295 18377
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 5350 18408 5356 18420
rect 4028 18380 5356 18408
rect 4028 18368 4034 18380
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 9398 18408 9404 18420
rect 9359 18380 9404 18408
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 11606 18408 11612 18420
rect 11567 18380 11612 18408
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 13170 18368 13176 18420
rect 13228 18408 13234 18420
rect 13449 18411 13507 18417
rect 13449 18408 13461 18411
rect 13228 18380 13461 18408
rect 13228 18368 13234 18380
rect 13449 18377 13461 18380
rect 13495 18377 13507 18411
rect 13906 18408 13912 18420
rect 13867 18380 13912 18408
rect 13449 18371 13507 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14826 18368 14832 18420
rect 14884 18408 14890 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14884 18380 14933 18408
rect 14884 18368 14890 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 16301 18411 16359 18417
rect 16301 18408 16313 18411
rect 15896 18380 16313 18408
rect 15896 18368 15902 18380
rect 16301 18377 16313 18380
rect 16347 18377 16359 18411
rect 16301 18371 16359 18377
rect 16761 18411 16819 18417
rect 16761 18377 16773 18411
rect 16807 18408 16819 18411
rect 16850 18408 16856 18420
rect 16807 18380 16856 18408
rect 16807 18377 16819 18380
rect 16761 18371 16819 18377
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 17681 18411 17739 18417
rect 17681 18408 17693 18411
rect 17460 18380 17693 18408
rect 17460 18368 17466 18380
rect 17681 18377 17693 18380
rect 17727 18377 17739 18411
rect 17681 18371 17739 18377
rect 20165 18411 20223 18417
rect 20165 18377 20177 18411
rect 20211 18408 20223 18411
rect 21266 18408 21272 18420
rect 20211 18380 21272 18408
rect 20211 18377 20223 18380
rect 20165 18371 20223 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 24581 18411 24639 18417
rect 24581 18377 24593 18411
rect 24627 18408 24639 18411
rect 24670 18408 24676 18420
rect 24627 18380 24676 18408
rect 24627 18377 24639 18380
rect 24581 18371 24639 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 2038 18340 2044 18352
rect 1999 18312 2044 18340
rect 2038 18300 2044 18312
rect 2096 18300 2102 18352
rect 3878 18300 3884 18352
rect 3936 18340 3942 18352
rect 9030 18340 9036 18352
rect 3936 18312 9036 18340
rect 3936 18300 3942 18312
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 16022 18340 16028 18352
rect 9646 18312 11744 18340
rect 15935 18312 16028 18340
rect 2056 18204 2084 18300
rect 8478 18272 8484 18284
rect 8439 18244 8484 18272
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9646 18272 9674 18312
rect 8904 18244 9674 18272
rect 8904 18232 8910 18244
rect 10042 18232 10048 18284
rect 10100 18272 10106 18284
rect 11716 18272 11744 18312
rect 16022 18300 16028 18312
rect 16080 18340 16086 18352
rect 17420 18340 17448 18368
rect 16080 18312 17448 18340
rect 16080 18300 16086 18312
rect 18966 18300 18972 18352
rect 19024 18340 19030 18352
rect 22370 18340 22376 18352
rect 19024 18312 22376 18340
rect 19024 18300 19030 18312
rect 22370 18300 22376 18312
rect 22428 18340 22434 18352
rect 22465 18343 22523 18349
rect 22465 18340 22477 18343
rect 22428 18312 22477 18340
rect 22428 18300 22434 18312
rect 22465 18309 22477 18312
rect 22511 18309 22523 18343
rect 22465 18303 22523 18309
rect 12250 18272 12256 18284
rect 10100 18244 10145 18272
rect 11716 18244 12256 18272
rect 10100 18232 10106 18244
rect 12250 18232 12256 18244
rect 12308 18272 12314 18284
rect 12518 18275 12576 18281
rect 12518 18272 12530 18275
rect 12308 18244 12530 18272
rect 12308 18232 12314 18244
rect 12518 18241 12530 18244
rect 12564 18241 12576 18275
rect 12518 18235 12576 18241
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18272 19303 18275
rect 20070 18272 20076 18284
rect 19291 18244 20076 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 22002 18272 22008 18284
rect 20956 18244 22008 18272
rect 20956 18232 20962 18244
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 23711 18244 24225 18272
rect 2225 18207 2283 18213
rect 2225 18204 2237 18207
rect 2056 18176 2237 18204
rect 2225 18173 2237 18176
rect 2271 18173 2283 18207
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 2225 18167 2283 18173
rect 6564 18176 6837 18204
rect 3878 18096 3884 18148
rect 3936 18136 3942 18148
rect 4065 18139 4123 18145
rect 4065 18136 4077 18139
rect 3936 18108 4077 18136
rect 3936 18096 3942 18108
rect 4065 18105 4077 18108
rect 4111 18105 4123 18139
rect 4065 18099 4123 18105
rect 4154 18096 4160 18148
rect 4212 18136 4218 18148
rect 4709 18139 4767 18145
rect 4212 18108 4257 18136
rect 4212 18096 4218 18108
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 5258 18136 5264 18148
rect 4755 18108 5264 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 3234 18028 3240 18080
rect 3292 18068 3298 18080
rect 3789 18071 3847 18077
rect 3789 18068 3801 18071
rect 3292 18040 3801 18068
rect 3292 18028 3298 18040
rect 3789 18037 3801 18040
rect 3835 18037 3847 18071
rect 3789 18031 3847 18037
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4985 18071 5043 18077
rect 4985 18068 4997 18071
rect 4304 18040 4997 18068
rect 4304 18028 4310 18040
rect 4985 18037 4997 18040
rect 5031 18037 5043 18071
rect 5350 18068 5356 18080
rect 5311 18040 5356 18068
rect 4985 18031 5043 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 5534 18068 5540 18080
rect 5495 18040 5540 18068
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 6086 18068 6092 18080
rect 6047 18040 6092 18068
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6362 18028 6368 18080
rect 6420 18068 6426 18080
rect 6564 18077 6592 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 6914 18164 6920 18216
rect 6972 18204 6978 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6972 18176 7297 18204
rect 6972 18164 6978 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 14052 18207 14110 18213
rect 13228 18176 13273 18204
rect 13228 18164 13234 18176
rect 14052 18173 14064 18207
rect 14098 18204 14110 18207
rect 15102 18204 15108 18216
rect 14098 18176 14504 18204
rect 15063 18176 15108 18204
rect 14098 18173 14110 18176
rect 14052 18167 14110 18173
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 8297 18139 8355 18145
rect 8297 18136 8309 18139
rect 7984 18108 8309 18136
rect 7984 18096 7990 18108
rect 8297 18105 8309 18108
rect 8343 18136 8355 18139
rect 8573 18139 8631 18145
rect 8573 18136 8585 18139
rect 8343 18108 8585 18136
rect 8343 18105 8355 18108
rect 8297 18099 8355 18105
rect 8573 18105 8585 18108
rect 8619 18105 8631 18139
rect 9122 18136 9128 18148
rect 9083 18108 9128 18136
rect 8573 18099 8631 18105
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 6420 18040 6561 18068
rect 6420 18028 6426 18040
rect 6549 18037 6561 18040
rect 6595 18037 6607 18071
rect 7098 18068 7104 18080
rect 7059 18040 7104 18068
rect 6549 18031 6607 18037
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 8588 18068 8616 18099
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 9858 18136 9864 18148
rect 9324 18108 9864 18136
rect 9324 18068 9352 18108
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 10134 18136 10140 18148
rect 10095 18108 10140 18136
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 10686 18136 10692 18148
rect 10647 18108 10692 18136
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 12158 18096 12164 18148
rect 12216 18136 12222 18148
rect 12253 18139 12311 18145
rect 12253 18136 12265 18139
rect 12216 18108 12265 18136
rect 12216 18096 12222 18108
rect 12253 18105 12265 18108
rect 12299 18136 12311 18139
rect 12621 18139 12679 18145
rect 12621 18136 12633 18139
rect 12299 18108 12633 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 12621 18105 12633 18108
rect 12667 18136 12679 18139
rect 13906 18136 13912 18148
rect 12667 18108 13912 18136
rect 12667 18105 12679 18108
rect 12621 18099 12679 18105
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 14476 18080 14504 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 16904 18207 16962 18213
rect 16904 18173 16916 18207
rect 16950 18204 16962 18207
rect 16950 18176 17448 18204
rect 16950 18173 16962 18176
rect 16904 18167 16962 18173
rect 14826 18096 14832 18148
rect 14884 18136 14890 18148
rect 15426 18139 15484 18145
rect 15426 18136 15438 18139
rect 14884 18108 15438 18136
rect 14884 18096 14890 18108
rect 15426 18105 15438 18108
rect 15472 18105 15484 18139
rect 15426 18099 15484 18105
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 16991 18139 17049 18145
rect 16991 18136 17003 18139
rect 15896 18108 17003 18136
rect 15896 18096 15902 18108
rect 16991 18105 17003 18108
rect 17037 18105 17049 18139
rect 16991 18099 17049 18105
rect 9766 18068 9772 18080
rect 8588 18040 9352 18068
rect 9727 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 12066 18068 12072 18080
rect 11379 18040 12072 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 14139 18071 14197 18077
rect 14139 18068 14151 18071
rect 13504 18040 14151 18068
rect 13504 18028 13510 18040
rect 14139 18037 14151 18040
rect 14185 18037 14197 18071
rect 14458 18068 14464 18080
rect 14419 18040 14464 18068
rect 14139 18031 14197 18037
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 17420 18077 17448 18176
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 18268 18207 18326 18213
rect 18268 18204 18280 18207
rect 18104 18176 18280 18204
rect 18104 18164 18110 18176
rect 18268 18173 18280 18176
rect 18314 18204 18326 18207
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 18314 18176 18705 18204
rect 18314 18173 18326 18176
rect 18268 18167 18326 18173
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 19392 18176 19656 18204
rect 19392 18164 19398 18176
rect 18371 18139 18429 18145
rect 18371 18105 18383 18139
rect 18417 18136 18429 18139
rect 19426 18136 19432 18148
rect 18417 18108 19432 18136
rect 18417 18105 18429 18108
rect 18371 18099 18429 18105
rect 19426 18096 19432 18108
rect 19484 18096 19490 18148
rect 19628 18145 19656 18176
rect 23566 18164 23572 18216
rect 23624 18204 23630 18216
rect 23711 18213 23739 18244
rect 24213 18241 24225 18244
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 23696 18207 23754 18213
rect 23696 18204 23708 18207
rect 23624 18176 23708 18204
rect 23624 18164 23630 18176
rect 23696 18173 23708 18176
rect 23742 18173 23754 18207
rect 23696 18167 23754 18173
rect 24118 18164 24124 18216
rect 24176 18204 24182 18216
rect 24708 18207 24766 18213
rect 24708 18204 24720 18207
rect 24176 18176 24720 18204
rect 24176 18164 24182 18176
rect 24708 18173 24720 18176
rect 24754 18204 24766 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24754 18176 25145 18204
rect 24754 18173 24766 18176
rect 24708 18167 24766 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 19607 18139 19665 18145
rect 19607 18105 19619 18139
rect 19653 18136 19665 18139
rect 20441 18139 20499 18145
rect 20441 18136 20453 18139
rect 19653 18108 20453 18136
rect 19653 18105 19665 18108
rect 19607 18099 19665 18105
rect 20441 18105 20453 18108
rect 20487 18105 20499 18139
rect 20441 18099 20499 18105
rect 21177 18139 21235 18145
rect 21177 18105 21189 18139
rect 21223 18105 21235 18139
rect 21177 18099 21235 18105
rect 17405 18071 17463 18077
rect 17405 18037 17417 18071
rect 17451 18068 17463 18071
rect 17494 18068 17500 18080
rect 17451 18040 17500 18068
rect 17451 18037 17463 18040
rect 17405 18031 17463 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 19153 18071 19211 18077
rect 19153 18037 19165 18071
rect 19199 18068 19211 18071
rect 19242 18068 19248 18080
rect 19199 18040 19248 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 19242 18028 19248 18040
rect 19300 18068 19306 18080
rect 19334 18068 19340 18080
rect 19300 18040 19340 18068
rect 19300 18028 19306 18040
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21192 18068 21220 18099
rect 21266 18096 21272 18148
rect 21324 18136 21330 18148
rect 21821 18139 21879 18145
rect 21324 18108 21369 18136
rect 21324 18096 21330 18108
rect 21821 18105 21833 18139
rect 21867 18136 21879 18139
rect 22094 18136 22100 18148
rect 21867 18108 22100 18136
rect 21867 18105 21879 18108
rect 21821 18099 21879 18105
rect 22094 18096 22100 18108
rect 22152 18096 22158 18148
rect 22186 18068 22192 18080
rect 21192 18040 22192 18068
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 22830 18068 22836 18080
rect 22428 18040 22836 18068
rect 22428 18028 22434 18040
rect 22830 18028 22836 18040
rect 22888 18028 22894 18080
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 23799 18071 23857 18077
rect 23799 18068 23811 18071
rect 23256 18040 23811 18068
rect 23256 18028 23262 18040
rect 23799 18037 23811 18040
rect 23845 18037 23857 18071
rect 23799 18031 23857 18037
rect 24578 18028 24584 18080
rect 24636 18068 24642 18080
rect 24811 18071 24869 18077
rect 24811 18068 24823 18071
rect 24636 18040 24823 18068
rect 24636 18028 24642 18040
rect 24811 18037 24823 18040
rect 24857 18037 24869 18071
rect 24811 18031 24869 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1535 17867 1593 17873
rect 1535 17833 1547 17867
rect 1581 17864 1593 17867
rect 3878 17864 3884 17876
rect 1581 17836 3884 17864
rect 1581 17833 1593 17836
rect 1535 17827 1593 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4212 17836 4997 17864
rect 4212 17824 4218 17836
rect 4985 17833 4997 17836
rect 5031 17864 5043 17867
rect 5350 17864 5356 17876
rect 5031 17836 5356 17864
rect 5031 17833 5043 17836
rect 4985 17827 5043 17833
rect 5350 17824 5356 17836
rect 5408 17824 5414 17876
rect 5994 17864 6000 17876
rect 5955 17836 6000 17864
rect 5994 17824 6000 17836
rect 6052 17824 6058 17876
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10100 17836 10701 17864
rect 10100 17824 10106 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 12158 17864 12164 17876
rect 12119 17836 12164 17864
rect 10689 17827 10747 17833
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12676 17836 12725 17864
rect 12676 17824 12682 17836
rect 12713 17833 12725 17836
rect 12759 17864 12771 17867
rect 13078 17864 13084 17876
rect 12759 17836 13084 17864
rect 12759 17833 12771 17836
rect 12713 17827 12771 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 19061 17867 19119 17873
rect 19061 17864 19073 17867
rect 15442 17836 19073 17864
rect 2498 17756 2504 17808
rect 2556 17796 2562 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 2556 17768 3433 17796
rect 2556 17756 2562 17768
rect 3421 17765 3433 17768
rect 3467 17796 3479 17799
rect 3789 17799 3847 17805
rect 3789 17796 3801 17799
rect 3467 17768 3801 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3789 17765 3801 17768
rect 3835 17796 3847 17799
rect 4246 17796 4252 17808
rect 3835 17768 4252 17796
rect 3835 17765 3847 17768
rect 3789 17759 3847 17765
rect 4246 17756 4252 17768
rect 4304 17756 4310 17808
rect 4430 17805 4436 17808
rect 4427 17796 4436 17805
rect 4391 17768 4436 17796
rect 4427 17759 4436 17768
rect 4430 17756 4436 17759
rect 4488 17756 4494 17808
rect 9582 17796 9588 17808
rect 5736 17768 9588 17796
rect 1464 17731 1522 17737
rect 1464 17697 1476 17731
rect 1510 17728 1522 17731
rect 1670 17728 1676 17740
rect 1510 17700 1676 17728
rect 1510 17697 1522 17700
rect 1464 17691 1522 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2682 17728 2688 17740
rect 2643 17700 2688 17728
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17728 2927 17731
rect 5736 17728 5764 17768
rect 9582 17756 9588 17768
rect 9640 17756 9646 17808
rect 9858 17796 9864 17808
rect 9819 17768 9864 17796
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 12250 17756 12256 17808
rect 12308 17796 12314 17808
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12308 17768 13001 17796
rect 12308 17756 12314 17768
rect 12989 17765 13001 17768
rect 13035 17765 13047 17799
rect 13446 17796 13452 17808
rect 13407 17768 13452 17796
rect 12989 17759 13047 17765
rect 13446 17756 13452 17768
rect 13504 17796 13510 17808
rect 13622 17799 13680 17805
rect 13622 17796 13634 17799
rect 13504 17768 13634 17796
rect 13504 17756 13510 17768
rect 13622 17765 13634 17768
rect 13668 17765 13680 17799
rect 13622 17759 13680 17765
rect 13734 17799 13792 17805
rect 13734 17765 13746 17799
rect 13780 17796 13792 17799
rect 13906 17796 13912 17808
rect 13780 17768 13912 17796
rect 13780 17765 13792 17768
rect 13734 17759 13792 17765
rect 13906 17756 13912 17768
rect 13964 17756 13970 17808
rect 14090 17756 14096 17808
rect 14148 17796 14154 17808
rect 14277 17799 14335 17805
rect 14277 17796 14289 17799
rect 14148 17768 14289 17796
rect 14148 17756 14154 17768
rect 14277 17765 14289 17768
rect 14323 17765 14335 17799
rect 14277 17759 14335 17765
rect 2915 17700 5764 17728
rect 5813 17731 5871 17737
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 5813 17697 5825 17731
rect 5859 17728 5871 17731
rect 6270 17728 6276 17740
rect 5859 17700 6276 17728
rect 5859 17697 5871 17700
rect 5813 17691 5871 17697
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 2884 17660 2912 17691
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6549 17731 6607 17737
rect 6549 17697 6561 17731
rect 6595 17728 6607 17731
rect 7098 17728 7104 17740
rect 6595 17700 7104 17728
rect 6595 17697 6607 17700
rect 6549 17691 6607 17697
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8909 17700 9413 17728
rect 2096 17632 2912 17660
rect 3145 17663 3203 17669
rect 2096 17620 2102 17632
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3191 17632 4077 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 4065 17629 4077 17632
rect 4111 17660 4123 17663
rect 5629 17663 5687 17669
rect 5629 17660 5641 17663
rect 4111 17632 5641 17660
rect 4111 17629 4123 17632
rect 4065 17623 4123 17629
rect 5629 17629 5641 17632
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 8018 17660 8024 17672
rect 6420 17632 8024 17660
rect 6420 17620 6426 17632
rect 8018 17620 8024 17632
rect 8076 17660 8082 17672
rect 8909 17660 8937 17700
rect 9401 17697 9413 17700
rect 9447 17728 9459 17731
rect 9490 17728 9496 17740
rect 9447 17700 9496 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 8076 17632 8937 17660
rect 8076 17620 8082 17632
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9364 17632 9781 17660
rect 9364 17620 9370 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 10870 17660 10876 17672
rect 10459 17632 10876 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11572 17632 11805 17660
rect 11572 17620 11578 17632
rect 11793 17629 11805 17632
rect 11839 17660 11851 17663
rect 15442 17660 15470 17836
rect 19061 17833 19073 17836
rect 19107 17833 19119 17867
rect 19061 17827 19119 17833
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 20622 17864 20628 17876
rect 19484 17836 20628 17864
rect 19484 17824 19490 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 21082 17864 21088 17876
rect 21043 17836 21088 17864
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 16022 17796 16028 17808
rect 15983 17768 16028 17796
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 18874 17796 18880 17808
rect 18835 17768 18880 17796
rect 18874 17756 18880 17768
rect 18932 17756 18938 17808
rect 20070 17796 20076 17808
rect 19306 17768 19564 17796
rect 20031 17768 20076 17796
rect 17402 17728 17408 17740
rect 17363 17700 17408 17728
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 17862 17728 17868 17740
rect 17823 17700 17868 17728
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18966 17728 18972 17740
rect 18927 17700 18972 17728
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 15930 17660 15936 17672
rect 11839 17632 15470 17660
rect 15891 17632 15936 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 16132 17632 17969 17660
rect 1946 17552 1952 17604
rect 2004 17592 2010 17604
rect 4246 17592 4252 17604
rect 2004 17564 4252 17592
rect 2004 17552 2010 17564
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 5261 17595 5319 17601
rect 5261 17592 5273 17595
rect 4448 17564 5273 17592
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 2038 17524 2044 17536
rect 1903 17496 2044 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 2038 17484 2044 17496
rect 2096 17524 2102 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 2096 17496 2237 17524
rect 2096 17484 2102 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 2225 17487 2283 17493
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4448 17524 4476 17564
rect 5261 17561 5273 17564
rect 5307 17561 5319 17595
rect 8297 17595 8355 17601
rect 8297 17592 8309 17595
rect 5261 17555 5319 17561
rect 5920 17564 8309 17592
rect 4120 17496 4476 17524
rect 4120 17484 4126 17496
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 5920 17524 5948 17564
rect 8297 17561 8309 17564
rect 8343 17561 8355 17595
rect 8297 17555 8355 17561
rect 15102 17552 15108 17604
rect 15160 17592 15166 17604
rect 15565 17595 15623 17601
rect 15565 17592 15577 17595
rect 15160 17564 15577 17592
rect 15160 17552 15166 17564
rect 15565 17561 15577 17564
rect 15611 17592 15623 17595
rect 16132 17592 16160 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 19306 17660 19334 17768
rect 19536 17737 19564 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 21637 17799 21695 17805
rect 21637 17765 21649 17799
rect 21683 17796 21695 17799
rect 21818 17796 21824 17808
rect 21683 17768 21824 17796
rect 21683 17765 21695 17768
rect 21637 17759 21695 17765
rect 21818 17756 21824 17768
rect 21876 17756 21882 17808
rect 19521 17731 19579 17737
rect 19521 17697 19533 17731
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 18196 17632 19334 17660
rect 19536 17660 19564 17691
rect 22830 17688 22836 17740
rect 22888 17728 22894 17740
rect 23052 17731 23110 17737
rect 23052 17728 23064 17731
rect 22888 17700 23064 17728
rect 22888 17688 22894 17700
rect 23052 17697 23064 17700
rect 23098 17697 23110 17731
rect 23052 17691 23110 17697
rect 24029 17731 24087 17737
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24118 17728 24124 17740
rect 24075 17700 24124 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 24118 17688 24124 17700
rect 24176 17688 24182 17740
rect 20070 17660 20076 17672
rect 19536 17632 20076 17660
rect 18196 17620 18202 17632
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17660 21603 17663
rect 21910 17660 21916 17672
rect 21591 17632 21916 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 23198 17660 23204 17672
rect 22020 17632 23204 17660
rect 15611 17564 16160 17592
rect 15611 17561 15623 17564
rect 15565 17555 15623 17561
rect 16206 17552 16212 17604
rect 16264 17592 16270 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 16264 17564 16497 17592
rect 16264 17552 16270 17564
rect 16485 17561 16497 17564
rect 16531 17592 16543 17595
rect 16853 17595 16911 17601
rect 16853 17592 16865 17595
rect 16531 17564 16865 17592
rect 16531 17561 16543 17564
rect 16485 17555 16543 17561
rect 16853 17561 16865 17564
rect 16899 17561 16911 17595
rect 17310 17592 17316 17604
rect 17223 17564 17316 17592
rect 16853 17555 16911 17561
rect 17310 17552 17316 17564
rect 17368 17592 17374 17604
rect 22020 17592 22048 17632
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 17368 17564 22048 17592
rect 17368 17552 17374 17564
rect 22094 17552 22100 17604
rect 22152 17592 22158 17604
rect 22738 17592 22744 17604
rect 22152 17564 22744 17592
rect 22152 17552 22158 17564
rect 22738 17552 22744 17564
rect 22796 17552 22802 17604
rect 6822 17524 6828 17536
rect 5132 17496 5948 17524
rect 6783 17496 6828 17524
rect 5132 17484 5138 17496
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 8021 17527 8079 17533
rect 8021 17493 8033 17527
rect 8067 17524 8079 17527
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8067 17496 8769 17524
rect 8067 17493 8079 17496
rect 8021 17487 8079 17493
rect 8757 17493 8769 17496
rect 8803 17524 8815 17527
rect 8938 17524 8944 17536
rect 8803 17496 8944 17524
rect 8803 17493 8815 17496
rect 8757 17487 8815 17493
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 13538 17524 13544 17536
rect 10836 17496 13544 17524
rect 10836 17484 10842 17496
rect 13538 17484 13544 17496
rect 13596 17524 13602 17536
rect 14553 17527 14611 17533
rect 14553 17524 14565 17527
rect 13596 17496 14565 17524
rect 13596 17484 13602 17496
rect 14553 17493 14565 17496
rect 14599 17524 14611 17527
rect 14826 17524 14832 17536
rect 14599 17496 14832 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 15013 17527 15071 17533
rect 15013 17493 15025 17527
rect 15059 17524 15071 17527
rect 15930 17524 15936 17536
rect 15059 17496 15936 17524
rect 15059 17493 15071 17496
rect 15013 17487 15071 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 22002 17484 22008 17536
rect 22060 17524 22066 17536
rect 23155 17527 23213 17533
rect 23155 17524 23167 17527
rect 22060 17496 23167 17524
rect 22060 17484 22066 17496
rect 23155 17493 23167 17496
rect 23201 17493 23213 17527
rect 23155 17487 23213 17493
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 24167 17527 24225 17533
rect 24167 17524 24179 17527
rect 23348 17496 24179 17524
rect 23348 17484 23354 17496
rect 24167 17493 24179 17496
rect 24213 17493 24225 17527
rect 24167 17487 24225 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4341 17323 4399 17329
rect 4341 17289 4353 17323
rect 4387 17320 4399 17323
rect 5442 17320 5448 17332
rect 4387 17292 5448 17320
rect 4387 17289 4399 17292
rect 4341 17283 4399 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8573 17323 8631 17329
rect 8573 17320 8585 17323
rect 8260 17292 8585 17320
rect 8260 17280 8266 17292
rect 8573 17289 8585 17292
rect 8619 17320 8631 17323
rect 11514 17320 11520 17332
rect 8619 17292 8892 17320
rect 11475 17292 11520 17320
rect 8619 17289 8631 17292
rect 8573 17283 8631 17289
rect 1394 17212 1400 17264
rect 1452 17252 1458 17264
rect 4985 17255 5043 17261
rect 4985 17252 4997 17255
rect 1452 17224 4997 17252
rect 1452 17212 1458 17224
rect 4985 17221 4997 17224
rect 5031 17252 5043 17255
rect 5031 17224 5304 17252
rect 5031 17221 5043 17224
rect 4985 17215 5043 17221
rect 1670 17184 1676 17196
rect 1583 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17184 1734 17196
rect 3970 17184 3976 17196
rect 1728 17156 3976 17184
rect 1728 17144 1734 17156
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 5276 17193 5304 17224
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5350 17144 5356 17196
rect 5408 17184 5414 17196
rect 5905 17187 5963 17193
rect 5905 17184 5917 17187
rect 5408 17156 5917 17184
rect 5408 17144 5414 17156
rect 5905 17153 5917 17156
rect 5951 17184 5963 17187
rect 8570 17184 8576 17196
rect 5951 17156 8576 17184
rect 5951 17153 5963 17156
rect 5905 17147 5963 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 8864 17193 8892 17292
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 13633 17323 13691 17329
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13906 17320 13912 17332
rect 13679 17292 13912 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16022 17320 16028 17332
rect 15979 17292 16028 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 18322 17320 18328 17332
rect 18283 17292 18328 17320
rect 18322 17280 18328 17292
rect 18380 17320 18386 17332
rect 18966 17320 18972 17332
rect 18380 17292 18972 17320
rect 18380 17280 18386 17292
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22511 17323 22569 17329
rect 22511 17320 22523 17323
rect 22244 17292 22523 17320
rect 22244 17280 22250 17292
rect 22511 17289 22523 17292
rect 22557 17289 22569 17323
rect 22511 17283 22569 17289
rect 13081 17255 13139 17261
rect 13081 17221 13093 17255
rect 13127 17252 13139 17255
rect 13170 17252 13176 17264
rect 13127 17224 13176 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 13170 17212 13176 17224
rect 13228 17212 13234 17264
rect 13262 17212 13268 17264
rect 13320 17252 13326 17264
rect 17773 17255 17831 17261
rect 17773 17252 17785 17255
rect 13320 17224 14504 17252
rect 13320 17212 13326 17224
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 9122 17184 9128 17196
rect 9083 17156 9128 17184
rect 8849 17147 8907 17153
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10008 17156 10425 17184
rect 10008 17144 10014 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10686 17184 10692 17196
rect 10647 17156 10692 17184
rect 10413 17147 10471 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17184 12587 17187
rect 13998 17184 14004 17196
rect 12575 17156 14004 17184
rect 12575 17153 12587 17156
rect 12529 17147 12587 17153
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 2096 17088 2329 17116
rect 2096 17076 2102 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17116 2651 17119
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 2639 17088 3433 17116
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 3421 17085 3433 17088
rect 3467 17116 3479 17119
rect 5074 17116 5080 17128
rect 3467 17088 5080 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7742 17116 7748 17128
rect 7055 17088 7748 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7742 17076 7748 17088
rect 7800 17116 7806 17128
rect 14476 17125 14504 17224
rect 15028 17224 17785 17252
rect 8205 17119 8263 17125
rect 8205 17116 8217 17119
rect 7800 17088 8217 17116
rect 7800 17076 7806 17088
rect 8205 17085 8217 17088
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 14461 17119 14519 17125
rect 14461 17085 14473 17119
rect 14507 17116 14519 17119
rect 14734 17116 14740 17128
rect 14507 17088 14740 17116
rect 14507 17085 14519 17088
rect 14461 17079 14519 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 14826 17076 14832 17128
rect 14884 17116 14890 17128
rect 15028 17125 15056 17224
rect 17773 17221 17785 17224
rect 17819 17252 17831 17255
rect 17862 17252 17868 17264
rect 17819 17224 17868 17252
rect 17819 17221 17831 17224
rect 17773 17215 17831 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 22278 17252 22284 17264
rect 18012 17224 22284 17252
rect 18012 17212 18018 17224
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 24118 17212 24124 17264
rect 24176 17252 24182 17264
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 24176 17224 24501 17252
rect 24176 17212 24182 17224
rect 24489 17221 24501 17224
rect 24535 17221 24547 17255
rect 24489 17215 24547 17221
rect 16574 17184 16580 17196
rect 16535 17156 16580 17184
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17184 18935 17187
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 18923 17156 20177 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 20165 17153 20177 17156
rect 20211 17184 20223 17187
rect 24026 17184 24032 17196
rect 20211 17156 24032 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 14884 17088 15025 17116
rect 14884 17076 14890 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 22278 17076 22284 17128
rect 22336 17116 22342 17128
rect 23750 17125 23756 17128
rect 22408 17119 22466 17125
rect 22408 17116 22420 17119
rect 22336 17088 22420 17116
rect 22336 17076 22342 17088
rect 22408 17085 22420 17088
rect 22454 17085 22466 17119
rect 23728 17119 23756 17125
rect 23728 17116 23740 17119
rect 23663 17088 23740 17116
rect 22408 17079 22466 17085
rect 23728 17085 23740 17088
rect 23808 17116 23814 17128
rect 24121 17119 24179 17125
rect 24121 17116 24133 17119
rect 23808 17088 24133 17116
rect 23728 17079 23756 17085
rect 23750 17076 23756 17079
rect 23808 17076 23814 17088
rect 24121 17085 24133 17088
rect 24167 17085 24179 17119
rect 24121 17079 24179 17085
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 3783 17051 3841 17057
rect 3783 17048 3795 17051
rect 3375 17020 3795 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 3783 17017 3795 17020
rect 3829 17048 3841 17051
rect 5353 17051 5411 17057
rect 3829 17020 4476 17048
rect 3829 17017 3841 17020
rect 3783 17011 3841 17017
rect 4448 16992 4476 17020
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 5442 17048 5448 17060
rect 5399 17020 5448 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 7330 17051 7388 17057
rect 6113 17020 6684 17048
rect 2682 16940 2688 16992
rect 2740 16980 2746 16992
rect 2961 16983 3019 16989
rect 2961 16980 2973 16983
rect 2740 16952 2973 16980
rect 2740 16940 2746 16952
rect 2961 16949 2973 16952
rect 3007 16980 3019 16983
rect 3602 16980 3608 16992
rect 3007 16952 3608 16980
rect 3007 16949 3019 16952
rect 2961 16943 3019 16949
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 4430 16940 4436 16992
rect 4488 16980 4494 16992
rect 4709 16983 4767 16989
rect 4709 16980 4721 16983
rect 4488 16952 4721 16980
rect 4488 16940 4494 16952
rect 4709 16949 4721 16952
rect 4755 16980 4767 16983
rect 6113 16980 6141 17020
rect 6270 16980 6276 16992
rect 4755 16952 6141 16980
rect 6231 16952 6276 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 6270 16940 6276 16952
rect 6328 16940 6334 16992
rect 6656 16989 6684 17020
rect 7330 17017 7342 17051
rect 7376 17048 7388 17051
rect 7466 17048 7472 17060
rect 7376 17020 7472 17048
rect 7376 17017 7388 17020
rect 7330 17011 7388 17017
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 7006 16980 7012 16992
rect 6687 16952 7012 16980
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 7006 16940 7012 16952
rect 7064 16980 7070 16992
rect 7345 16980 7373 17011
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 8938 17048 8944 17060
rect 8899 17020 8944 17048
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17017 10563 17051
rect 10505 17011 10563 17017
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12618 17048 12624 17060
rect 12299 17020 12624 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 7064 16952 7373 16980
rect 8956 16980 8984 17008
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 8956 16952 9781 16980
rect 7064 16940 7070 16952
rect 9769 16949 9781 16952
rect 9815 16980 9827 16983
rect 9858 16980 9864 16992
rect 9815 16952 9864 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 9858 16940 9864 16952
rect 9916 16980 9922 16992
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 9916 16952 10149 16980
rect 9916 16940 9922 16952
rect 10137 16949 10149 16952
rect 10183 16980 10195 16983
rect 10520 16980 10548 17011
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 14918 17008 14924 17060
rect 14976 17048 14982 17060
rect 16206 17048 16212 17060
rect 14976 17020 16212 17048
rect 14976 17008 14982 17020
rect 16206 17008 16212 17020
rect 16264 17008 16270 17060
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 16356 17020 16401 17048
rect 16356 17008 16362 17020
rect 20714 17008 20720 17060
rect 20772 17048 20778 17060
rect 20901 17051 20959 17057
rect 20901 17048 20913 17051
rect 20772 17020 20913 17048
rect 20772 17008 20778 17020
rect 20901 17017 20913 17020
rect 20947 17017 20959 17051
rect 20901 17011 20959 17017
rect 20990 17008 20996 17060
rect 21048 17048 21054 17060
rect 21545 17051 21603 17057
rect 21048 17020 21141 17048
rect 21048 17008 21054 17020
rect 21545 17017 21557 17051
rect 21591 17048 21603 17051
rect 21634 17048 21640 17060
rect 21591 17020 21640 17048
rect 21591 17017 21603 17020
rect 21545 17011 21603 17017
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 10183 16952 10548 16980
rect 11885 16983 11943 16989
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 12158 16980 12164 16992
rect 11931 16952 12164 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 12158 16940 12164 16952
rect 12216 16980 12222 16992
rect 12802 16980 12808 16992
rect 12216 16952 12808 16980
rect 12216 16940 12222 16952
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13998 16980 14004 16992
rect 13959 16952 14004 16980
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14826 16980 14832 16992
rect 14787 16952 14832 16980
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 18785 16983 18843 16989
rect 18785 16980 18797 16983
rect 18695 16952 18797 16980
rect 18785 16949 18797 16952
rect 18831 16980 18843 16983
rect 19242 16980 19248 16992
rect 18831 16952 19248 16980
rect 18831 16949 18843 16952
rect 18785 16943 18843 16949
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 20438 16980 20444 16992
rect 19843 16952 20444 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 20530 16940 20536 16992
rect 20588 16980 20594 16992
rect 20625 16983 20683 16989
rect 20625 16980 20637 16983
rect 20588 16952 20637 16980
rect 20588 16940 20594 16952
rect 20625 16949 20637 16952
rect 20671 16980 20683 16983
rect 21008 16980 21036 17008
rect 21818 16980 21824 16992
rect 20671 16952 21036 16980
rect 21779 16952 21824 16980
rect 20671 16949 20683 16952
rect 20625 16943 20683 16949
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 22830 16940 22836 16992
rect 22888 16980 22894 16992
rect 23017 16983 23075 16989
rect 23017 16980 23029 16983
rect 22888 16952 23029 16980
rect 22888 16940 22894 16952
rect 23017 16949 23029 16952
rect 23063 16949 23075 16983
rect 23017 16943 23075 16949
rect 23198 16940 23204 16992
rect 23256 16980 23262 16992
rect 23799 16983 23857 16989
rect 23799 16980 23811 16983
rect 23256 16952 23811 16980
rect 23256 16940 23262 16952
rect 23799 16949 23811 16952
rect 23845 16949 23857 16983
rect 23799 16943 23857 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 4614 16736 4620 16788
rect 4672 16776 4678 16788
rect 5353 16779 5411 16785
rect 5353 16776 5365 16779
rect 4672 16748 5365 16776
rect 4672 16736 4678 16748
rect 5353 16745 5365 16748
rect 5399 16776 5411 16779
rect 5534 16776 5540 16788
rect 5399 16748 5540 16776
rect 5399 16745 5411 16748
rect 5353 16739 5411 16745
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 7742 16776 7748 16788
rect 7703 16748 7748 16776
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 9364 16748 9413 16776
rect 9364 16736 9370 16748
rect 9401 16745 9413 16748
rect 9447 16745 9459 16779
rect 9401 16739 9459 16745
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10689 16779 10747 16785
rect 10689 16776 10701 16779
rect 10008 16748 10701 16776
rect 10008 16736 10014 16748
rect 10689 16745 10701 16748
rect 10735 16745 10747 16779
rect 10689 16739 10747 16745
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14884 16748 15025 16776
rect 14884 16736 14890 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 5258 16708 5264 16720
rect 2056 16680 5264 16708
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 2056 16640 2084 16680
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 9490 16708 9496 16720
rect 5828 16680 9496 16708
rect 1510 16612 2084 16640
rect 2685 16643 2743 16649
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 2866 16640 2872 16652
rect 2731 16612 2872 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 1946 16572 1952 16584
rect 1859 16544 1952 16572
rect 1946 16532 1952 16544
rect 2004 16572 2010 16584
rect 2498 16572 2504 16584
rect 2004 16544 2504 16572
rect 2004 16532 2010 16544
rect 2498 16532 2504 16544
rect 2556 16572 2562 16584
rect 2700 16572 2728 16603
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 4062 16640 4068 16652
rect 3191 16612 4068 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 2556 16544 2728 16572
rect 2976 16572 3004 16603
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 5828 16640 5856 16680
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 9548 16680 9781 16708
rect 9548 16668 9554 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 9769 16671 9827 16677
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10042 16708 10048 16720
rect 9916 16680 10048 16708
rect 9916 16668 9922 16680
rect 10042 16668 10048 16680
rect 10100 16668 10106 16720
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 13817 16711 13875 16717
rect 13817 16708 13829 16711
rect 13504 16680 13829 16708
rect 13504 16668 13510 16680
rect 13817 16677 13829 16680
rect 13863 16677 13875 16711
rect 13817 16671 13875 16677
rect 14369 16711 14427 16717
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14918 16708 14924 16720
rect 14415 16680 14924 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 5994 16640 6000 16652
rect 4304 16612 5856 16640
rect 5955 16612 6000 16640
rect 4304 16600 4310 16612
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 6144 16612 6377 16640
rect 6144 16600 6150 16612
rect 6365 16609 6377 16612
rect 6411 16640 6423 16643
rect 6822 16640 6828 16652
rect 6411 16612 6828 16640
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7650 16640 7656 16652
rect 7611 16612 7656 16640
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16640 8079 16643
rect 8386 16640 8392 16652
rect 8067 16612 8392 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 12066 16640 12072 16652
rect 11112 16612 12072 16640
rect 11112 16600 11118 16612
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 12618 16640 12624 16652
rect 12579 16612 12624 16640
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 15028 16640 15056 16739
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16776 16451 16779
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16439 16748 16681 16776
rect 16439 16745 16451 16748
rect 16393 16739 16451 16745
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 17920 16748 18061 16776
rect 17920 16736 17926 16748
rect 18049 16745 18061 16748
rect 18095 16745 18107 16779
rect 18049 16739 18107 16745
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 20990 16776 20996 16788
rect 19291 16748 20996 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21910 16776 21916 16788
rect 21871 16748 21916 16776
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 24121 16779 24179 16785
rect 24121 16776 24133 16779
rect 24084 16748 24133 16776
rect 24084 16736 24090 16748
rect 24121 16745 24133 16748
rect 24167 16745 24179 16779
rect 24121 16739 24179 16745
rect 15835 16711 15893 16717
rect 15835 16677 15847 16711
rect 15881 16708 15893 16711
rect 16114 16708 16120 16720
rect 15881 16680 16120 16708
rect 15881 16677 15893 16680
rect 15835 16671 15893 16677
rect 16114 16668 16120 16680
rect 16172 16708 16178 16720
rect 18687 16711 18745 16717
rect 18687 16708 18699 16711
rect 16172 16680 18699 16708
rect 16172 16668 16178 16680
rect 18687 16677 18699 16680
rect 18733 16677 18745 16711
rect 18687 16671 18745 16677
rect 19613 16711 19671 16717
rect 19613 16677 19625 16711
rect 19659 16708 19671 16711
rect 20070 16708 20076 16720
rect 19659 16680 20076 16708
rect 19659 16677 19671 16680
rect 19613 16671 19671 16677
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 20806 16708 20812 16720
rect 20496 16680 20812 16708
rect 20496 16668 20502 16680
rect 20806 16668 20812 16680
rect 20864 16708 20870 16720
rect 21085 16711 21143 16717
rect 21085 16708 21097 16711
rect 20864 16680 21097 16708
rect 20864 16668 20870 16680
rect 21085 16677 21097 16680
rect 21131 16708 21143 16711
rect 21818 16708 21824 16720
rect 21131 16680 21824 16708
rect 21131 16677 21143 16680
rect 21085 16671 21143 16677
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 22554 16708 22560 16720
rect 22515 16680 22560 16708
rect 22554 16668 22560 16680
rect 22612 16668 22618 16720
rect 22646 16668 22652 16720
rect 22704 16708 22710 16720
rect 22704 16680 22749 16708
rect 22704 16668 22710 16680
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15028 16612 15485 16640
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 17218 16640 17224 16652
rect 17179 16612 17224 16640
rect 15473 16603 15531 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 24210 16640 24216 16652
rect 24171 16612 24216 16640
rect 24210 16600 24216 16612
rect 24268 16600 24274 16652
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16609 24547 16643
rect 24489 16603 24547 16609
rect 3878 16572 3884 16584
rect 2976 16544 3884 16572
rect 2556 16532 2562 16544
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 6638 16572 6644 16584
rect 6599 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10870 16572 10876 16584
rect 10459 16544 10876 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 1535 16507 1593 16513
rect 1535 16473 1547 16507
rect 1581 16504 1593 16507
rect 4062 16504 4068 16516
rect 1581 16476 4068 16504
rect 1581 16473 1593 16476
rect 1535 16467 1593 16473
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 4706 16464 4712 16516
rect 4764 16504 4770 16516
rect 4985 16507 5043 16513
rect 4985 16504 4997 16507
rect 4764 16476 4997 16504
rect 4764 16464 4770 16476
rect 4985 16473 4997 16476
rect 5031 16504 5043 16507
rect 5629 16507 5687 16513
rect 5629 16504 5641 16507
rect 5031 16476 5641 16504
rect 5031 16473 5043 16476
rect 4985 16467 5043 16473
rect 5629 16473 5641 16476
rect 5675 16473 5687 16507
rect 5629 16467 5687 16473
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 8294 16504 8300 16516
rect 7800 16476 8300 16504
rect 7800 16464 7806 16476
rect 8294 16464 8300 16476
rect 8352 16464 8358 16516
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 11072 16504 11100 16600
rect 12710 16572 12716 16584
rect 12671 16544 12716 16572
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 13722 16572 13728 16584
rect 13683 16544 13728 16572
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16572 17831 16575
rect 18322 16572 18328 16584
rect 17819 16544 18328 16572
rect 17819 16541 17831 16544
rect 17773 16535 17831 16541
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 20438 16572 20444 16584
rect 19576 16544 20444 16572
rect 19576 16532 19582 16544
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 20982 16575 21040 16581
rect 20982 16572 20994 16575
rect 20916 16544 20994 16572
rect 8536 16476 11100 16504
rect 8536 16464 8542 16476
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 13320 16476 13814 16504
rect 13320 16464 13326 16476
rect 2317 16439 2375 16445
rect 2317 16405 2329 16439
rect 2363 16436 2375 16439
rect 2958 16436 2964 16448
rect 2363 16408 2964 16436
rect 2363 16405 2375 16408
rect 2317 16399 2375 16405
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3108 16408 3433 16436
rect 3108 16396 3114 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 7064 16408 7113 16436
rect 7064 16396 7070 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 7650 16396 7656 16448
rect 7708 16436 7714 16448
rect 8496 16436 8524 16464
rect 7708 16408 8524 16436
rect 8665 16439 8723 16445
rect 7708 16396 7714 16408
rect 8665 16405 8677 16439
rect 8711 16436 8723 16439
rect 8754 16436 8760 16448
rect 8711 16408 8760 16436
rect 8711 16405 8723 16408
rect 8665 16399 8723 16405
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 8938 16436 8944 16448
rect 8899 16408 8944 16436
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13786 16436 13814 16476
rect 17359 16439 17417 16445
rect 17359 16436 17371 16439
rect 13786 16408 17371 16436
rect 17359 16405 17371 16408
rect 17405 16405 17417 16439
rect 20714 16436 20720 16448
rect 20675 16408 20720 16436
rect 17359 16399 17417 16405
rect 20714 16396 20720 16408
rect 20772 16396 20778 16448
rect 20916 16436 20944 16544
rect 20982 16541 20994 16544
rect 21028 16541 21040 16575
rect 21634 16572 21640 16584
rect 21547 16544 21640 16572
rect 20982 16535 21040 16541
rect 21634 16532 21640 16544
rect 21692 16572 21698 16584
rect 22094 16572 22100 16584
rect 21692 16544 22100 16572
rect 21692 16532 21698 16544
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 22738 16532 22744 16584
rect 22796 16572 22802 16584
rect 22833 16575 22891 16581
rect 22833 16572 22845 16575
rect 22796 16544 22845 16572
rect 22796 16532 22802 16544
rect 22833 16541 22845 16544
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24504 16504 24532 16603
rect 24176 16476 24532 16504
rect 24176 16464 24182 16476
rect 20990 16436 20996 16448
rect 20903 16408 20996 16436
rect 20990 16396 20996 16408
rect 21048 16436 21054 16448
rect 23198 16436 23204 16448
rect 21048 16408 23204 16436
rect 21048 16396 21054 16408
rect 23198 16396 23204 16408
rect 23256 16396 23262 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1946 16192 1952 16244
rect 2004 16232 2010 16244
rect 2133 16235 2191 16241
rect 2133 16232 2145 16235
rect 2004 16204 2145 16232
rect 2004 16192 2010 16204
rect 2133 16201 2145 16204
rect 2179 16201 2191 16235
rect 2133 16195 2191 16201
rect 2593 16235 2651 16241
rect 2593 16201 2605 16235
rect 2639 16232 2651 16235
rect 2866 16232 2872 16244
rect 2639 16204 2872 16232
rect 2639 16201 2651 16204
rect 2593 16195 2651 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4430 16232 4436 16244
rect 4203 16204 4436 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4430 16192 4436 16204
rect 4488 16192 4494 16244
rect 8202 16232 8208 16244
rect 7668 16204 8208 16232
rect 5994 16164 6000 16176
rect 5955 16136 6000 16164
rect 5994 16124 6000 16136
rect 6052 16164 6058 16176
rect 7668 16164 7696 16204
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 9858 16232 9864 16244
rect 9815 16204 9864 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 12066 16232 12072 16244
rect 12027 16204 12072 16232
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 12618 16232 12624 16244
rect 12579 16204 12624 16232
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 14090 16232 14096 16244
rect 13228 16204 14096 16232
rect 13228 16192 13234 16204
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 14737 16235 14795 16241
rect 14737 16201 14749 16235
rect 14783 16232 14795 16235
rect 15286 16232 15292 16244
rect 14783 16204 15292 16232
rect 14783 16201 14795 16204
rect 14737 16195 14795 16201
rect 6052 16136 7696 16164
rect 7745 16167 7803 16173
rect 6052 16124 6058 16136
rect 7745 16133 7757 16167
rect 7791 16164 7803 16167
rect 8754 16164 8760 16176
rect 7791 16136 8760 16164
rect 7791 16133 7803 16136
rect 7745 16127 7803 16133
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 12802 16124 12808 16176
rect 12860 16164 12866 16176
rect 14752 16164 14780 16195
rect 15286 16192 15292 16204
rect 15344 16232 15350 16244
rect 16114 16232 16120 16244
rect 15344 16204 16120 16232
rect 15344 16192 15350 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 17218 16232 17224 16244
rect 17179 16204 17224 16232
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 20530 16232 20536 16244
rect 20491 16204 20536 16232
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 24811 16235 24869 16241
rect 24811 16232 24823 16235
rect 20772 16204 24823 16232
rect 20772 16192 20778 16204
rect 24811 16201 24823 16204
rect 24857 16201 24869 16235
rect 24811 16195 24869 16201
rect 16482 16164 16488 16176
rect 12860 16136 14780 16164
rect 16395 16136 16488 16164
rect 12860 16124 12866 16136
rect 16482 16124 16488 16136
rect 16540 16164 16546 16176
rect 17954 16164 17960 16176
rect 16540 16136 17960 16164
rect 16540 16124 16546 16136
rect 1670 16096 1676 16108
rect 1412 16068 1676 16096
rect 1412 16037 1440 16068
rect 1670 16056 1676 16068
rect 1728 16096 1734 16108
rect 8938 16096 8944 16108
rect 1728 16068 8944 16096
rect 1728 16056 1734 16068
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 9122 16096 9128 16108
rect 9083 16068 9128 16096
rect 9122 16056 9128 16068
rect 9180 16096 9186 16108
rect 9950 16096 9956 16108
rect 9180 16068 9956 16096
rect 9180 16056 9186 16068
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13446 16096 13452 16108
rect 13219 16068 13452 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13446 16056 13452 16068
rect 13504 16096 13510 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13504 16068 14289 16096
rect 13504 16056 13510 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 15378 16056 15384 16108
rect 15436 16096 15442 16108
rect 16715 16099 16773 16105
rect 16715 16096 16727 16099
rect 15436 16068 16727 16096
rect 15436 16056 15442 16068
rect 16715 16065 16727 16068
rect 16761 16065 16773 16099
rect 16715 16059 16773 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 2866 16028 2872 16040
rect 2827 16000 2872 16028
rect 1397 15991 1455 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7926 16028 7932 16040
rect 6871 16000 7932 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8478 16028 8484 16040
rect 8159 16000 8484 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 16028 14887 16031
rect 14918 16028 14924 16040
rect 14875 16000 14924 16028
rect 14875 15997 14887 16000
rect 14829 15991 14887 15997
rect 14918 15988 14924 16000
rect 14976 16028 14982 16040
rect 16628 16031 16686 16037
rect 14976 16000 15976 16028
rect 14976 15988 14982 16000
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15960 3479 15963
rect 3510 15960 3516 15972
rect 3467 15932 3516 15960
rect 3467 15929 3479 15932
rect 3421 15923 3479 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 4614 15960 4620 15972
rect 4575 15932 4620 15960
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 4706 15920 4712 15972
rect 4764 15960 4770 15972
rect 5258 15960 5264 15972
rect 4764 15932 4809 15960
rect 5219 15932 5264 15960
rect 4764 15920 4770 15932
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 7146 15963 7204 15969
rect 7146 15929 7158 15963
rect 7192 15929 7204 15963
rect 7146 15923 7204 15929
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15929 8723 15963
rect 8665 15923 8723 15929
rect 106 15852 112 15904
rect 164 15892 170 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 164 15864 1593 15892
rect 164 15852 170 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 3694 15892 3700 15904
rect 3655 15864 3700 15892
rect 1581 15855 1639 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 5994 15892 6000 15904
rect 5675 15864 6000 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7006 15892 7012 15904
rect 6687 15864 7012 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7006 15852 7012 15864
rect 7064 15892 7070 15904
rect 7161 15892 7189 15923
rect 8386 15892 8392 15904
rect 7064 15864 7189 15892
rect 8347 15864 8392 15892
rect 7064 15852 7070 15864
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 8680 15892 8708 15923
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 10226 15960 10232 15972
rect 8812 15932 9536 15960
rect 10187 15932 10232 15960
rect 8812 15920 8818 15932
rect 9306 15892 9312 15904
rect 8680 15864 9312 15892
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 9508 15892 9536 15932
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15929 10379 15963
rect 10870 15960 10876 15972
rect 10831 15932 10876 15960
rect 10321 15923 10379 15929
rect 9766 15892 9772 15904
rect 9508 15864 9772 15892
rect 9766 15852 9772 15864
rect 9824 15892 9830 15904
rect 10336 15892 10364 15923
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 13354 15960 13360 15972
rect 13315 15932 13360 15960
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 14001 15963 14059 15969
rect 13504 15932 13549 15960
rect 13504 15920 13510 15932
rect 14001 15929 14013 15963
rect 14047 15960 14059 15963
rect 14734 15960 14740 15972
rect 14047 15932 14740 15960
rect 14047 15929 14059 15932
rect 14001 15923 14059 15929
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 15191 15963 15249 15969
rect 15191 15929 15203 15963
rect 15237 15960 15249 15963
rect 15286 15960 15292 15972
rect 15237 15932 15292 15960
rect 15237 15929 15249 15932
rect 15191 15923 15249 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 15948 15960 15976 16000
rect 16628 15997 16640 16031
rect 16674 16028 16686 16031
rect 16868 16028 16896 16136
rect 17954 16124 17960 16136
rect 18012 16124 18018 16176
rect 20806 16164 20812 16176
rect 20767 16136 20812 16164
rect 20806 16124 20812 16136
rect 20864 16124 20870 16176
rect 21082 16124 21088 16176
rect 21140 16164 21146 16176
rect 22465 16167 22523 16173
rect 22465 16164 22477 16167
rect 21140 16136 22477 16164
rect 21140 16124 21146 16136
rect 22465 16133 22477 16136
rect 22511 16133 22523 16167
rect 22465 16127 22523 16133
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 19613 16099 19671 16105
rect 17920 16068 18552 16096
rect 17920 16056 17926 16068
rect 16674 16000 16896 16028
rect 17773 16031 17831 16037
rect 16674 15997 16686 16000
rect 16628 15991 16686 15997
rect 17773 15997 17785 16031
rect 17819 16028 17831 16031
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17819 16000 18337 16028
rect 17819 15997 17831 16000
rect 17773 15991 17831 15997
rect 18325 15997 18337 16000
rect 18371 16028 18383 16031
rect 18414 16028 18420 16040
rect 18371 16000 18420 16028
rect 18371 15997 18383 16000
rect 18325 15991 18383 15997
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18524 16037 18552 16068
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 19978 16096 19984 16108
rect 19659 16068 19984 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 21910 16096 21916 16108
rect 21499 16068 21916 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 22480 16096 22508 16127
rect 22554 16124 22560 16176
rect 22612 16164 22618 16176
rect 22833 16167 22891 16173
rect 22833 16164 22845 16167
rect 22612 16136 22845 16164
rect 22612 16124 22618 16136
rect 22833 16133 22845 16136
rect 22879 16133 22891 16167
rect 22833 16127 22891 16133
rect 24210 16124 24216 16176
rect 24268 16164 24274 16176
rect 24489 16167 24547 16173
rect 24489 16164 24501 16167
rect 24268 16136 24501 16164
rect 24268 16124 24274 16136
rect 24489 16133 24501 16136
rect 24535 16133 24547 16167
rect 24489 16127 24547 16133
rect 22646 16096 22652 16108
rect 22480 16068 22652 16096
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 22922 16056 22928 16108
rect 22980 16096 22986 16108
rect 23106 16096 23112 16108
rect 22980 16068 23112 16096
rect 22980 16056 22986 16068
rect 23106 16056 23112 16068
rect 23164 16096 23170 16108
rect 23164 16068 24751 16096
rect 23164 16056 23170 16068
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 24723 16037 24751 16068
rect 23712 16031 23770 16037
rect 23712 16028 23724 16031
rect 22888 16000 23724 16028
rect 22888 15988 22894 16000
rect 23712 15997 23724 16000
rect 23758 16028 23770 16031
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 23758 16000 24133 16028
rect 23758 15997 23770 16000
rect 23712 15991 23770 15997
rect 24121 15997 24133 16000
rect 24167 15997 24179 16031
rect 24121 15991 24179 15997
rect 24708 16031 24766 16037
rect 24708 15997 24720 16031
rect 24754 16028 24766 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24754 16000 25145 16028
rect 24754 15997 24766 16000
rect 24708 15991 24766 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 19934 15963 19992 15969
rect 19934 15960 19946 15963
rect 15948 15932 18092 15960
rect 11149 15895 11207 15901
rect 11149 15892 11161 15895
rect 9824 15864 11161 15892
rect 9824 15852 9830 15864
rect 11149 15861 11161 15864
rect 11195 15861 11207 15895
rect 15746 15892 15752 15904
rect 15707 15864 15752 15892
rect 11149 15855 11207 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 18064 15892 18092 15932
rect 19536 15932 19946 15960
rect 19536 15904 19564 15932
rect 19934 15929 19946 15932
rect 19980 15929 19992 15963
rect 19934 15923 19992 15929
rect 21545 15963 21603 15969
rect 21545 15929 21557 15963
rect 21591 15929 21603 15963
rect 22094 15960 22100 15972
rect 22055 15932 22100 15960
rect 21545 15923 21603 15929
rect 18141 15895 18199 15901
rect 18141 15892 18153 15895
rect 18064 15864 18153 15892
rect 18141 15861 18153 15864
rect 18187 15861 18199 15895
rect 18141 15855 18199 15861
rect 19153 15895 19211 15901
rect 19153 15861 19165 15895
rect 19199 15892 19211 15895
rect 19242 15892 19248 15904
rect 19199 15864 19248 15892
rect 19199 15861 19211 15864
rect 19153 15855 19211 15861
rect 19242 15852 19248 15864
rect 19300 15892 19306 15904
rect 19518 15892 19524 15904
rect 19300 15864 19524 15892
rect 19300 15852 19306 15864
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 21266 15892 21272 15904
rect 21179 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15892 21330 15904
rect 21560 15892 21588 15923
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 22554 15920 22560 15972
rect 22612 15960 22618 15972
rect 23799 15963 23857 15969
rect 23799 15960 23811 15963
rect 22612 15932 23811 15960
rect 22612 15920 22618 15932
rect 23799 15929 23811 15932
rect 23845 15929 23857 15963
rect 23799 15923 23857 15929
rect 22186 15892 22192 15904
rect 21324 15864 22192 15892
rect 21324 15852 21330 15864
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 22646 15892 22652 15904
rect 22428 15864 22652 15892
rect 22428 15852 22434 15864
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 7064 15660 7113 15688
rect 7064 15648 7070 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 12802 15688 12808 15700
rect 7699 15660 9904 15688
rect 12763 15660 12808 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 9876 15632 9904 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 13446 15688 13452 15700
rect 13403 15660 13452 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 13722 15688 13728 15700
rect 13683 15660 13728 15688
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 14323 15691 14381 15697
rect 14323 15688 14335 15691
rect 14056 15660 14335 15688
rect 14056 15648 14062 15660
rect 14323 15657 14335 15660
rect 14369 15657 14381 15691
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14323 15651 14381 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 15442 15660 17233 15688
rect 3142 15620 3148 15632
rect 3103 15592 3148 15620
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 7926 15620 7932 15632
rect 7887 15592 7932 15620
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 9490 15620 9496 15632
rect 9451 15592 9496 15620
rect 9490 15580 9496 15592
rect 9548 15580 9554 15632
rect 9858 15620 9864 15632
rect 9771 15592 9864 15620
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 15442 15620 15470 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 19613 15691 19671 15697
rect 19613 15657 19625 15691
rect 19659 15688 19671 15691
rect 21266 15688 21272 15700
rect 19659 15660 21272 15688
rect 19659 15657 19671 15660
rect 19613 15651 19671 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 22002 15688 22008 15700
rect 21963 15660 22008 15688
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22244 15660 22692 15688
rect 22244 15648 22250 15660
rect 15746 15620 15752 15632
rect 13786 15592 15470 15620
rect 15707 15592 15752 15620
rect 1464 15555 1522 15561
rect 1464 15521 1476 15555
rect 1510 15552 1522 15555
rect 2222 15552 2228 15564
rect 1510 15524 2228 15552
rect 1510 15521 1522 15524
rect 1464 15515 1522 15521
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15552 2467 15555
rect 3694 15552 3700 15564
rect 2455 15524 3700 15552
rect 2455 15521 2467 15524
rect 2409 15515 2467 15521
rect 3694 15512 3700 15524
rect 3752 15512 3758 15564
rect 4062 15552 4068 15564
rect 4023 15524 4068 15552
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 5074 15512 5080 15564
rect 5132 15552 5138 15564
rect 5169 15555 5227 15561
rect 5169 15552 5181 15555
rect 5132 15524 5181 15552
rect 5132 15512 5138 15524
rect 5169 15521 5181 15524
rect 5215 15521 5227 15555
rect 5169 15515 5227 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 5994 15552 6000 15564
rect 5767 15524 6000 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5994 15512 6000 15524
rect 6052 15552 6058 15564
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 6052 15524 6285 15552
rect 6052 15512 6058 15524
rect 6273 15521 6285 15524
rect 6319 15552 6331 15555
rect 6641 15555 6699 15561
rect 6641 15552 6653 15555
rect 6319 15524 6653 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 6641 15521 6653 15524
rect 6687 15552 6699 15555
rect 8386 15552 8392 15564
rect 6687 15524 8392 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8608 15555 8666 15561
rect 8608 15552 8620 15555
rect 8536 15524 8620 15552
rect 8536 15512 8542 15524
rect 8608 15521 8620 15524
rect 8654 15521 8666 15555
rect 8608 15515 8666 15521
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11204 15524 11253 15552
rect 11204 15512 11210 15524
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12437 15555 12495 15561
rect 12437 15552 12449 15555
rect 12308 15524 12449 15552
rect 12308 15512 12314 15524
rect 12437 15521 12449 15524
rect 12483 15552 12495 15555
rect 13786 15552 13814 15592
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 19055 15623 19113 15629
rect 19055 15589 19067 15623
rect 19101 15620 19113 15623
rect 19518 15620 19524 15632
rect 19101 15592 19524 15620
rect 19101 15589 19113 15592
rect 19055 15583 19113 15589
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 20717 15623 20775 15629
rect 20717 15589 20729 15623
rect 20763 15620 20775 15623
rect 20990 15620 20996 15632
rect 20763 15592 20996 15620
rect 20763 15589 20775 15592
rect 20717 15583 20775 15589
rect 20990 15580 20996 15592
rect 21048 15580 21054 15632
rect 21082 15580 21088 15632
rect 21140 15620 21146 15632
rect 22554 15620 22560 15632
rect 21140 15592 21185 15620
rect 22515 15592 22560 15620
rect 21140 15580 21146 15592
rect 22554 15580 22560 15592
rect 22612 15580 22618 15632
rect 22664 15629 22692 15660
rect 23014 15648 23020 15700
rect 23072 15688 23078 15700
rect 24118 15688 24124 15700
rect 23072 15660 24124 15688
rect 23072 15648 23078 15660
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 22649 15623 22707 15629
rect 22649 15589 22661 15623
rect 22695 15620 22707 15623
rect 23198 15620 23204 15632
rect 22695 15592 23204 15620
rect 22695 15589 22707 15592
rect 22649 15583 22707 15589
rect 23198 15580 23204 15592
rect 23256 15580 23262 15632
rect 12483 15524 13814 15552
rect 14252 15555 14310 15561
rect 12483 15521 12495 15524
rect 12437 15515 12495 15521
rect 14252 15521 14264 15555
rect 14298 15552 14310 15555
rect 14366 15552 14372 15564
rect 14298 15524 14372 15552
rect 14298 15521 14310 15524
rect 14252 15515 14310 15521
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15552 17739 15555
rect 17862 15552 17868 15564
rect 17727 15524 17868 15552
rect 17727 15521 17739 15524
rect 17681 15515 17739 15521
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15484 2007 15487
rect 2777 15487 2835 15493
rect 2777 15484 2789 15487
rect 1995 15456 2789 15484
rect 1995 15453 2007 15456
rect 1949 15447 2007 15453
rect 2777 15453 2789 15456
rect 2823 15484 2835 15487
rect 2866 15484 2872 15496
rect 2823 15456 2872 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 4614 15484 4620 15496
rect 3016 15456 4620 15484
rect 3016 15444 3022 15456
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15484 5963 15487
rect 6733 15487 6791 15493
rect 6733 15484 6745 15487
rect 5951 15456 6745 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 6733 15453 6745 15456
rect 6779 15484 6791 15487
rect 8110 15484 8116 15496
rect 6779 15456 8116 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15453 9827 15487
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 9769 15447 9827 15453
rect 1535 15419 1593 15425
rect 1535 15385 1547 15419
rect 1581 15416 1593 15419
rect 9490 15416 9496 15428
rect 1581 15388 9496 15416
rect 1581 15385 1593 15388
rect 1535 15379 1593 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 9784 15416 9812 15447
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 15654 15484 15660 15496
rect 15615 15456 15660 15484
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 17236 15484 17264 15515
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 18138 15484 18144 15496
rect 17236 15456 18144 15484
rect 10870 15416 10876 15428
rect 9784 15388 10876 15416
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 16206 15416 16212 15428
rect 16167 15388 16212 15416
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 2314 15348 2320 15360
rect 2275 15320 2320 15348
rect 2314 15308 2320 15320
rect 2372 15348 2378 15360
rect 2547 15351 2605 15357
rect 2547 15348 2559 15351
rect 2372 15320 2559 15348
rect 2372 15308 2378 15320
rect 2547 15317 2559 15320
rect 2593 15317 2605 15351
rect 2682 15348 2688 15360
rect 2643 15320 2688 15348
rect 2547 15311 2605 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 3418 15348 3424 15360
rect 3379 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4246 15348 4252 15360
rect 3927 15320 4252 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5074 15348 5080 15360
rect 5035 15320 5080 15348
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 8294 15348 8300 15360
rect 8255 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 8711 15351 8769 15357
rect 8711 15317 8723 15351
rect 8757 15348 8769 15351
rect 8846 15348 8852 15360
rect 8757 15320 8852 15348
rect 8757 15317 8769 15320
rect 8711 15311 8769 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10134 15348 10140 15360
rect 9456 15320 10140 15348
rect 9456 15308 9462 15320
rect 10134 15308 10140 15320
rect 10192 15348 10198 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 10192 15320 10701 15348
rect 10192 15308 10198 15320
rect 10689 15317 10701 15320
rect 10735 15317 10747 15351
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 10689 15311 10747 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11238 15308 11244 15360
rect 11296 15348 11302 15360
rect 11379 15351 11437 15357
rect 11379 15348 11391 15351
rect 11296 15320 11391 15348
rect 11296 15308 11302 15320
rect 11379 15317 11391 15320
rect 11425 15317 11437 15351
rect 11379 15311 11437 15317
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 17126 15348 17132 15360
rect 12584 15320 17132 15348
rect 12584 15308 12590 15320
rect 17126 15308 17132 15320
rect 17184 15348 17190 15360
rect 17236 15348 17264 15456
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18690 15484 18696 15496
rect 18651 15456 18696 15484
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21818 15484 21824 15496
rect 21039 15456 21824 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 22738 15484 22744 15496
rect 22204 15456 22744 15484
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 19058 15416 19064 15428
rect 18012 15388 19064 15416
rect 18012 15376 18018 15388
rect 19058 15376 19064 15388
rect 19116 15376 19122 15428
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 21545 15419 21603 15425
rect 21545 15416 21557 15419
rect 20772 15388 21557 15416
rect 20772 15376 20778 15388
rect 21545 15385 21557 15388
rect 21591 15416 21603 15419
rect 22094 15416 22100 15428
rect 21591 15388 22100 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 18506 15348 18512 15360
rect 17184 15320 17264 15348
rect 18467 15320 18512 15348
rect 17184 15308 17190 15320
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 20898 15308 20904 15360
rect 20956 15348 20962 15360
rect 22204 15348 22232 15456
rect 22738 15444 22744 15456
rect 22796 15484 22802 15496
rect 22833 15487 22891 15493
rect 22833 15484 22845 15487
rect 22796 15456 22845 15484
rect 22796 15444 22802 15456
rect 22833 15453 22845 15456
rect 22879 15453 22891 15487
rect 22833 15447 22891 15453
rect 20956 15320 22232 15348
rect 20956 15308 20962 15320
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1673 15147 1731 15153
rect 1673 15113 1685 15147
rect 1719 15144 1731 15147
rect 1854 15144 1860 15156
rect 1719 15116 1860 15144
rect 1719 15113 1731 15116
rect 1673 15107 1731 15113
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 2774 15144 2780 15156
rect 2735 15116 2780 15144
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3605 15147 3663 15153
rect 3605 15113 3617 15147
rect 3651 15144 3663 15147
rect 3878 15144 3884 15156
rect 3651 15116 3884 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 8110 15144 8116 15156
rect 8071 15116 8116 15144
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9916 15116 10057 15144
rect 9916 15104 9922 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 12250 15144 12256 15156
rect 12211 15116 12256 15144
rect 10045 15107 10103 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 13078 15144 13084 15156
rect 13039 15116 13084 15144
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 14277 15147 14335 15153
rect 14277 15113 14289 15147
rect 14323 15144 14335 15147
rect 14366 15144 14372 15156
rect 14323 15116 14372 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 17126 15144 17132 15156
rect 17087 15116 17132 15144
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 17589 15147 17647 15153
rect 17589 15113 17601 15147
rect 17635 15144 17647 15147
rect 17862 15144 17868 15156
rect 17635 15116 17868 15144
rect 17635 15113 17647 15116
rect 17589 15107 17647 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18414 15144 18420 15156
rect 18371 15116 18420 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18414 15104 18420 15116
rect 18472 15144 18478 15156
rect 19334 15144 19340 15156
rect 18472 15116 19340 15144
rect 18472 15104 18478 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20717 15147 20775 15153
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 21082 15144 21088 15156
rect 20763 15116 21088 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 21818 15144 21824 15156
rect 21779 15116 21824 15144
rect 21818 15104 21824 15116
rect 21876 15144 21882 15156
rect 22511 15147 22569 15153
rect 22511 15144 22523 15147
rect 21876 15116 22523 15144
rect 21876 15104 21882 15116
rect 22511 15113 22523 15116
rect 22557 15113 22569 15147
rect 23198 15144 23204 15156
rect 23159 15116 23204 15144
rect 22511 15107 22569 15113
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 1872 15076 1900 15104
rect 2409 15079 2467 15085
rect 2409 15076 2421 15079
rect 1872 15048 2421 15076
rect 2409 15045 2421 15048
rect 2455 15076 2467 15079
rect 2682 15076 2688 15088
rect 2455 15048 2688 15076
rect 2455 15045 2467 15048
rect 2409 15039 2467 15045
rect 2682 15036 2688 15048
rect 2740 15036 2746 15088
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2792 15008 2820 15104
rect 3142 15085 3148 15088
rect 3126 15079 3148 15085
rect 3126 15045 3138 15079
rect 3126 15039 3148 15045
rect 3142 15036 3148 15039
rect 3200 15036 3206 15088
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 7837 15079 7895 15085
rect 3844 15048 4936 15076
rect 3844 15036 3850 15048
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 1811 14980 3341 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 3329 14977 3341 14980
rect 3375 15008 3387 15011
rect 3973 15011 4031 15017
rect 3973 15008 3985 15011
rect 3375 14980 3985 15008
rect 3375 14977 3387 14980
rect 3329 14971 3387 14977
rect 3973 14977 3985 14980
rect 4019 15008 4031 15011
rect 4154 15008 4160 15020
rect 4019 14980 4160 15008
rect 4019 14977 4031 14980
rect 3973 14971 4031 14977
rect 4154 14968 4160 14980
rect 4212 14968 4218 15020
rect 1544 14943 1602 14949
rect 1544 14909 1556 14943
rect 1590 14940 1602 14943
rect 2314 14940 2320 14952
rect 1590 14912 2320 14940
rect 1590 14909 1602 14912
rect 1544 14903 1602 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 3191 14943 3249 14949
rect 3191 14940 3203 14943
rect 2464 14912 3203 14940
rect 2464 14900 2470 14912
rect 3191 14909 3203 14912
rect 3237 14940 3249 14943
rect 3418 14940 3424 14952
rect 3237 14912 3424 14940
rect 3237 14909 3249 14912
rect 3191 14903 3249 14909
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 4908 14940 4936 15048
rect 7837 15045 7849 15079
rect 7883 15076 7895 15079
rect 10413 15079 10471 15085
rect 10413 15076 10425 15079
rect 7883 15048 10425 15076
rect 7883 15045 7895 15048
rect 7837 15039 7895 15045
rect 10413 15045 10425 15048
rect 10459 15076 10471 15079
rect 10778 15076 10784 15088
rect 10459 15048 10784 15076
rect 10459 15045 10471 15048
rect 10413 15039 10471 15045
rect 10778 15036 10784 15048
rect 10836 15036 10842 15088
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 16669 15079 16727 15085
rect 16669 15076 16681 15079
rect 15712 15048 16681 15076
rect 15712 15036 15718 15048
rect 16669 15045 16681 15048
rect 16715 15076 16727 15079
rect 21726 15076 21732 15088
rect 16715 15048 21732 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 21726 15036 21732 15048
rect 21784 15036 21790 15088
rect 22370 15076 22376 15088
rect 22204 15048 22376 15076
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6917 15011 6975 15017
rect 6917 15008 6929 15011
rect 5951 14980 6929 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6917 14977 6929 14980
rect 6963 15008 6975 15011
rect 8294 15008 8300 15020
rect 6963 14980 8300 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 10042 15008 10048 15020
rect 9815 14980 10048 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 10042 14968 10048 14980
rect 10100 15008 10106 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10100 14980 10977 15008
rect 10100 14968 10106 14980
rect 10965 14977 10977 14980
rect 11011 15008 11023 15011
rect 11146 15008 11152 15020
rect 11011 14980 11152 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11146 14968 11152 14980
rect 11204 15008 11210 15020
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 11204 14980 11621 15008
rect 11204 14968 11210 14980
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 12676 14980 13676 15008
rect 12676 14968 12682 14980
rect 5166 14940 5172 14952
rect 4908 14912 5172 14940
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5442 14900 5448 14952
rect 5500 14940 5506 14952
rect 5721 14943 5779 14949
rect 5721 14940 5733 14943
rect 5500 14912 5733 14940
rect 5500 14900 5506 14912
rect 5721 14909 5733 14912
rect 5767 14940 5779 14943
rect 5994 14940 6000 14952
rect 5767 14912 6000 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 7024 14912 7322 14940
rect 1397 14875 1455 14881
rect 1397 14841 1409 14875
rect 1443 14872 1455 14875
rect 2038 14872 2044 14884
rect 1443 14844 2044 14872
rect 1443 14841 1455 14844
rect 1397 14835 1455 14841
rect 2038 14832 2044 14844
rect 2096 14872 2102 14884
rect 2774 14872 2780 14884
rect 2096 14844 2780 14872
rect 2096 14832 2102 14844
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 2866 14832 2872 14884
rect 2924 14872 2930 14884
rect 2960 14875 3018 14881
rect 2960 14872 2972 14875
rect 2924 14844 2972 14872
rect 2924 14832 2930 14844
rect 2960 14841 2972 14844
rect 3006 14841 3018 14875
rect 2960 14835 3018 14841
rect 7024 14816 7052 14912
rect 7294 14881 7322 14912
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13648 14949 13676 14980
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 14792 14980 15945 15008
rect 14792 14968 14798 14980
rect 15933 14977 15945 14980
rect 15979 15008 15991 15011
rect 17586 15008 17592 15020
rect 15979 14980 17592 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 15008 19211 15011
rect 19886 15008 19892 15020
rect 19199 14980 19892 15008
rect 19199 14977 19211 14980
rect 19153 14971 19211 14977
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 15008 20407 15011
rect 20530 15008 20536 15020
rect 20395 14980 20536 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 20530 14968 20536 14980
rect 20588 15008 20594 15020
rect 21082 15008 21088 15020
rect 20588 14980 21088 15008
rect 20588 14968 20594 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 13173 14943 13231 14949
rect 13173 14940 13185 14943
rect 13136 14912 13185 14940
rect 13136 14900 13142 14912
rect 13173 14909 13185 14912
rect 13219 14909 13231 14943
rect 13173 14903 13231 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 18414 14940 18420 14952
rect 18375 14912 18420 14940
rect 13633 14903 13691 14909
rect 18414 14900 18420 14912
rect 18472 14900 18478 14952
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 18874 14940 18880 14952
rect 18564 14912 18880 14940
rect 18564 14900 18570 14912
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 22204 14940 22232 15048
rect 22370 15036 22376 15048
rect 22428 15076 22434 15088
rect 22833 15079 22891 15085
rect 22833 15076 22845 15079
rect 22428 15048 22845 15076
rect 22428 15036 22434 15048
rect 22833 15045 22845 15048
rect 22879 15045 22891 15079
rect 22833 15039 22891 15045
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 22554 15008 22560 15020
rect 22327 14980 22560 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 22204 14912 22385 14940
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 23696 14943 23754 14949
rect 23696 14940 23708 14943
rect 23624 14912 23708 14940
rect 23624 14900 23630 14912
rect 23696 14909 23708 14912
rect 23742 14940 23754 14943
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23742 14912 24133 14940
rect 23742 14909 23754 14912
rect 23696 14903 23754 14909
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 7279 14875 7337 14881
rect 7279 14841 7291 14875
rect 7325 14841 7337 14875
rect 9122 14872 9128 14884
rect 9083 14844 9128 14872
rect 7279 14835 7337 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 9214 14832 9220 14884
rect 9272 14872 9278 14884
rect 9272 14844 9317 14872
rect 9272 14832 9278 14844
rect 9950 14832 9956 14884
rect 10008 14872 10014 14884
rect 10689 14875 10747 14881
rect 10689 14872 10701 14875
rect 10008 14844 10701 14872
rect 10008 14832 10014 14844
rect 10689 14841 10701 14844
rect 10735 14841 10747 14875
rect 10689 14835 10747 14841
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 4246 14804 4252 14816
rect 3936 14776 4252 14804
rect 3936 14764 3942 14776
rect 4246 14764 4252 14776
rect 4304 14804 4310 14816
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4304 14776 4353 14804
rect 4304 14764 4310 14776
rect 4341 14773 4353 14776
rect 4387 14804 4399 14807
rect 4709 14807 4767 14813
rect 4709 14804 4721 14807
rect 4387 14776 4721 14804
rect 4387 14773 4399 14776
rect 4341 14767 4399 14773
rect 4709 14773 4721 14776
rect 4755 14773 4767 14807
rect 4709 14767 4767 14773
rect 6273 14807 6331 14813
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6319 14776 6561 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7006 14804 7012 14816
rect 6595 14776 7012 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 8536 14776 8585 14804
rect 8536 14764 8542 14776
rect 8573 14773 8585 14776
rect 8619 14773 8631 14807
rect 10704 14804 10732 14835
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 10836 14844 10881 14872
rect 10836 14832 10842 14844
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 14366 14872 14372 14884
rect 12584 14844 14372 14872
rect 12584 14832 12590 14844
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 14737 14875 14795 14881
rect 14737 14841 14749 14875
rect 14783 14872 14795 14875
rect 15654 14872 15660 14884
rect 14783 14844 15660 14872
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 15654 14832 15660 14844
rect 15712 14832 15718 14884
rect 15746 14832 15752 14884
rect 15804 14872 15810 14884
rect 15804 14844 15849 14872
rect 15804 14832 15810 14844
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 19797 14875 19855 14881
rect 19797 14872 19809 14875
rect 18748 14844 19809 14872
rect 18748 14832 18754 14844
rect 19797 14841 19809 14844
rect 19843 14841 19855 14875
rect 20898 14872 20904 14884
rect 20859 14844 20904 14872
rect 19797 14835 19855 14841
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 20993 14875 21051 14881
rect 20993 14841 21005 14875
rect 21039 14872 21051 14875
rect 21082 14872 21088 14884
rect 21039 14844 21088 14872
rect 21039 14841 21051 14844
rect 20993 14835 21051 14841
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 21545 14875 21603 14881
rect 21545 14841 21557 14875
rect 21591 14872 21603 14875
rect 21634 14872 21640 14884
rect 21591 14844 21640 14872
rect 21591 14841 21603 14844
rect 21545 14835 21603 14841
rect 21634 14832 21640 14844
rect 21692 14832 21698 14884
rect 11054 14804 11060 14816
rect 10704 14776 11060 14804
rect 8573 14767 8631 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12713 14807 12771 14813
rect 12713 14773 12725 14807
rect 12759 14804 12771 14807
rect 12802 14804 12808 14816
rect 12759 14776 12808 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15473 14807 15531 14813
rect 15473 14804 15485 14807
rect 15151 14776 15485 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15473 14773 15485 14776
rect 15519 14804 15531 14807
rect 15764 14804 15792 14832
rect 19518 14804 19524 14816
rect 15519 14776 15792 14804
rect 19479 14776 19524 14804
rect 15519 14773 15531 14776
rect 15473 14767 15531 14773
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 21174 14764 21180 14816
rect 21232 14804 21238 14816
rect 23799 14807 23857 14813
rect 23799 14804 23811 14807
rect 21232 14776 23811 14804
rect 21232 14764 21238 14776
rect 23799 14773 23811 14776
rect 23845 14773 23857 14807
rect 23799 14767 23857 14773
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24581 14807 24639 14813
rect 24581 14804 24593 14807
rect 23992 14776 24593 14804
rect 23992 14764 23998 14776
rect 24581 14773 24593 14776
rect 24627 14804 24639 14807
rect 24670 14804 24676 14816
rect 24627 14776 24676 14804
rect 24627 14773 24639 14776
rect 24581 14767 24639 14773
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14600 2286 14612
rect 2590 14600 2596 14612
rect 2280 14572 2596 14600
rect 2280 14560 2286 14572
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 4982 14600 4988 14612
rect 3099 14572 4988 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5166 14600 5172 14612
rect 5127 14572 5172 14600
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 5920 14572 8938 14600
rect 1535 14535 1593 14541
rect 1535 14501 1547 14535
rect 1581 14532 1593 14535
rect 5920 14532 5948 14572
rect 1581 14504 5948 14532
rect 1581 14501 1593 14504
rect 1535 14495 1593 14501
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 7146 14535 7204 14541
rect 7146 14532 7158 14535
rect 7064 14504 7158 14532
rect 7064 14492 7070 14504
rect 7146 14501 7158 14504
rect 7192 14501 7204 14535
rect 8478 14532 8484 14544
rect 8439 14504 8484 14532
rect 7146 14495 7204 14501
rect 8478 14492 8484 14504
rect 8536 14492 8542 14544
rect 8910 14532 8938 14572
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9493 14603 9551 14609
rect 9493 14600 9505 14603
rect 9180 14572 9505 14600
rect 9180 14560 9186 14572
rect 9493 14569 9505 14572
rect 9539 14600 9551 14603
rect 10781 14603 10839 14609
rect 9539 14572 10456 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9398 14532 9404 14544
rect 8910 14504 9404 14532
rect 9398 14492 9404 14504
rect 9456 14492 9462 14544
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 10428 14541 10456 14572
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 10870 14600 10876 14612
rect 10827 14572 10876 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 16942 14600 16948 14612
rect 12032 14572 16804 14600
rect 16903 14572 16948 14600
rect 12032 14560 12038 14572
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9824 14504 9873 14532
rect 9824 14492 9830 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 9861 14495 9919 14501
rect 10413 14535 10471 14541
rect 10413 14501 10425 14535
rect 10459 14532 10471 14535
rect 10686 14532 10692 14544
rect 10459 14504 10692 14532
rect 10459 14501 10471 14504
rect 10413 14495 10471 14501
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 11790 14532 11796 14544
rect 11703 14504 11796 14532
rect 11790 14492 11796 14504
rect 11848 14532 11854 14544
rect 13811 14535 13869 14541
rect 11848 14504 12388 14532
rect 11848 14492 11854 14504
rect 1448 14467 1506 14473
rect 1448 14433 1460 14467
rect 1494 14464 1506 14467
rect 2130 14464 2136 14476
rect 1494 14436 2136 14464
rect 1494 14433 1506 14436
rect 1448 14427 1506 14433
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 2409 14467 2467 14473
rect 2409 14464 2421 14467
rect 2240 14436 2421 14464
rect 2240 14340 2268 14436
rect 2409 14433 2421 14436
rect 2455 14433 2467 14467
rect 3510 14464 3516 14476
rect 2409 14427 2467 14433
rect 2792 14436 3516 14464
rect 2792 14405 2820 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4614 14464 4620 14476
rect 4111 14436 4620 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 5442 14464 5448 14476
rect 4847 14436 5448 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5994 14464 6000 14476
rect 5675 14436 6000 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 8662 14473 8668 14476
rect 6825 14467 6883 14473
rect 6825 14464 6837 14467
rect 6696 14436 6837 14464
rect 6696 14424 6702 14436
rect 6825 14433 6837 14436
rect 6871 14464 6883 14467
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 6871 14436 8033 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8640 14467 8668 14473
rect 8640 14464 8652 14467
rect 8575 14436 8652 14464
rect 8021 14427 8079 14433
rect 8640 14433 8652 14436
rect 8720 14464 8726 14476
rect 9030 14464 9036 14476
rect 8720 14436 9036 14464
rect 8640 14427 8668 14433
rect 8662 14424 8668 14427
rect 8720 14424 8726 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 11974 14464 11980 14476
rect 11935 14436 11980 14464
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 12360 14473 12388 14504
rect 13811 14501 13823 14535
rect 13857 14532 13869 14535
rect 13906 14532 13912 14544
rect 13857 14504 13912 14532
rect 13857 14501 13869 14504
rect 13811 14495 13869 14501
rect 13906 14492 13912 14504
rect 13964 14492 13970 14544
rect 15470 14532 15476 14544
rect 15431 14504 15476 14532
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 16776 14532 16804 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 18690 14600 18696 14612
rect 18651 14572 18696 14600
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 20717 14603 20775 14609
rect 20717 14569 20729 14603
rect 20763 14600 20775 14603
rect 20898 14600 20904 14612
rect 20763 14572 20904 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 17494 14532 17500 14544
rect 16776 14504 17500 14532
rect 17494 14492 17500 14504
rect 17552 14532 17558 14544
rect 21082 14532 21088 14544
rect 17552 14504 18460 14532
rect 21043 14504 21088 14532
rect 17552 14492 17558 14504
rect 18432 14476 18460 14504
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 21634 14532 21640 14544
rect 21595 14504 21640 14532
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 21726 14492 21732 14544
rect 21784 14532 21790 14544
rect 23615 14535 23673 14541
rect 23615 14532 23627 14535
rect 21784 14504 23627 14532
rect 21784 14492 21790 14504
rect 23615 14501 23627 14504
rect 23661 14501 23673 14535
rect 23615 14495 23673 14501
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 12618 14464 12624 14476
rect 12391 14436 12624 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12618 14424 12624 14436
rect 12676 14464 12682 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 12676 14436 13185 14464
rect 12676 14424 12682 14436
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13446 14464 13452 14476
rect 13407 14436 13452 14464
rect 13173 14427 13231 14433
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14365 2835 14399
rect 2777 14359 2835 14365
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4212 14368 4445 14396
rect 4212 14356 4218 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 5408 14368 6285 14396
rect 5408 14356 5414 14368
rect 6273 14365 6285 14368
rect 6319 14396 6331 14399
rect 7190 14396 7196 14408
rect 6319 14368 7196 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 7190 14356 7196 14368
rect 7248 14396 7254 14408
rect 7650 14396 7656 14408
rect 7248 14368 7656 14396
rect 7248 14356 7254 14368
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 9548 14368 9781 14396
rect 9548 14356 9554 14368
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 12434 14396 12440 14408
rect 12395 14368 12440 14396
rect 9769 14359 9827 14365
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 13188 14396 13216 14427
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 17126 14464 17132 14476
rect 17087 14436 17132 14464
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 18414 14464 18420 14476
rect 18327 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18874 14464 18880 14476
rect 18835 14436 18880 14464
rect 18874 14424 18880 14436
rect 18932 14424 18938 14476
rect 22532 14467 22590 14473
rect 22532 14433 22544 14467
rect 22578 14464 22590 14467
rect 22738 14464 22744 14476
rect 22578 14436 22744 14464
rect 22578 14433 22590 14436
rect 22532 14427 22590 14433
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 23528 14467 23586 14473
rect 23528 14433 23540 14467
rect 23574 14464 23586 14467
rect 24118 14464 24124 14476
rect 23574 14436 24124 14464
rect 23574 14433 23586 14436
rect 23528 14427 23586 14433
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 13538 14396 13544 14408
rect 13188 14368 13544 14396
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 15378 14396 15384 14408
rect 15339 14368 15384 14396
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16758 14396 16764 14408
rect 16071 14368 16764 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20993 14399 21051 14405
rect 20993 14396 21005 14399
rect 20772 14368 21005 14396
rect 20772 14356 20778 14368
rect 20993 14365 21005 14368
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 2222 14288 2228 14340
rect 2280 14288 2286 14340
rect 2314 14288 2320 14340
rect 2372 14328 2378 14340
rect 2574 14331 2632 14337
rect 2574 14328 2586 14331
rect 2372 14300 2586 14328
rect 2372 14288 2378 14300
rect 2574 14297 2586 14300
rect 2620 14328 2632 14331
rect 3142 14328 3148 14340
rect 2620 14300 3148 14328
rect 2620 14297 2632 14300
rect 2574 14291 2632 14297
rect 3142 14288 3148 14300
rect 3200 14328 3206 14340
rect 4341 14331 4399 14337
rect 3200 14300 3924 14328
rect 3200 14288 3206 14300
rect 3896 14272 3924 14300
rect 4341 14297 4353 14331
rect 4387 14328 4399 14331
rect 4522 14328 4528 14340
rect 4387 14300 4528 14328
rect 4387 14297 4399 14300
rect 4341 14291 4399 14297
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 7745 14331 7803 14337
rect 7745 14297 7757 14331
rect 7791 14328 7803 14331
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 7791 14300 9045 14328
rect 7791 14297 7803 14300
rect 7745 14291 7803 14297
rect 9033 14297 9045 14300
rect 9079 14328 9091 14331
rect 9214 14328 9220 14340
rect 9079 14300 9220 14328
rect 9079 14297 9091 14300
rect 9033 14291 9091 14297
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 22603 14331 22661 14337
rect 22603 14328 22615 14331
rect 17736 14300 22615 14328
rect 17736 14288 17742 14300
rect 22603 14297 22615 14300
rect 22649 14297 22661 14331
rect 22603 14291 22661 14297
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4246 14269 4252 14272
rect 4230 14263 4252 14269
rect 4230 14229 4242 14263
rect 4230 14223 4252 14229
rect 4246 14220 4252 14223
rect 4304 14220 4310 14272
rect 6546 14260 6552 14272
rect 6507 14232 6552 14260
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 8711 14263 8769 14269
rect 8711 14229 8723 14263
rect 8757 14260 8769 14263
rect 8938 14260 8944 14272
rect 8757 14232 8944 14260
rect 8757 14229 8769 14232
rect 8711 14223 8769 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 19702 14260 19708 14272
rect 19663 14232 19708 14260
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 2682 14056 2688 14068
rect 2639 14028 2688 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 2004 13824 2145 13852
rect 2004 13812 2010 13824
rect 2133 13821 2145 13824
rect 2179 13852 2191 13855
rect 2608 13852 2636 14019
rect 2682 14016 2688 14028
rect 2740 14056 2746 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2740 14028 2881 14056
rect 2740 14016 2746 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 3218 14059 3276 14065
rect 3218 14025 3230 14059
rect 3264 14056 3276 14059
rect 3878 14056 3884 14068
rect 3264 14028 3884 14056
rect 3264 14025 3276 14028
rect 3218 14019 3276 14025
rect 2884 13988 2912 14019
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 6604 14028 7849 14056
rect 6604 14016 6610 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 8662 14056 8668 14068
rect 8623 14028 8668 14056
rect 7837 14019 7895 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9824 14028 10057 14056
rect 9824 14016 9830 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 11974 14056 11980 14068
rect 11935 14028 11980 14056
rect 10045 14019 10103 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 13817 14059 13875 14065
rect 13817 14025 13829 14059
rect 13863 14056 13875 14059
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 13863 14028 16405 14056
rect 13863 14025 13875 14028
rect 13817 14019 13875 14025
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 16393 14019 16451 14025
rect 16577 14059 16635 14065
rect 16577 14025 16589 14059
rect 16623 14056 16635 14059
rect 16942 14056 16948 14068
rect 16623 14028 16948 14056
rect 16623 14025 16635 14028
rect 16577 14019 16635 14025
rect 3329 13991 3387 13997
rect 3329 13988 3341 13991
rect 2884 13960 3341 13988
rect 3329 13957 3341 13960
rect 3375 13957 3387 13991
rect 5994 13988 6000 14000
rect 5907 13960 6000 13988
rect 3329 13951 3387 13957
rect 5994 13948 6000 13960
rect 6052 13988 6058 14000
rect 6730 13988 6736 14000
rect 6052 13960 6736 13988
rect 6052 13948 6058 13960
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 11992 13988 12020 14016
rect 7156 13960 12020 13988
rect 7156 13948 7162 13960
rect 12802 13948 12808 14000
rect 12860 13988 12866 14000
rect 13722 13988 13728 14000
rect 12860 13960 13728 13988
rect 12860 13948 12866 13960
rect 13722 13948 13728 13960
rect 13780 13988 13786 14000
rect 14093 13991 14151 13997
rect 14093 13988 14105 13991
rect 13780 13960 14105 13988
rect 13780 13948 13786 13960
rect 14093 13957 14105 13960
rect 14139 13957 14151 13991
rect 14093 13951 14151 13957
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 3602 13920 3608 13932
rect 3467 13892 3608 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 3602 13880 3608 13892
rect 3660 13920 3666 13932
rect 4154 13920 4160 13932
rect 3660 13892 4160 13920
rect 3660 13880 3666 13892
rect 4154 13880 4160 13892
rect 4212 13920 4218 13932
rect 4430 13920 4436 13932
rect 4212 13892 4436 13920
rect 4212 13880 4218 13892
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 5350 13920 5356 13932
rect 5184 13892 5356 13920
rect 5184 13861 5212 13892
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7926 13920 7932 13932
rect 7607 13892 7932 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8846 13880 8852 13932
rect 8904 13920 8910 13932
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 8904 13892 9137 13920
rect 8904 13880 8910 13892
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 9125 13883 9183 13889
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 12768 13892 14289 13920
rect 12768 13880 12774 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 16592 13920 16620 14019
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17460 14028 17785 14056
rect 17460 14016 17466 14028
rect 17773 14025 17785 14028
rect 17819 14056 17831 14059
rect 17862 14056 17868 14068
rect 17819 14028 17868 14056
rect 17819 14025 17831 14028
rect 17773 14019 17831 14025
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 18472 14028 19073 14056
rect 18472 14016 18478 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 20530 14056 20536 14068
rect 20491 14028 20536 14056
rect 19061 14019 19119 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 21140 14028 22385 14056
rect 21140 14016 21146 14028
rect 22373 14025 22385 14028
rect 22419 14025 22431 14059
rect 22373 14019 22431 14025
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 23937 14059 23995 14065
rect 23937 14056 23949 14059
rect 23900 14028 23949 14056
rect 23900 14016 23906 14028
rect 23937 14025 23949 14028
rect 23983 14025 23995 14059
rect 24946 14056 24952 14068
rect 24907 14028 24952 14056
rect 23937 14019 23995 14025
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13988 16911 13991
rect 17126 13988 17132 14000
rect 16899 13960 17132 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 24489 13991 24547 13997
rect 24489 13988 24501 13991
rect 19484 13960 24501 13988
rect 19484 13948 19490 13960
rect 17221 13923 17279 13929
rect 17221 13920 17233 13923
rect 15335 13892 16620 13920
rect 16776 13892 17233 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 2179 13824 2636 13852
rect 5169 13855 5227 13861
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 5169 13821 5181 13855
rect 5215 13821 5227 13855
rect 5442 13852 5448 13864
rect 5403 13824 5448 13852
rect 5169 13815 5227 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13852 7435 13855
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7423 13824 8217 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 8205 13821 8217 13824
rect 8251 13852 8263 13855
rect 8386 13852 8392 13864
rect 8251 13824 8392 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13596 13824 13829 13852
rect 13596 13812 13602 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 14047 13824 14105 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 14093 13821 14105 13824
rect 14139 13852 14151 13855
rect 15194 13852 15200 13864
rect 14139 13824 15200 13852
rect 14139 13821 14151 13824
rect 14093 13815 14151 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13852 16451 13855
rect 16776 13852 16804 13892
rect 17221 13889 17233 13892
rect 17267 13920 17279 13923
rect 17310 13920 17316 13932
rect 17267 13892 17316 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13920 19671 13923
rect 19702 13920 19708 13932
rect 19659 13892 19708 13920
rect 19659 13889 19671 13892
rect 19613 13883 19671 13889
rect 19702 13880 19708 13892
rect 19760 13920 19766 13932
rect 19760 13892 21312 13920
rect 19760 13880 19766 13892
rect 16439 13824 16804 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17920 13824 18061 13852
rect 17920 13812 17926 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18506 13812 18512 13864
rect 18564 13852 18570 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18564 13824 18613 13852
rect 18564 13812 18570 13824
rect 18601 13821 18613 13824
rect 18647 13852 18659 13855
rect 18874 13852 18880 13864
rect 18647 13824 18880 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 21174 13852 21180 13864
rect 21135 13824 21180 13852
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13784 2283 13787
rect 2406 13784 2412 13796
rect 2271 13756 2412 13784
rect 2271 13753 2283 13756
rect 2225 13747 2283 13753
rect 2406 13744 2412 13756
rect 2464 13744 2470 13796
rect 3050 13784 3056 13796
rect 3011 13756 3056 13784
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3786 13784 3792 13796
rect 3747 13756 3792 13784
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13784 5687 13787
rect 5994 13784 6000 13796
rect 5675 13756 6000 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 9214 13784 9220 13796
rect 9175 13756 9220 13784
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9769 13787 9827 13793
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 10686 13784 10692 13796
rect 9815 13756 10692 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 11333 13787 11391 13793
rect 10836 13756 10881 13784
rect 10836 13744 10842 13756
rect 11333 13753 11345 13787
rect 11379 13784 11391 13787
rect 11422 13784 11428 13796
rect 11379 13756 11428 13784
rect 11379 13753 11391 13756
rect 11333 13747 11391 13753
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13034 13787 13092 13793
rect 13034 13784 13046 13787
rect 12860 13756 13046 13784
rect 12860 13744 12866 13756
rect 13034 13753 13046 13756
rect 13080 13753 13092 13787
rect 14829 13787 14887 13793
rect 14829 13784 14841 13787
rect 13034 13747 13092 13753
rect 13648 13756 14841 13784
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3510 13716 3516 13728
rect 2832 13688 3516 13716
rect 2832 13676 2838 13688
rect 3510 13676 3516 13688
rect 3568 13676 3574 13728
rect 4522 13716 4528 13728
rect 4483 13688 4528 13716
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6236 13688 6561 13716
rect 6236 13676 6242 13688
rect 6549 13685 6561 13688
rect 6595 13716 6607 13719
rect 7006 13716 7012 13728
rect 6595 13688 7012 13716
rect 6595 13685 6607 13688
rect 6549 13679 6607 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8294 13716 8300 13728
rect 7892 13688 8300 13716
rect 7892 13676 7898 13688
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10796 13716 10824 13744
rect 10551 13688 10824 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 13648 13725 13676 13756
rect 14829 13753 14841 13756
rect 14875 13784 14887 13787
rect 15470 13784 15476 13796
rect 14875 13756 15476 13784
rect 14875 13753 14887 13756
rect 14829 13747 14887 13753
rect 15470 13744 15476 13756
rect 15528 13744 15534 13796
rect 15651 13787 15709 13793
rect 15651 13784 15663 13787
rect 15580 13756 15663 13784
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13412 13688 13645 13716
rect 13412 13676 13418 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15580 13716 15608 13756
rect 15651 13753 15663 13756
rect 15697 13784 15709 13787
rect 16022 13784 16028 13796
rect 15697 13756 16028 13784
rect 15697 13753 15709 13756
rect 15651 13747 15709 13753
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 19518 13784 19524 13796
rect 19431 13756 19524 13784
rect 16206 13716 16212 13728
rect 15252 13688 15608 13716
rect 16167 13688 16212 13716
rect 15252 13676 15258 13688
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 18322 13716 18328 13728
rect 18283 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 19444 13725 19472 13756
rect 19518 13744 19524 13756
rect 19576 13784 19582 13796
rect 19934 13787 19992 13793
rect 19934 13784 19946 13787
rect 19576 13756 19946 13784
rect 19576 13744 19582 13756
rect 19934 13753 19946 13756
rect 19980 13753 19992 13787
rect 19934 13747 19992 13753
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 19208 13688 19441 13716
rect 19208 13676 19214 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20588 13688 20821 13716
rect 20588 13676 20594 13688
rect 20809 13685 20821 13688
rect 20855 13716 20867 13719
rect 21174 13716 21180 13728
rect 20855 13688 21180 13716
rect 20855 13685 20867 13688
rect 20809 13679 20867 13685
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 21284 13716 21312 13892
rect 21450 13852 21456 13864
rect 21411 13824 21456 13852
rect 21450 13812 21456 13824
rect 21508 13812 21514 13864
rect 21910 13852 21916 13864
rect 21823 13824 21916 13852
rect 21910 13812 21916 13824
rect 21968 13852 21974 13864
rect 23014 13852 23020 13864
rect 21968 13824 23020 13852
rect 21968 13812 21974 13824
rect 23014 13812 23020 13824
rect 23072 13812 23078 13864
rect 23711 13861 23739 13960
rect 24489 13957 24501 13960
rect 24535 13957 24547 13991
rect 24489 13951 24547 13957
rect 25133 13923 25191 13929
rect 25133 13920 25145 13923
rect 24723 13892 25145 13920
rect 24723 13864 24751 13892
rect 25133 13889 25145 13892
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 23696 13855 23754 13861
rect 23696 13821 23708 13855
rect 23742 13821 23754 13855
rect 24670 13852 24676 13864
rect 24728 13861 24751 13864
rect 24728 13855 24766 13861
rect 24618 13824 24676 13852
rect 23696 13815 23754 13821
rect 24670 13812 24676 13824
rect 24754 13821 24766 13855
rect 24728 13815 24766 13821
rect 24728 13812 24734 13815
rect 22738 13784 22744 13796
rect 22699 13756 22744 13784
rect 22738 13744 22744 13756
rect 22796 13744 22802 13796
rect 21453 13719 21511 13725
rect 21453 13716 21465 13719
rect 21284 13688 21465 13716
rect 21453 13685 21465 13688
rect 21499 13685 21511 13719
rect 24118 13716 24124 13728
rect 24079 13688 24124 13716
rect 21453 13679 21511 13685
rect 24118 13676 24124 13688
rect 24176 13676 24182 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1535 13515 1593 13521
rect 1535 13481 1547 13515
rect 1581 13512 1593 13515
rect 1670 13512 1676 13524
rect 1581 13484 1676 13512
rect 1581 13481 1593 13484
rect 1535 13475 1593 13481
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 2188 13484 2237 13512
rect 2188 13472 2194 13484
rect 2225 13481 2237 13484
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3602 13512 3608 13524
rect 3559 13484 3608 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 9398 13512 9404 13524
rect 6595 13484 7604 13512
rect 9359 13484 9404 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 5258 13444 5264 13456
rect 1688 13416 5264 13444
rect 1464 13379 1522 13385
rect 1464 13345 1476 13379
rect 1510 13376 1522 13379
rect 1688 13376 1716 13416
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 5991 13447 6049 13453
rect 5991 13413 6003 13447
rect 6037 13444 6049 13447
rect 6178 13444 6184 13456
rect 6037 13416 6184 13444
rect 6037 13413 6049 13416
rect 5991 13407 6049 13413
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 7576 13453 7604 13484
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 10689 13515 10747 13521
rect 9968 13484 10640 13512
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 7742 13444 7748 13456
rect 7607 13416 7748 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 7742 13404 7748 13416
rect 7800 13444 7806 13456
rect 9968 13444 9996 13484
rect 7800 13416 9996 13444
rect 10090 13447 10148 13453
rect 7800 13404 7806 13416
rect 10090 13413 10102 13447
rect 10136 13413 10148 13447
rect 10612 13444 10640 13484
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 10778 13512 10784 13524
rect 10735 13484 10784 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 12802 13512 12808 13524
rect 12763 13484 12808 13512
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 13504 13484 14197 13512
rect 13504 13472 13510 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 15286 13512 15292 13524
rect 15151 13484 15292 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 20806 13472 20812 13524
rect 20864 13512 20870 13524
rect 22557 13515 22615 13521
rect 22557 13512 22569 13515
rect 20864 13484 22569 13512
rect 20864 13472 20870 13484
rect 22557 13481 22569 13484
rect 22603 13481 22615 13515
rect 24762 13512 24768 13524
rect 24723 13484 24768 13512
rect 22557 13475 22615 13481
rect 24762 13472 24768 13484
rect 24820 13472 24826 13524
rect 11238 13444 11244 13456
rect 10612 13416 11244 13444
rect 10090 13407 10148 13413
rect 1510 13348 1716 13376
rect 1510 13345 1522 13348
rect 1464 13339 1522 13345
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2188 13348 2421 13376
rect 2188 13336 2194 13348
rect 2409 13345 2421 13348
rect 2455 13376 2467 13379
rect 3050 13376 3056 13388
rect 2455 13348 3056 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 3694 13376 3700 13388
rect 3384 13348 3700 13376
rect 3384 13336 3390 13348
rect 3694 13336 3700 13348
rect 3752 13376 3758 13388
rect 3973 13379 4031 13385
rect 3973 13376 3985 13379
rect 3752 13348 3985 13376
rect 3752 13336 3758 13348
rect 3973 13345 3985 13348
rect 4019 13345 4031 13379
rect 3973 13339 4031 13345
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 4212 13348 6837 13376
rect 4212 13336 4218 13348
rect 6825 13345 6837 13348
rect 6871 13376 6883 13379
rect 7098 13376 7104 13388
rect 6871 13348 7104 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 10105 13376 10133 13407
rect 11238 13404 11244 13416
rect 11296 13444 11302 13456
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 11296 13416 11713 13444
rect 11296 13404 11302 13416
rect 11701 13413 11713 13416
rect 11747 13413 11759 13447
rect 13354 13444 13360 13456
rect 13315 13416 13360 13444
rect 11701 13407 11759 13413
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 14366 13404 14372 13456
rect 14424 13444 14430 13456
rect 15378 13444 15384 13456
rect 14424 13416 15384 13444
rect 14424 13404 14430 13416
rect 15378 13404 15384 13416
rect 15436 13444 15442 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15436 13416 15485 13444
rect 15436 13404 15442 13416
rect 15473 13413 15485 13416
rect 15519 13413 15531 13447
rect 15473 13407 15531 13413
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16942 13444 16948 13456
rect 16264 13416 16948 13444
rect 16264 13404 16270 13416
rect 16942 13404 16948 13416
rect 17000 13444 17006 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 17000 13416 17049 13444
rect 17000 13404 17006 13416
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 17037 13407 17095 13413
rect 19150 13404 19156 13456
rect 19208 13444 19214 13456
rect 19382 13447 19440 13453
rect 19382 13444 19394 13447
rect 19208 13416 19394 13444
rect 19208 13404 19214 13416
rect 19382 13413 19394 13416
rect 19428 13413 19440 13447
rect 22738 13444 22744 13456
rect 19382 13407 19440 13413
rect 19673 13416 22744 13444
rect 9732 13348 10133 13376
rect 9732 13336 9738 13348
rect 10686 13336 10692 13388
rect 10744 13376 10750 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10744 13348 10977 13376
rect 10744 13336 10750 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13376 17647 13379
rect 19673 13376 19701 13416
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 20898 13376 20904 13388
rect 17635 13348 19701 13376
rect 20859 13348 20904 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13308 2835 13311
rect 3418 13308 3424 13320
rect 2823 13280 3424 13308
rect 2823 13277 2835 13280
rect 2777 13271 2835 13277
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 4430 13308 4436 13320
rect 4391 13280 4436 13308
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 5994 13308 6000 13320
rect 5675 13280 6000 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 8478 13308 8484 13320
rect 7515 13280 8484 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 2685 13243 2743 13249
rect 2685 13240 2697 13243
rect 2464 13212 2697 13240
rect 2464 13200 2470 13212
rect 2685 13209 2697 13212
rect 2731 13240 2743 13243
rect 4341 13243 4399 13249
rect 4341 13240 4353 13243
rect 2731 13212 4353 13240
rect 2731 13209 2743 13212
rect 2685 13203 2743 13209
rect 4341 13209 4353 13212
rect 4387 13240 4399 13243
rect 4522 13240 4528 13252
rect 4387 13212 4528 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 4614 13200 4620 13252
rect 4672 13240 4678 13252
rect 5077 13243 5135 13249
rect 5077 13240 5089 13243
rect 4672 13212 5089 13240
rect 4672 13200 4678 13212
rect 5077 13209 5089 13212
rect 5123 13209 5135 13243
rect 5077 13203 5135 13209
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 7484 13240 7512 13271
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 8018 13240 8024 13252
rect 5408 13212 7512 13240
rect 7979 13212 8024 13240
rect 5408 13200 5414 13212
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 10980 13240 11008 13339
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13277 11943 13311
rect 13262 13308 13268 13320
rect 13175 13280 13268 13308
rect 11885 13271 11943 13277
rect 11900 13240 11928 13271
rect 13262 13268 13268 13280
rect 13320 13308 13326 13320
rect 13630 13308 13636 13320
rect 13320 13280 13636 13308
rect 13320 13268 13326 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 14274 13308 14280 13320
rect 13955 13280 14280 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 14274 13268 14280 13280
rect 14332 13308 14338 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 14332 13280 15393 13308
rect 14332 13268 14338 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16816 13280 16957 13308
rect 16816 13268 16822 13280
rect 16945 13277 16957 13280
rect 16991 13308 17003 13311
rect 17034 13308 17040 13320
rect 16991 13280 17040 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 10980 13212 11928 13240
rect 15933 13243 15991 13249
rect 15933 13209 15945 13243
rect 15979 13240 15991 13243
rect 17126 13240 17132 13252
rect 15979 13212 17132 13240
rect 15979 13209 15991 13212
rect 15933 13203 15991 13209
rect 17126 13200 17132 13212
rect 17184 13240 17190 13252
rect 17604 13240 17632 13339
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21232 13348 21373 13376
rect 21232 13336 21238 13348
rect 21361 13345 21373 13348
rect 21407 13376 21419 13379
rect 21910 13376 21916 13388
rect 21407 13348 21916 13376
rect 21407 13345 21419 13348
rect 21361 13339 21419 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22186 13336 22192 13388
rect 22244 13376 22250 13388
rect 22465 13379 22523 13385
rect 22465 13376 22477 13379
rect 22244 13348 22477 13376
rect 22244 13336 22250 13348
rect 22465 13345 22477 13348
rect 22511 13376 22523 13379
rect 22646 13376 22652 13388
rect 22511 13348 22652 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 23014 13376 23020 13388
rect 22975 13348 23020 13376
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24268 13348 24593 13376
rect 24268 13336 24274 13348
rect 24581 13345 24593 13348
rect 24627 13376 24639 13379
rect 24670 13376 24676 13388
rect 24627 13348 24676 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13308 19027 13311
rect 19061 13311 19119 13317
rect 19061 13308 19073 13311
rect 19015 13280 19073 13308
rect 19015 13277 19027 13280
rect 18969 13271 19027 13277
rect 19061 13277 19073 13280
rect 19107 13308 19119 13311
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 19107 13280 21465 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 17184 13212 17632 13240
rect 19981 13243 20039 13249
rect 17184 13200 17190 13212
rect 19981 13209 19993 13243
rect 20027 13240 20039 13243
rect 21082 13240 21088 13252
rect 20027 13212 21088 13240
rect 20027 13209 20039 13212
rect 19981 13203 20039 13209
rect 21082 13200 21088 13212
rect 21140 13200 21146 13252
rect 21174 13200 21180 13252
rect 21232 13240 21238 13252
rect 22462 13240 22468 13252
rect 21232 13212 22468 13240
rect 21232 13200 21238 13212
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 2547 13175 2605 13181
rect 2547 13172 2559 13175
rect 2372 13144 2559 13172
rect 2372 13132 2378 13144
rect 2547 13141 2559 13144
rect 2593 13141 2605 13175
rect 2547 13135 2605 13141
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3510 13172 3516 13184
rect 3099 13144 3516 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 3786 13132 3792 13144
rect 3844 13172 3850 13184
rect 4203 13175 4261 13181
rect 4203 13172 4215 13175
rect 3844 13144 4215 13172
rect 3844 13132 3850 13144
rect 4203 13141 4215 13144
rect 4249 13141 4261 13175
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4203 13135 4261 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 5166 13172 5172 13184
rect 5040 13144 5172 13172
rect 5040 13132 5046 13144
rect 5166 13132 5172 13144
rect 5224 13172 5230 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 5224 13144 5457 13172
rect 5224 13132 5230 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 5445 13135 5503 13141
rect 7285 13175 7343 13181
rect 7285 13141 7297 13175
rect 7331 13172 7343 13175
rect 8110 13172 8116 13184
rect 7331 13144 8116 13172
rect 7331 13141 7343 13144
rect 7285 13135 7343 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9214 13172 9220 13184
rect 9171 13144 9220 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 17678 13132 17684 13184
rect 17736 13172 17742 13184
rect 18049 13175 18107 13181
rect 18049 13172 18061 13175
rect 17736 13144 18061 13172
rect 17736 13132 17742 13144
rect 18049 13141 18061 13144
rect 18095 13172 18107 13175
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 18095 13144 18429 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18417 13141 18429 13144
rect 18463 13172 18475 13175
rect 18506 13172 18512 13184
rect 18463 13144 18512 13172
rect 18463 13141 18475 13144
rect 18417 13135 18475 13141
rect 18506 13132 18512 13144
rect 18564 13172 18570 13184
rect 20530 13172 20536 13184
rect 18564 13144 20536 13172
rect 18564 13132 18570 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 21266 13132 21272 13184
rect 21324 13172 21330 13184
rect 21913 13175 21971 13181
rect 21913 13172 21925 13175
rect 21324 13144 21925 13172
rect 21324 13132 21330 13144
rect 21913 13141 21925 13144
rect 21959 13141 21971 13175
rect 21913 13135 21971 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 2740 12940 2881 12968
rect 2740 12928 2746 12940
rect 2869 12937 2881 12940
rect 2915 12968 2927 12971
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2915 12940 3341 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3329 12937 3341 12940
rect 3375 12937 3387 12971
rect 3329 12931 3387 12937
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4430 12968 4436 12980
rect 4203 12940 4436 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4580 12940 4625 12968
rect 4580 12928 4586 12940
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6273 12971 6331 12977
rect 6273 12968 6285 12971
rect 6236 12940 6285 12968
rect 6236 12928 6242 12940
rect 6273 12937 6285 12940
rect 6319 12968 6331 12971
rect 7098 12968 7104 12980
rect 6319 12940 7104 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7742 12968 7748 12980
rect 7703 12940 7748 12968
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 8996 12940 11069 12968
rect 8996 12928 9002 12940
rect 11057 12937 11069 12940
rect 11103 12968 11115 12971
rect 11606 12968 11612 12980
rect 11103 12940 11612 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 15197 12971 15255 12977
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15378 12968 15384 12980
rect 15243 12940 15384 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 15565 12971 15623 12977
rect 15565 12937 15577 12971
rect 15611 12968 15623 12971
rect 16022 12968 16028 12980
rect 15611 12940 16028 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 22189 12971 22247 12977
rect 22189 12937 22201 12971
rect 22235 12968 22247 12971
rect 22925 12971 22983 12977
rect 22925 12968 22937 12971
rect 22235 12940 22937 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 22925 12937 22937 12940
rect 22971 12968 22983 12971
rect 23014 12968 23020 12980
rect 22971 12940 23020 12968
rect 22971 12937 22983 12940
rect 22925 12931 22983 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 2314 12860 2320 12912
rect 2372 12900 2378 12912
rect 3191 12903 3249 12909
rect 3191 12900 3203 12903
rect 2372 12872 3203 12900
rect 2372 12860 2378 12872
rect 3191 12869 3203 12872
rect 3237 12900 3249 12903
rect 3786 12900 3792 12912
rect 3237 12872 3792 12900
rect 3237 12869 3249 12872
rect 3191 12863 3249 12869
rect 3786 12860 3792 12872
rect 3844 12900 3850 12912
rect 4614 12900 4620 12912
rect 3844 12872 4620 12900
rect 3844 12860 3850 12872
rect 4614 12860 4620 12872
rect 4672 12900 4678 12912
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4672 12872 4813 12900
rect 4672 12860 4678 12872
rect 4801 12869 4813 12872
rect 4847 12869 4859 12903
rect 6546 12900 6552 12912
rect 4801 12863 4859 12869
rect 5000 12872 6552 12900
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 5000 12832 5028 12872
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 10686 12900 10692 12912
rect 10647 12872 10692 12900
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 11238 12900 11244 12912
rect 10836 12872 11244 12900
rect 10836 12860 10842 12872
rect 11238 12860 11244 12872
rect 11296 12900 11302 12912
rect 11425 12903 11483 12909
rect 11425 12900 11437 12903
rect 11296 12872 11437 12900
rect 11296 12860 11302 12872
rect 11425 12869 11437 12872
rect 11471 12869 11483 12903
rect 11425 12863 11483 12869
rect 14292 12872 17908 12900
rect 3757 12804 5028 12832
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3757 12764 3785 12804
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 9030 12832 9036 12844
rect 5316 12804 9036 12832
rect 5316 12792 5322 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9766 12832 9772 12844
rect 9539 12804 9772 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9766 12792 9772 12804
rect 9824 12832 9830 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 9824 12804 13001 12832
rect 9824 12792 9830 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 14292 12832 14320 12872
rect 12989 12795 13047 12801
rect 14200 12804 14320 12832
rect 3200 12736 3785 12764
rect 3200 12724 3206 12736
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 5040 12736 5181 12764
rect 5040 12724 5046 12736
rect 5169 12733 5181 12736
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 5721 12767 5779 12773
rect 5721 12764 5733 12767
rect 5500 12736 5733 12764
rect 5500 12724 5506 12736
rect 5721 12733 5733 12736
rect 5767 12764 5779 12767
rect 6362 12764 6368 12776
rect 5767 12736 6368 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 6968 12767 7026 12773
rect 6968 12733 6980 12767
rect 7014 12764 7026 12767
rect 7466 12764 7472 12776
rect 7014 12736 7472 12764
rect 7014 12733 7026 12736
rect 6968 12727 7026 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 11422 12764 11428 12776
rect 10796 12736 11428 12764
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 3326 12696 3332 12708
rect 3099 12668 3332 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 3789 12699 3847 12705
rect 3789 12665 3801 12699
rect 3835 12696 3847 12699
rect 5460 12696 5488 12724
rect 3835 12668 5488 12696
rect 5905 12699 5963 12705
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 7055 12699 7113 12705
rect 5951 12668 6408 12696
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 1670 12628 1676 12640
rect 1631 12600 1676 12628
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 2222 12588 2228 12640
rect 2280 12628 2286 12640
rect 2409 12631 2467 12637
rect 2409 12628 2421 12631
rect 2280 12600 2421 12628
rect 2280 12588 2286 12600
rect 2409 12597 2421 12600
rect 2455 12597 2467 12631
rect 6380 12628 6408 12668
rect 7055 12665 7067 12699
rect 7101 12696 7113 12699
rect 7650 12696 7656 12708
rect 7101 12668 7656 12696
rect 7101 12665 7113 12668
rect 7055 12659 7113 12665
rect 7650 12656 7656 12668
rect 7708 12656 7714 12708
rect 8018 12696 8024 12708
rect 7979 12668 8024 12696
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 8113 12699 8171 12705
rect 8113 12665 8125 12699
rect 8159 12696 8171 12699
rect 8386 12696 8392 12708
rect 8159 12668 8392 12696
rect 8159 12665 8171 12668
rect 8113 12659 8171 12665
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12696 8723 12699
rect 10134 12696 10140 12708
rect 8711 12668 9996 12696
rect 10095 12668 10140 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 6914 12628 6920 12640
rect 6380 12600 6920 12628
rect 2409 12591 2467 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7466 12628 7472 12640
rect 7427 12600 7472 12628
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 9766 12628 9772 12640
rect 7616 12600 9772 12628
rect 7616 12588 7622 12600
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9968 12628 9996 12668
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 10594 12696 10600 12708
rect 10275 12668 10600 12696
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 10796 12628 10824 12736
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12216 12736 12449 12764
rect 12216 12724 12222 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12894 12764 12900 12776
rect 12855 12736 12900 12764
rect 12437 12727 12495 12733
rect 12452 12696 12480 12727
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 14200 12773 14228 12804
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 17034 12832 17040 12844
rect 15988 12804 17040 12832
rect 15988 12792 15994 12804
rect 17034 12792 17040 12804
rect 17092 12832 17098 12844
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 17092 12804 17233 12832
rect 17092 12792 17098 12804
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17880 12832 17908 12872
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 22462 12900 22468 12912
rect 18104 12872 22468 12900
rect 18104 12860 18110 12872
rect 22462 12860 22468 12872
rect 22520 12860 22526 12912
rect 18598 12832 18604 12844
rect 17880 12804 18604 12832
rect 17221 12795 17279 12801
rect 18598 12792 18604 12804
rect 18656 12832 18662 12844
rect 21358 12832 21364 12844
rect 18656 12804 21364 12832
rect 18656 12792 18662 12804
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 21542 12832 21548 12844
rect 21503 12804 21548 12832
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13004 12736 14013 12764
rect 13004 12696 13032 12736
rect 14001 12733 14013 12736
rect 14047 12764 14059 12767
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 14047 12736 14197 12764
rect 14047 12733 14059 12736
rect 14001 12727 14059 12733
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14185 12727 14243 12733
rect 14338 12736 14565 12764
rect 14338 12696 14366 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15654 12764 15660 12776
rect 14875 12736 15660 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 18084 12767 18142 12773
rect 18084 12764 18096 12767
rect 15993 12736 18096 12764
rect 12452 12668 13032 12696
rect 13786 12668 14366 12696
rect 9968 12600 10824 12628
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11020 12600 11897 12628
rect 11020 12588 11026 12600
rect 11885 12597 11897 12600
rect 11931 12628 11943 12631
rect 12894 12628 12900 12640
rect 11931 12600 12900 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 13541 12631 13599 12637
rect 13541 12628 13553 12631
rect 13504 12600 13553 12628
rect 13504 12588 13510 12600
rect 13541 12597 13553 12600
rect 13587 12628 13599 12631
rect 13786 12628 13814 12668
rect 14458 12656 14464 12708
rect 14516 12696 14522 12708
rect 15993 12696 16021 12736
rect 18084 12733 18096 12736
rect 18130 12764 18142 12767
rect 18506 12764 18512 12776
rect 18130 12736 18512 12764
rect 18130 12733 18142 12736
rect 18084 12727 18142 12733
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 20806 12764 20812 12776
rect 19383 12736 20812 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 14516 12668 16021 12696
rect 14516 12656 14522 12668
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 18187 12699 18245 12705
rect 18187 12696 18199 12699
rect 16448 12668 18199 12696
rect 16448 12656 16454 12668
rect 18187 12665 18199 12668
rect 18233 12665 18245 12699
rect 19658 12699 19716 12705
rect 19658 12696 19670 12699
rect 18187 12659 18245 12665
rect 19168 12668 19670 12696
rect 19168 12640 19196 12668
rect 19658 12665 19670 12668
rect 19704 12696 19716 12699
rect 20533 12699 20591 12705
rect 20533 12696 20545 12699
rect 19704 12668 20545 12696
rect 19704 12665 19716 12668
rect 19658 12659 19716 12665
rect 20533 12665 20545 12668
rect 20579 12665 20591 12699
rect 21174 12696 21180 12708
rect 21135 12668 21180 12696
rect 20533 12659 20591 12665
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 21266 12656 21272 12708
rect 21324 12696 21330 12708
rect 21324 12668 21369 12696
rect 21324 12656 21330 12668
rect 16022 12628 16028 12640
rect 13587 12600 13814 12628
rect 15983 12600 16028 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 16574 12628 16580 12640
rect 16535 12600 16580 12628
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 19150 12628 19156 12640
rect 19111 12600 19156 12628
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 20254 12628 20260 12640
rect 20215 12600 20260 12628
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21284 12628 21312 12656
rect 20772 12600 21312 12628
rect 20772 12588 20778 12600
rect 22186 12588 22192 12640
rect 22244 12628 22250 12640
rect 22465 12631 22523 12637
rect 22465 12628 22477 12631
rect 22244 12600 22477 12628
rect 22244 12588 22250 12600
rect 22465 12597 22477 12600
rect 22511 12597 22523 12631
rect 23658 12628 23664 12640
rect 23619 12600 23664 12628
rect 22465 12591 22523 12597
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 24210 12588 24216 12640
rect 24268 12628 24274 12640
rect 24581 12631 24639 12637
rect 24581 12628 24593 12631
rect 24268 12600 24593 12628
rect 24268 12588 24274 12600
rect 24581 12597 24593 12600
rect 24627 12597 24639 12631
rect 24581 12591 24639 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 4430 12424 4436 12436
rect 4126 12396 4436 12424
rect 1397 12359 1455 12365
rect 1397 12325 1409 12359
rect 1443 12356 1455 12359
rect 4126 12356 4154 12396
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 4614 12424 4620 12436
rect 4575 12396 4620 12424
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 8386 12424 8392 12436
rect 7883 12396 8392 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8536 12396 8581 12424
rect 8536 12384 8542 12396
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8904 12396 9045 12424
rect 8904 12384 8910 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 13630 12424 13636 12436
rect 13591 12396 13636 12424
rect 9033 12387 9091 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 15654 12424 15660 12436
rect 15615 12396 15660 12424
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19208 12396 19257 12424
rect 19208 12384 19214 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 20714 12424 20720 12436
rect 19843 12396 20720 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 21174 12384 21180 12436
rect 21232 12424 21238 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21232 12396 21925 12424
rect 21232 12384 21238 12396
rect 21913 12393 21925 12396
rect 21959 12424 21971 12427
rect 23658 12424 23664 12436
rect 21959 12396 23664 12424
rect 21959 12393 21971 12396
rect 21913 12387 21971 12393
rect 23658 12384 23664 12396
rect 23716 12384 23722 12436
rect 1443 12328 4154 12356
rect 4295 12359 4353 12365
rect 1443 12325 1455 12328
rect 1397 12319 1455 12325
rect 4295 12325 4307 12359
rect 4341 12356 4353 12359
rect 5350 12356 5356 12368
rect 4341 12328 5356 12356
rect 4341 12325 4353 12328
rect 4295 12319 4353 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5531 12359 5589 12365
rect 5531 12325 5543 12359
rect 5577 12356 5589 12359
rect 7098 12356 7104 12368
rect 5577 12328 7104 12356
rect 5577 12325 5589 12328
rect 5531 12319 5589 12325
rect 7098 12316 7104 12328
rect 7156 12356 7162 12368
rect 7238 12359 7296 12365
rect 7238 12356 7250 12359
rect 7156 12328 7250 12356
rect 7156 12316 7162 12328
rect 7238 12325 7250 12328
rect 7284 12356 7296 12359
rect 7558 12356 7564 12368
rect 7284 12328 7564 12356
rect 7284 12325 7296 12328
rect 7238 12319 7296 12325
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 9401 12359 9459 12365
rect 9401 12356 9413 12359
rect 7708 12328 9413 12356
rect 7708 12316 7714 12328
rect 9401 12325 9413 12328
rect 9447 12356 9459 12359
rect 10134 12356 10140 12368
rect 9447 12328 10140 12356
rect 9447 12325 9459 12328
rect 9401 12319 9459 12325
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 10870 12356 10876 12368
rect 10831 12328 10876 12356
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 11422 12356 11428 12368
rect 11383 12328 11428 12356
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 12437 12359 12495 12365
rect 12437 12356 12449 12359
rect 11848 12328 12449 12356
rect 11848 12316 11854 12328
rect 12437 12325 12449 12328
rect 12483 12325 12495 12359
rect 12437 12319 12495 12325
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 16574 12356 16580 12368
rect 16439 12328 16580 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 16945 12359 17003 12365
rect 16945 12325 16957 12359
rect 16991 12356 17003 12359
rect 17126 12356 17132 12368
rect 16991 12328 17132 12356
rect 16991 12325 17003 12328
rect 16945 12319 17003 12325
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 20254 12316 20260 12368
rect 20312 12356 20318 12368
rect 20622 12356 20628 12368
rect 20312 12328 20628 12356
rect 20312 12316 20318 12328
rect 20622 12316 20628 12328
rect 20680 12356 20686 12368
rect 21085 12359 21143 12365
rect 21085 12356 21097 12359
rect 20680 12328 21097 12356
rect 20680 12316 20686 12328
rect 21085 12325 21097 12328
rect 21131 12325 21143 12359
rect 21085 12319 21143 12325
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2096 12260 2421 12288
rect 2096 12248 2102 12260
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2409 12251 2467 12257
rect 4062 12248 4068 12300
rect 4120 12288 4126 12300
rect 4192 12291 4250 12297
rect 4192 12288 4204 12291
rect 4120 12260 4204 12288
rect 4120 12248 4126 12260
rect 4192 12257 4204 12260
rect 4238 12257 4250 12291
rect 4192 12251 4250 12257
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 6052 12260 8125 12288
rect 6052 12248 6058 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 9744 12291 9802 12297
rect 9744 12257 9756 12291
rect 9790 12288 9802 12291
rect 9858 12288 9864 12300
rect 9790 12260 9864 12288
rect 9790 12257 9802 12260
rect 9744 12251 9802 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 14252 12291 14310 12297
rect 14252 12257 14264 12291
rect 14298 12288 14310 12291
rect 14366 12288 14372 12300
rect 14298 12260 14372 12288
rect 14298 12257 14310 12260
rect 14252 12251 14310 12257
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 17770 12288 17776 12300
rect 17731 12260 17776 12288
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 20806 12288 20812 12300
rect 20211 12260 20812 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 22462 12288 22468 12300
rect 22520 12297 22526 12300
rect 22520 12291 22558 12297
rect 22410 12260 22468 12288
rect 22462 12248 22468 12260
rect 22546 12288 22558 12291
rect 23512 12291 23570 12297
rect 23512 12288 23524 12291
rect 22546 12260 23524 12288
rect 22546 12257 22558 12260
rect 22520 12251 22558 12257
rect 23512 12257 23524 12260
rect 23558 12257 23570 12291
rect 23512 12251 23570 12257
rect 22520 12248 22526 12251
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2240 12192 2789 12220
rect 2240 12096 2268 12192
rect 2777 12189 2789 12192
rect 2823 12220 2835 12223
rect 3418 12220 3424 12232
rect 2823 12192 3424 12220
rect 2823 12189 2835 12192
rect 2777 12183 2835 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4396 12192 5181 12220
rect 4396 12180 4402 12192
rect 5169 12189 5181 12192
rect 5215 12220 5227 12223
rect 6454 12220 6460 12232
rect 5215 12192 6460 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 6914 12220 6920 12232
rect 6875 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 12342 12220 12348 12232
rect 10827 12192 11468 12220
rect 12303 12192 12348 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 11440 12164 11468 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 13354 12220 13360 12232
rect 13267 12192 13360 12220
rect 12621 12183 12679 12189
rect 2406 12112 2412 12164
rect 2464 12152 2470 12164
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 2464 12124 2697 12152
rect 2464 12112 2470 12124
rect 2685 12121 2697 12124
rect 2731 12152 2743 12155
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 2731 12124 3801 12152
rect 2731 12121 2743 12124
rect 2685 12115 2743 12121
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 3789 12115 3847 12121
rect 4126 12124 4997 12152
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 2547 12087 2605 12093
rect 2547 12084 2559 12087
rect 2372 12056 2559 12084
rect 2372 12044 2378 12056
rect 2547 12053 2559 12056
rect 2593 12053 2605 12087
rect 2547 12047 2605 12053
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3053 12087 3111 12093
rect 3053 12084 3065 12087
rect 3016 12056 3065 12084
rect 3016 12044 3022 12056
rect 3053 12053 3065 12056
rect 3099 12053 3111 12087
rect 3053 12047 3111 12053
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 4126 12084 4154 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 7892 12124 10149 12152
rect 7892 12112 7898 12124
rect 10137 12121 10149 12124
rect 10183 12152 10195 12155
rect 10686 12152 10692 12164
rect 10183 12124 10692 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10686 12112 10692 12124
rect 10744 12112 10750 12164
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 12636 12152 12664 12183
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 16301 12223 16359 12229
rect 13412 12192 13814 12220
rect 13412 12180 13418 12192
rect 11480 12124 12664 12152
rect 13786 12152 13814 12192
rect 16301 12189 16313 12223
rect 16347 12220 16359 12223
rect 16666 12220 16672 12232
rect 16347 12192 16672 12220
rect 16347 12189 16359 12192
rect 16301 12183 16359 12189
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 18230 12220 18236 12232
rect 16776 12192 18236 12220
rect 16776 12152 16804 12192
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 20993 12223 21051 12229
rect 20993 12220 21005 12223
rect 20763 12192 21005 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 20993 12189 21005 12192
rect 21039 12220 21051 12223
rect 23615 12223 23673 12229
rect 23615 12220 23627 12223
rect 21039 12192 23627 12220
rect 21039 12189 21051 12192
rect 20993 12183 21051 12189
rect 23615 12189 23627 12192
rect 23661 12189 23673 12223
rect 23615 12183 23673 12189
rect 13786 12124 16804 12152
rect 18785 12155 18843 12161
rect 11480 12112 11486 12124
rect 18785 12121 18797 12155
rect 18831 12152 18843 12155
rect 18892 12152 18920 12183
rect 21266 12152 21272 12164
rect 18831 12124 21272 12152
rect 18831 12121 18843 12124
rect 18785 12115 18843 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 21542 12152 21548 12164
rect 21503 12124 21548 12152
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 6086 12084 6092 12096
rect 3384 12056 4154 12084
rect 6047 12056 6092 12084
rect 3384 12044 3390 12056
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6362 12044 6368 12096
rect 6420 12084 6426 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 6420 12056 6469 12084
rect 6420 12044 6426 12056
rect 6457 12053 6469 12056
rect 6503 12084 6515 12087
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6503 12056 6837 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 6825 12053 6837 12056
rect 6871 12084 6883 12087
rect 8110 12084 8116 12096
rect 6871 12056 8116 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 9815 12087 9873 12093
rect 9815 12053 9827 12087
rect 9861 12084 9873 12087
rect 9950 12084 9956 12096
rect 9861 12056 9956 12084
rect 9861 12053 9873 12056
rect 9815 12047 9873 12053
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10502 12084 10508 12096
rect 10463 12056 10508 12084
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 14323 12087 14381 12093
rect 14323 12053 14335 12087
rect 14369 12084 14381 12087
rect 15378 12084 15384 12096
rect 14369 12056 15384 12084
rect 14369 12053 14381 12056
rect 14323 12047 14381 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16022 12084 16028 12096
rect 15983 12056 16028 12084
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 17911 12087 17969 12093
rect 17911 12053 17923 12087
rect 17957 12084 17969 12087
rect 18966 12084 18972 12096
rect 17957 12056 18972 12084
rect 17957 12053 17969 12056
rect 17911 12047 17969 12053
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 22603 12087 22661 12093
rect 22603 12084 22615 12087
rect 19116 12056 22615 12084
rect 19116 12044 19122 12056
rect 22603 12053 22615 12056
rect 22649 12053 22661 12087
rect 22603 12047 22661 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1946 11880 1952 11892
rect 1907 11852 1952 11880
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 2096 11852 2329 11880
rect 2096 11840 2102 11852
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 4028 11852 4629 11880
rect 4028 11840 4034 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6362 11880 6368 11892
rect 6319 11852 6368 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 2222 11821 2228 11824
rect 2206 11815 2228 11821
rect 2206 11812 2218 11815
rect 2135 11784 2218 11812
rect 2206 11781 2218 11784
rect 2280 11812 2286 11824
rect 3053 11815 3111 11821
rect 3053 11812 3065 11815
rect 2280 11784 3065 11812
rect 2206 11775 2228 11781
rect 2222 11772 2228 11775
rect 2280 11772 2286 11784
rect 3053 11781 3065 11784
rect 3099 11781 3111 11815
rect 3053 11775 3111 11781
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2409 11747 2467 11753
rect 2409 11744 2421 11747
rect 2372 11716 2421 11744
rect 2372 11704 2378 11716
rect 2409 11713 2421 11716
rect 2455 11744 2467 11747
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 2455 11716 3433 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 3421 11713 3433 11716
rect 3467 11713 3479 11747
rect 4338 11744 4344 11756
rect 4299 11716 4344 11744
rect 3421 11707 3479 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 6288 11744 6316 11843
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 8389 11883 8447 11889
rect 8389 11880 8401 11883
rect 6972 11852 8401 11880
rect 6972 11840 6978 11852
rect 8389 11849 8401 11852
rect 8435 11849 8447 11883
rect 8389 11843 8447 11849
rect 9677 11883 9735 11889
rect 9677 11849 9689 11883
rect 9723 11880 9735 11883
rect 9858 11880 9864 11892
rect 9723 11852 9864 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 10870 11880 10876 11892
rect 10735 11852 10876 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10870 11840 10876 11852
rect 10928 11880 10934 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10928 11852 10977 11880
rect 10928 11840 10934 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 11422 11880 11428 11892
rect 11383 11852 11428 11880
rect 10965 11843 11023 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12434 11880 12440 11892
rect 12299 11852 12440 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12802 11880 12808 11892
rect 12763 11852 12808 11880
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 15470 11880 15476 11892
rect 13924 11852 15476 11880
rect 5092 11716 6316 11744
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 2004 11648 2053 11676
rect 2004 11636 2010 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 3786 11676 3792 11688
rect 3747 11648 3792 11676
rect 2041 11639 2099 11645
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 5092 11676 5120 11716
rect 4203 11648 5120 11676
rect 5445 11679 5503 11685
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5534 11676 5540 11688
rect 5491 11648 5540 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5736 11685 5764 11716
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 11790 11744 11796 11756
rect 10744 11716 11796 11744
rect 10744 11704 10750 11716
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 12452 11744 12480 11840
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 13924 11821 13952 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15841 11883 15899 11889
rect 15841 11849 15853 11883
rect 15887 11880 15899 11883
rect 16574 11880 16580 11892
rect 15887 11852 16580 11880
rect 15887 11849 15899 11852
rect 15841 11843 15899 11849
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 19392 11852 19441 11880
rect 19392 11840 19398 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 19429 11843 19487 11849
rect 13909 11815 13967 11821
rect 13909 11812 13921 11815
rect 13780 11784 13921 11812
rect 13780 11772 13786 11784
rect 13909 11781 13921 11784
rect 13955 11781 13967 11815
rect 13909 11775 13967 11781
rect 14642 11772 14648 11824
rect 14700 11812 14706 11824
rect 17405 11815 17463 11821
rect 17405 11812 17417 11815
rect 14700 11784 17417 11812
rect 14700 11772 14706 11784
rect 17405 11781 17417 11784
rect 17451 11812 17463 11815
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 17451 11784 17693 11812
rect 17451 11781 17463 11784
rect 17405 11775 17463 11781
rect 17681 11781 17693 11784
rect 17727 11781 17739 11815
rect 17681 11775 17739 11781
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12452 11716 13001 11744
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 15105 11747 15163 11753
rect 15105 11744 15117 11747
rect 14332 11716 15117 11744
rect 14332 11704 14338 11716
rect 15105 11713 15117 11716
rect 15151 11744 15163 11747
rect 16022 11744 16028 11756
rect 15151 11716 16028 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16390 11744 16396 11756
rect 16351 11716 16396 11744
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16666 11744 16672 11756
rect 16627 11716 16672 11744
rect 16666 11704 16672 11716
rect 16724 11744 16730 11756
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 16724 11716 18429 11744
rect 16724 11704 16730 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 5951 11648 6837 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 6825 11645 6837 11648
rect 6871 11676 6883 11679
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 6871 11648 8033 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 8021 11645 8033 11648
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 8824 11679 8882 11685
rect 8824 11645 8836 11679
rect 8870 11676 8882 11679
rect 8870 11648 8984 11676
rect 8870 11645 8882 11648
rect 8824 11639 8882 11645
rect 2774 11608 2780 11620
rect 2735 11580 2780 11608
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6362 11608 6368 11620
rect 6144 11580 6368 11608
rect 6144 11568 6150 11580
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 7098 11608 7104 11620
rect 6656 11580 7104 11608
rect 6656 11552 6684 11580
rect 7098 11568 7104 11580
rect 7156 11617 7162 11620
rect 7156 11611 7204 11617
rect 7156 11577 7158 11611
rect 7192 11577 7204 11611
rect 8956 11608 8984 11648
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9180 11648 9781 11676
rect 9180 11636 9186 11648
rect 9769 11645 9781 11648
rect 9815 11676 9827 11679
rect 10502 11676 10508 11688
rect 9815 11648 10508 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 19444 11676 19472 11843
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20625 11883 20683 11889
rect 20625 11880 20637 11883
rect 20588 11852 20637 11880
rect 20588 11840 20594 11852
rect 20625 11849 20637 11852
rect 20671 11849 20683 11883
rect 22462 11880 22468 11892
rect 22423 11852 22468 11880
rect 20625 11843 20683 11849
rect 20640 11744 20668 11843
rect 22462 11840 22468 11852
rect 22520 11880 22526 11892
rect 23753 11883 23811 11889
rect 23753 11880 23765 11883
rect 22520 11852 23765 11880
rect 22520 11840 22526 11852
rect 23753 11849 23765 11852
rect 23799 11849 23811 11883
rect 24762 11880 24768 11892
rect 24723 11852 24768 11880
rect 23753 11843 23811 11849
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 20640 11716 21680 11744
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19444 11648 19625 11676
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 20070 11676 20076 11688
rect 20031 11648 20076 11676
rect 19613 11639 19671 11645
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 21082 11676 21088 11688
rect 20864 11648 21088 11676
rect 20864 11636 20870 11648
rect 21082 11636 21088 11648
rect 21140 11676 21146 11688
rect 21652 11685 21680 11716
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 21140 11648 21189 11676
rect 21140 11636 21146 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 21637 11679 21695 11685
rect 21637 11645 21649 11679
rect 21683 11645 21695 11679
rect 24578 11676 24584 11688
rect 24539 11648 24584 11676
rect 21637 11639 21695 11645
rect 24578 11636 24584 11648
rect 24636 11676 24642 11688
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24636 11648 25145 11676
rect 24636 11636 24642 11648
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 9217 11611 9275 11617
rect 9217 11608 9229 11611
rect 8956 11580 9229 11608
rect 7156 11571 7204 11577
rect 9217 11577 9229 11580
rect 9263 11608 9275 11611
rect 9490 11608 9496 11620
rect 9263 11580 9496 11608
rect 9263 11577 9275 11580
rect 9217 11571 9275 11577
rect 7156 11568 7162 11571
rect 9490 11568 9496 11580
rect 9548 11568 9554 11620
rect 9858 11568 9864 11620
rect 9916 11608 9922 11620
rect 10131 11611 10189 11617
rect 10131 11608 10143 11611
rect 9916 11580 10143 11608
rect 9916 11568 9922 11580
rect 10131 11577 10143 11580
rect 10177 11608 10189 11611
rect 12802 11608 12808 11620
rect 10177 11580 12808 11608
rect 10177 11577 10189 11580
rect 10131 11571 10189 11577
rect 12802 11568 12808 11580
rect 12860 11608 12866 11620
rect 13354 11617 13360 11620
rect 13310 11611 13360 11617
rect 13310 11608 13322 11611
rect 12860 11580 13322 11608
rect 12860 11568 12866 11580
rect 13310 11577 13322 11580
rect 13356 11577 13360 11611
rect 13310 11571 13360 11577
rect 13354 11568 13360 11571
rect 13412 11568 13418 11620
rect 14277 11611 14335 11617
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 14366 11608 14372 11620
rect 14323 11580 14372 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14826 11617 14832 11620
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 14818 11611 14832 11617
rect 14818 11608 14830 11611
rect 14691 11580 14830 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 14818 11577 14830 11580
rect 14818 11571 14832 11577
rect 14826 11568 14832 11571
rect 14884 11568 14890 11620
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 16209 11611 16267 11617
rect 16209 11608 16221 11611
rect 14976 11580 16221 11608
rect 14976 11568 14982 11580
rect 16209 11577 16221 11580
rect 16255 11608 16267 11611
rect 16485 11611 16543 11617
rect 16485 11608 16497 11611
rect 16255 11580 16497 11608
rect 16255 11577 16267 11580
rect 16209 11571 16267 11577
rect 16485 11577 16497 11580
rect 16531 11577 16543 11611
rect 16485 11571 16543 11577
rect 17681 11611 17739 11617
rect 17681 11577 17693 11611
rect 17727 11608 17739 11611
rect 18141 11611 18199 11617
rect 18141 11608 18153 11611
rect 17727 11580 18153 11608
rect 17727 11577 17739 11580
rect 17681 11571 17739 11577
rect 18141 11577 18153 11580
rect 18187 11577 18199 11611
rect 18141 11571 18199 11577
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 18288 11580 18333 11608
rect 18288 11568 18294 11580
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 21542 11608 21548 11620
rect 19392 11580 21548 11608
rect 19392 11568 19398 11580
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 6638 11540 6644 11552
rect 5123 11512 6644 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 6638 11500 6644 11512
rect 6696 11500 6702 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 7834 11540 7840 11552
rect 7791 11512 7840 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8895 11543 8953 11549
rect 8895 11509 8907 11543
rect 8941 11540 8953 11543
rect 9030 11540 9036 11552
rect 8941 11512 9036 11540
rect 8941 11509 8953 11512
rect 8895 11503 8953 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 17770 11540 17776 11552
rect 17731 11512 17776 11540
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 19150 11540 19156 11552
rect 19111 11512 19156 11540
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19889 11543 19947 11549
rect 19889 11509 19901 11543
rect 19935 11540 19947 11543
rect 19978 11540 19984 11552
rect 19935 11512 19984 11540
rect 19935 11509 19947 11512
rect 19889 11503 19947 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 20864 11512 21005 11540
rect 20864 11500 20870 11512
rect 20993 11509 21005 11512
rect 21039 11509 21051 11543
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 20993 11503 21051 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 23753 11543 23811 11549
rect 23753 11509 23765 11543
rect 23799 11540 23811 11543
rect 23937 11543 23995 11549
rect 23937 11540 23949 11543
rect 23799 11512 23949 11540
rect 23799 11509 23811 11512
rect 23753 11503 23811 11509
rect 23937 11509 23949 11512
rect 23983 11540 23995 11543
rect 24670 11540 24676 11552
rect 23983 11512 24676 11540
rect 23983 11509 23995 11512
rect 23937 11503 23995 11509
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4396 11308 5273 11336
rect 4396 11296 4402 11308
rect 5261 11305 5273 11308
rect 5307 11336 5319 11339
rect 5534 11336 5540 11348
rect 5307 11308 5540 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 6012 11308 8861 11336
rect 6012 11277 6040 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 12342 11336 12348 11348
rect 9088 11308 12348 11336
rect 9088 11296 9094 11308
rect 12342 11296 12348 11308
rect 12400 11336 12406 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12400 11308 12449 11336
rect 12400 11296 12406 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 12437 11299 12495 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14550 11336 14556 11348
rect 13955 11308 14556 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14550 11296 14556 11308
rect 14608 11336 14614 11348
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14608 11308 14841 11336
rect 14608 11296 14614 11308
rect 14829 11305 14841 11308
rect 14875 11336 14887 11339
rect 14918 11336 14924 11348
rect 14875 11308 14924 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16666 11296 16672 11308
rect 16724 11336 16730 11348
rect 18141 11339 18199 11345
rect 16724 11308 17632 11336
rect 16724 11296 16730 11308
rect 3099 11271 3157 11277
rect 3099 11237 3111 11271
rect 3145 11268 3157 11271
rect 5997 11271 6055 11277
rect 5997 11268 6009 11271
rect 3145 11240 6009 11268
rect 3145 11237 3157 11240
rect 3099 11231 3157 11237
rect 5997 11237 6009 11240
rect 6043 11237 6055 11271
rect 5997 11231 6055 11237
rect 6098 11271 6156 11277
rect 6098 11237 6110 11271
rect 6144 11268 6156 11271
rect 6362 11268 6368 11280
rect 6144 11240 6368 11268
rect 6144 11237 6156 11240
rect 6098 11231 6156 11237
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 6454 11228 6460 11280
rect 6512 11268 6518 11280
rect 7285 11271 7343 11277
rect 7285 11268 7297 11271
rect 6512 11240 7297 11268
rect 6512 11228 6518 11240
rect 7285 11237 7297 11240
rect 7331 11237 7343 11271
rect 7285 11231 7343 11237
rect 7653 11271 7711 11277
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7834 11268 7840 11280
rect 7699 11240 7840 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7834 11228 7840 11240
rect 7892 11228 7898 11280
rect 9858 11268 9864 11280
rect 9819 11240 9864 11268
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 10137 11271 10195 11277
rect 10137 11268 10149 11271
rect 10008 11240 10149 11268
rect 10008 11228 10014 11240
rect 10137 11237 10149 11240
rect 10183 11237 10195 11271
rect 10137 11231 10195 11237
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11268 10287 11271
rect 10594 11268 10600 11280
rect 10275 11240 10600 11268
rect 10275 11237 10287 11240
rect 10229 11231 10287 11237
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 10781 11271 10839 11277
rect 10781 11237 10793 11271
rect 10827 11268 10839 11271
rect 11422 11268 11428 11280
rect 10827 11240 11428 11268
rect 10827 11237 10839 11240
rect 10781 11231 10839 11237
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 15378 11268 15384 11280
rect 15339 11240 15384 11268
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 17604 11277 17632 11308
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 18230 11336 18236 11348
rect 18187 11308 18236 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 18506 11336 18512 11348
rect 18467 11308 18512 11336
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 20622 11336 20628 11348
rect 20583 11308 20628 11336
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 17037 11271 17095 11277
rect 17037 11268 17049 11271
rect 15528 11240 17049 11268
rect 15528 11228 15534 11240
rect 17037 11237 17049 11240
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 17589 11271 17647 11277
rect 17589 11237 17601 11271
rect 17635 11237 17647 11271
rect 21082 11268 21088 11280
rect 21043 11240 21088 11268
rect 17589 11231 17647 11237
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 1302 11160 1308 11212
rect 1360 11200 1366 11212
rect 1489 11203 1547 11209
rect 1489 11200 1501 11203
rect 1360 11172 1501 11200
rect 1360 11160 1366 11172
rect 1489 11169 1501 11172
rect 1535 11169 1547 11203
rect 1489 11163 1547 11169
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 2996 11203 3054 11209
rect 2996 11200 3008 11203
rect 2924 11172 3008 11200
rect 2924 11160 2930 11172
rect 2996 11169 3008 11172
rect 3042 11169 3054 11203
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 2996 11163 3054 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 11974 11200 11980 11212
rect 11935 11172 11980 11200
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12115 11203 12173 11209
rect 12115 11169 12127 11203
rect 12161 11200 12173 11203
rect 12161 11172 13814 11200
rect 12161 11169 12173 11172
rect 12115 11163 12173 11169
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2314 11132 2320 11144
rect 2179 11104 2320 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 2777 11135 2835 11141
rect 2777 11132 2789 11135
rect 2372 11104 2789 11132
rect 2372 11092 2378 11104
rect 2777 11101 2789 11104
rect 2823 11101 2835 11135
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 2777 11095 2835 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 7374 11132 7380 11144
rect 6425 11104 7380 11132
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 2406 11064 2412 11076
rect 1636 11036 2412 11064
rect 1636 11024 1642 11036
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 4154 11064 4160 11076
rect 3844 11036 4160 11064
rect 3844 11024 3850 11036
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 6425 11064 6453 11104
rect 7374 11092 7380 11104
rect 7432 11132 7438 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7432 11104 7573 11132
rect 7432 11092 7438 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8018 11132 8024 11144
rect 7883 11104 8024 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 4488 11036 6453 11064
rect 6549 11067 6607 11073
rect 4488 11024 4494 11036
rect 6549 11033 6561 11067
rect 6595 11064 6607 11067
rect 7852 11064 7880 11095
rect 8018 11092 8024 11104
rect 8076 11132 8082 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8076 11104 9229 11132
rect 8076 11092 8082 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 13786 11132 13814 11172
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18414 11200 18420 11212
rect 17920 11172 18420 11200
rect 17920 11160 17926 11172
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 16758 11132 16764 11144
rect 13786 11104 16764 11132
rect 12989 11095 13047 11101
rect 6595 11036 7880 11064
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 10962 11064 10968 11076
rect 8996 11036 10968 11064
rect 8996 11024 9002 11036
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 13004 11008 13032 11095
rect 16758 11092 16764 11104
rect 16816 11132 16822 11144
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 16816 11104 16957 11132
rect 16816 11092 16822 11104
rect 16945 11101 16957 11104
rect 16991 11101 17003 11135
rect 16945 11095 17003 11101
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 18892 11132 18920 11163
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 22500 11203 22558 11209
rect 22500 11200 22512 11203
rect 22336 11172 22512 11200
rect 22336 11160 22342 11172
rect 22500 11169 22512 11172
rect 22546 11200 22558 11203
rect 23106 11200 23112 11212
rect 22546 11172 23112 11200
rect 22546 11169 22558 11172
rect 22500 11163 22558 11169
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 17644 11104 19625 11132
rect 17644 11092 17650 11104
rect 19613 11101 19625 11104
rect 19659 11132 19671 11135
rect 20070 11132 20076 11144
rect 19659 11104 20076 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 20070 11092 20076 11104
rect 20128 11092 20134 11144
rect 20438 11092 20444 11144
rect 20496 11132 20502 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20496 11104 21005 11132
rect 20496 11092 20502 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11132 21695 11135
rect 22002 11132 22008 11144
rect 21683 11104 22008 11132
rect 21683 11101 21695 11104
rect 21637 11095 21695 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23532 11104 23577 11132
rect 23532 11092 23538 11104
rect 15930 11064 15936 11076
rect 15891 11036 15936 11064
rect 15930 11024 15936 11036
rect 15988 11024 15994 11076
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 22186 11064 22192 11076
rect 17184 11036 22192 11064
rect 17184 11024 17190 11036
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3384 10968 3433 10996
rect 3384 10956 3390 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 5534 10996 5540 11008
rect 5495 10968 5540 10996
rect 3421 10959 3479 10965
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 6696 10968 6929 10996
rect 6696 10956 6702 10968
rect 6917 10965 6929 10968
rect 6963 10965 6975 10999
rect 6917 10959 6975 10965
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 8481 10999 8539 11005
rect 8481 10996 8493 10999
rect 7064 10968 8493 10996
rect 7064 10956 7070 10968
rect 8481 10965 8493 10968
rect 8527 10965 8539 10999
rect 8481 10959 8539 10965
rect 12897 10999 12955 11005
rect 12897 10965 12909 10999
rect 12943 10996 12955 10999
rect 12986 10996 12992 11008
rect 12943 10968 12992 10996
rect 12943 10965 12955 10968
rect 12897 10959 12955 10965
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 14148 10968 14289 10996
rect 14148 10956 14154 10968
rect 14277 10965 14289 10968
rect 14323 10996 14335 10999
rect 19058 10996 19064 11008
rect 14323 10968 19064 10996
rect 14323 10965 14335 10968
rect 14277 10959 14335 10965
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 22603 10999 22661 11005
rect 22603 10996 22615 10999
rect 21048 10968 22615 10996
rect 21048 10956 21054 10968
rect 22603 10965 22615 10968
rect 22649 10965 22661 10999
rect 22603 10959 22661 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 1946 10792 1952 10804
rect 1535 10764 1952 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 1946 10752 1952 10764
rect 2004 10792 2010 10804
rect 3418 10792 3424 10804
rect 2004 10764 3424 10792
rect 2004 10752 2010 10764
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4338 10792 4344 10804
rect 4295 10764 4344 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 5074 10792 5080 10804
rect 5035 10764 5080 10792
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 10008 10764 11345 10792
rect 10008 10752 10014 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 12667 10795 12725 10801
rect 12667 10761 12679 10795
rect 12713 10792 12725 10795
rect 14642 10792 14648 10804
rect 12713 10764 14648 10792
rect 12713 10761 12725 10764
rect 12667 10755 12725 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15436 10764 16313 10792
rect 15436 10752 15442 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 18472 10764 19257 10792
rect 18472 10752 18478 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 19245 10755 19303 10761
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10792 20775 10795
rect 21082 10792 21088 10804
rect 20763 10764 21088 10792
rect 20763 10761 20775 10764
rect 20717 10755 20775 10761
rect 21082 10752 21088 10764
rect 21140 10752 21146 10804
rect 9493 10727 9551 10733
rect 9493 10693 9505 10727
rect 9539 10724 9551 10727
rect 10594 10724 10600 10736
rect 9539 10696 10600 10724
rect 9539 10693 9551 10696
rect 9493 10687 9551 10693
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 13354 10724 13360 10736
rect 13315 10696 13360 10724
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 14550 10684 14556 10736
rect 14608 10724 14614 10736
rect 14737 10727 14795 10733
rect 14737 10724 14749 10727
rect 14608 10696 14749 10724
rect 14608 10684 14614 10696
rect 14737 10693 14749 10696
rect 14783 10724 14795 10727
rect 15470 10724 15476 10736
rect 14783 10696 15476 10724
rect 14783 10693 14795 10696
rect 14737 10687 14795 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 15930 10724 15936 10736
rect 15891 10696 15936 10724
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 17083 10727 17141 10733
rect 17083 10693 17095 10727
rect 17129 10724 17141 10727
rect 24762 10724 24768 10736
rect 17129 10696 21680 10724
rect 24723 10696 24768 10724
rect 17129 10693 17141 10696
rect 17083 10687 17141 10693
rect 3050 10616 3056 10668
rect 3108 10656 3114 10668
rect 4614 10656 4620 10668
rect 3108 10628 4620 10656
rect 3108 10616 3114 10628
rect 4614 10616 4620 10628
rect 4672 10656 4678 10668
rect 5534 10656 5540 10668
rect 4672 10628 5540 10656
rect 4672 10616 4678 10628
rect 5534 10616 5540 10628
rect 5592 10656 5598 10668
rect 8478 10656 8484 10668
rect 5592 10628 8484 10656
rect 5592 10616 5598 10628
rect 1670 10588 1676 10600
rect 1631 10560 1676 10588
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1912 10560 1961 10588
rect 1912 10548 1918 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5736 10597 5764 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 9122 10656 9128 10668
rect 9083 10628 9128 10656
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 9876 10628 10977 10656
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 5132 10560 5181 10588
rect 5132 10548 5138 10560
rect 5169 10557 5181 10560
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8260 10560 8401 10588
rect 8260 10548 8266 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8938 10588 8944 10600
rect 8899 10560 8944 10588
rect 8389 10551 8447 10557
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 3050 10520 3056 10532
rect 3011 10492 3056 10520
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 3145 10523 3203 10529
rect 3145 10489 3157 10523
rect 3191 10520 3203 10523
rect 3694 10520 3700 10532
rect 3191 10492 3556 10520
rect 3655 10492 3700 10520
rect 3191 10489 3203 10492
rect 3145 10483 3203 10489
rect 1302 10412 1308 10464
rect 1360 10452 1366 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 1360 10424 2421 10452
rect 1360 10412 1366 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2866 10452 2872 10464
rect 2827 10424 2872 10452
rect 2409 10415 2467 10421
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 3528 10452 3556 10492
rect 3694 10480 3700 10492
rect 3752 10480 3758 10532
rect 5905 10523 5963 10529
rect 4126 10492 5212 10520
rect 4126 10452 4154 10492
rect 5184 10464 5212 10492
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 6086 10520 6092 10532
rect 5951 10492 6092 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 6086 10480 6092 10492
rect 6144 10480 6150 10532
rect 6914 10520 6920 10532
rect 6875 10492 6920 10520
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 7009 10523 7067 10529
rect 7009 10489 7021 10523
rect 7055 10489 7067 10523
rect 7558 10520 7564 10532
rect 7519 10492 7564 10520
rect 7009 10483 7067 10489
rect 3528 10424 4154 10452
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 5224 10424 6193 10452
rect 5224 10412 5230 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6181 10415 6239 10421
rect 6546 10412 6552 10424
rect 6604 10452 6610 10464
rect 7024 10452 7052 10483
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 7929 10523 7987 10529
rect 7929 10489 7941 10523
rect 7975 10520 7987 10523
rect 8110 10520 8116 10532
rect 7975 10492 8116 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 8110 10480 8116 10492
rect 8168 10520 8174 10532
rect 8956 10520 8984 10548
rect 8168 10492 8984 10520
rect 8168 10480 8174 10492
rect 9582 10480 9588 10532
rect 9640 10520 9646 10532
rect 9876 10520 9904 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10656 13691 10659
rect 14090 10656 14096 10668
rect 13679 10628 14096 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 14274 10656 14280 10668
rect 14235 10628 14280 10656
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 15562 10656 15568 10668
rect 15243 10628 15568 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 15562 10616 15568 10628
rect 15620 10656 15626 10668
rect 16761 10659 16819 10665
rect 16761 10656 16773 10659
rect 15620 10628 16773 10656
rect 15620 10616 15626 10628
rect 16761 10625 16773 10628
rect 16807 10625 16819 10659
rect 16761 10619 16819 10625
rect 17218 10616 17224 10668
rect 17276 10656 17282 10668
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17276 10628 18061 10656
rect 17276 10616 17282 10628
rect 18049 10625 18061 10628
rect 18095 10656 18107 10659
rect 18506 10656 18512 10668
rect 18095 10628 18512 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10656 19855 10659
rect 19978 10656 19984 10668
rect 19843 10628 19984 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 21652 10665 21680 10696
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 21910 10656 21916 10668
rect 21683 10628 21916 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 22002 10616 22008 10668
rect 22060 10656 22066 10668
rect 22060 10628 22105 10656
rect 22060 10616 22066 10628
rect 12596 10591 12654 10597
rect 12596 10557 12608 10591
rect 12642 10588 12654 10591
rect 12710 10588 12716 10600
rect 12642 10560 12716 10588
rect 12642 10557 12654 10560
rect 12596 10551 12654 10557
rect 12710 10548 12716 10560
rect 12768 10588 12774 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12768 10560 13001 10588
rect 12768 10548 12774 10560
rect 12989 10557 13001 10560
rect 13035 10588 13047 10591
rect 16850 10588 16856 10600
rect 13035 10560 13400 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 10045 10523 10103 10529
rect 10045 10520 10057 10523
rect 9640 10492 10057 10520
rect 9640 10480 9646 10492
rect 10045 10489 10057 10492
rect 10091 10489 10103 10523
rect 10045 10483 10103 10489
rect 10137 10523 10195 10529
rect 10137 10489 10149 10523
rect 10183 10489 10195 10523
rect 10686 10520 10692 10532
rect 10647 10492 10692 10520
rect 10137 10483 10195 10489
rect 9858 10452 9864 10464
rect 6604 10424 7052 10452
rect 9771 10424 9864 10452
rect 6604 10412 6610 10424
rect 9858 10412 9864 10424
rect 9916 10452 9922 10464
rect 10152 10452 10180 10483
rect 10686 10480 10692 10492
rect 10744 10480 10750 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 12032 10492 12081 10520
rect 12032 10480 12038 10492
rect 12069 10489 12081 10492
rect 12115 10520 12127 10523
rect 13078 10520 13084 10532
rect 12115 10492 13084 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 13372 10520 13400 10560
rect 16408 10560 16856 10588
rect 13722 10520 13728 10532
rect 13372 10492 13492 10520
rect 13683 10492 13728 10520
rect 9916 10424 10180 10452
rect 13464 10452 13492 10492
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 15378 10520 15384 10532
rect 15339 10492 15384 10520
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 15528 10492 15573 10520
rect 15528 10480 15534 10492
rect 16408 10452 16436 10560
rect 16850 10548 16856 10560
rect 16908 10588 16914 10600
rect 16980 10591 17038 10597
rect 16980 10588 16992 10591
rect 16908 10560 16992 10588
rect 16908 10548 16914 10560
rect 16980 10557 16992 10560
rect 17026 10588 17038 10591
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 17026 10560 17417 10588
rect 17026 10557 17038 10560
rect 16980 10551 17038 10557
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19058 10588 19064 10600
rect 19015 10560 19064 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19058 10548 19064 10560
rect 19116 10588 19122 10600
rect 19116 10560 21496 10588
rect 19116 10548 19122 10560
rect 18370 10523 18428 10529
rect 18370 10489 18382 10523
rect 18416 10489 18428 10523
rect 18370 10483 18428 10489
rect 20118 10523 20176 10529
rect 20118 10489 20130 10523
rect 20164 10489 20176 10523
rect 20118 10483 20176 10489
rect 17770 10452 17776 10464
rect 13464 10424 16436 10452
rect 17731 10424 17776 10452
rect 9916 10412 9922 10424
rect 17770 10412 17776 10424
rect 17828 10452 17834 10464
rect 18385 10452 18413 10483
rect 19150 10452 19156 10464
rect 17828 10424 19156 10452
rect 17828 10412 17834 10424
rect 19150 10412 19156 10424
rect 19208 10452 19214 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19208 10424 19625 10452
rect 19208 10412 19214 10424
rect 19613 10421 19625 10424
rect 19659 10452 19671 10455
rect 20133 10452 20161 10483
rect 21468 10461 21496 10560
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24176 10560 24593 10588
rect 24176 10548 24182 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24627 10560 25145 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 21729 10523 21787 10529
rect 21729 10489 21741 10523
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 19659 10424 20161 10452
rect 21453 10455 21511 10461
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 21453 10421 21465 10455
rect 21499 10452 21511 10455
rect 21744 10452 21772 10483
rect 21499 10424 21772 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22557 10455 22615 10461
rect 22557 10452 22569 10455
rect 22336 10424 22569 10452
rect 22336 10412 22342 10424
rect 22557 10421 22569 10424
rect 22603 10421 22615 10455
rect 22557 10415 22615 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2225 10251 2283 10257
rect 2225 10248 2237 10251
rect 1728 10220 2237 10248
rect 1728 10208 1734 10220
rect 2225 10217 2237 10220
rect 2271 10217 2283 10251
rect 2225 10211 2283 10217
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 3108 10220 4261 10248
rect 3108 10208 3114 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 6454 10248 6460 10260
rect 5675 10220 6460 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6604 10220 6684 10248
rect 6604 10208 6610 10220
rect 3142 10180 3148 10192
rect 2516 10152 3148 10180
rect 2516 10124 2544 10152
rect 3142 10140 3148 10152
rect 3200 10140 3206 10192
rect 3418 10180 3424 10192
rect 3379 10152 3424 10180
rect 3418 10140 3424 10152
rect 3476 10180 3482 10192
rect 3789 10183 3847 10189
rect 3789 10180 3801 10183
rect 3476 10152 3801 10180
rect 3476 10140 3482 10152
rect 3789 10149 3801 10152
rect 3835 10149 3847 10183
rect 3789 10143 3847 10149
rect 5071 10183 5129 10189
rect 5071 10149 5083 10183
rect 5117 10180 5129 10183
rect 5534 10180 5540 10192
rect 5117 10152 5540 10180
rect 5117 10149 5129 10152
rect 5071 10143 5129 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 6656 10189 6684 10220
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 7469 10251 7527 10257
rect 7469 10248 7481 10251
rect 7432 10220 7481 10248
rect 7432 10208 7438 10220
rect 7469 10217 7481 10220
rect 7515 10217 7527 10251
rect 7834 10248 7840 10260
rect 7795 10220 7840 10248
rect 7469 10211 7527 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 12986 10248 12992 10260
rect 9646 10220 11560 10248
rect 12947 10220 12992 10248
rect 6641 10183 6699 10189
rect 6641 10149 6653 10183
rect 6687 10149 6699 10183
rect 6641 10143 6699 10149
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 9214 10180 9220 10192
rect 6880 10152 9220 10180
rect 6880 10140 6886 10152
rect 9214 10140 9220 10152
rect 9272 10180 9278 10192
rect 9646 10180 9674 10220
rect 9950 10180 9956 10192
rect 9272 10152 9674 10180
rect 9911 10152 9956 10180
rect 9272 10140 9278 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 11532 10189 11560 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13722 10208 13728 10260
rect 13780 10248 13786 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13780 10220 13921 10248
rect 13780 10208 13786 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 15381 10251 15439 10257
rect 15381 10248 15393 10251
rect 14700 10220 15393 10248
rect 14700 10208 14706 10220
rect 15381 10217 15393 10220
rect 15427 10217 15439 10251
rect 16758 10248 16764 10260
rect 16719 10220 16764 10248
rect 15381 10211 15439 10217
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 17218 10248 17224 10260
rect 17179 10220 17224 10248
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20438 10208 20444 10260
rect 20496 10248 20502 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20496 10220 20637 10248
rect 20496 10208 20502 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 21910 10248 21916 10260
rect 21871 10220 21916 10248
rect 20625 10211 20683 10217
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 11517 10183 11575 10189
rect 11517 10149 11529 10183
rect 11563 10180 11575 10183
rect 11698 10180 11704 10192
rect 11563 10152 11704 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 18414 10180 18420 10192
rect 12912 10152 18420 10180
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2038 10112 2044 10124
rect 1510 10084 2044 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 2958 10112 2964 10124
rect 2919 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 4246 10112 4252 10124
rect 4126 10084 4252 10112
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 4126 10044 4154 10084
rect 4246 10072 4252 10084
rect 4304 10112 4310 10124
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 4304 10084 5917 10112
rect 4304 10072 4310 10084
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 8018 10112 8024 10124
rect 7248 10084 8024 10112
rect 7248 10072 7254 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8478 10112 8484 10124
rect 8439 10084 8484 10112
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 12912 10121 12940 10152
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 19058 10180 19064 10192
rect 19019 10152 19064 10180
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 21082 10180 21088 10192
rect 21043 10152 21088 10180
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12676 10084 12909 10112
rect 12676 10072 12682 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 13354 10112 13360 10124
rect 13315 10084 13360 10112
rect 12897 10075 12955 10081
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 14792 10084 15301 10112
rect 14792 10072 14798 10084
rect 15289 10081 15301 10084
rect 15335 10112 15347 10115
rect 15654 10112 15660 10124
rect 15335 10084 15660 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 17310 10112 17316 10124
rect 17271 10084 17316 10112
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 17773 10115 17831 10121
rect 17773 10112 17785 10115
rect 17644 10084 17785 10112
rect 17644 10072 17650 10084
rect 17773 10081 17785 10084
rect 17819 10112 17831 10115
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 17819 10084 18521 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 22462 10112 22468 10124
rect 22520 10121 22526 10124
rect 22520 10115 22558 10121
rect 22410 10084 22468 10112
rect 18509 10075 18567 10081
rect 22462 10072 22468 10084
rect 22546 10112 22558 10115
rect 24210 10112 24216 10124
rect 22546 10084 24216 10112
rect 22546 10081 22558 10084
rect 22520 10075 22558 10081
rect 22520 10072 22526 10075
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 4706 10044 4712 10056
rect 3191 10016 4154 10044
rect 4667 10016 4712 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 8754 10044 8760 10056
rect 6595 10016 7598 10044
rect 8715 10016 8760 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 1535 9979 1593 9985
rect 1535 9945 1547 9979
rect 1581 9976 1593 9979
rect 6564 9976 6592 10007
rect 1581 9948 6592 9976
rect 1581 9945 1593 9948
rect 1535 9939 1593 9945
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 7064 9948 7113 9976
rect 7064 9936 7070 9948
rect 7101 9945 7113 9948
rect 7147 9945 7159 9979
rect 7570 9976 7598 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9732 10016 9873 10044
rect 9732 10004 9738 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 11422 10044 11428 10056
rect 11383 10016 11428 10044
rect 10137 10007 10195 10013
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 7570 9948 9045 9976
rect 7101 9939 7159 9945
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 10152 9976 10180 10007
rect 11422 10004 11428 10016
rect 11480 10004 11486 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11572 10016 11713 10044
rect 11572 10004 11578 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 11701 10007 11759 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 18966 10044 18972 10056
rect 18927 10016 18972 10044
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 19610 10044 19616 10056
rect 19571 10016 19616 10044
rect 19610 10004 19616 10016
rect 19668 10004 19674 10056
rect 20990 10044 20996 10056
rect 20951 10016 20996 10044
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21266 10044 21272 10056
rect 21227 10016 21272 10044
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 11054 9976 11060 9988
rect 9033 9939 9091 9945
rect 9140 9948 11060 9976
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 6362 9908 6368 9920
rect 6275 9880 6368 9908
rect 6362 9868 6368 9880
rect 6420 9908 6426 9920
rect 6822 9908 6828 9920
rect 6420 9880 6828 9908
rect 6420 9868 6426 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7116 9908 7144 9939
rect 9140 9908 9168 9948
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 7116 9880 9168 9908
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 10686 9908 10692 9920
rect 9539 9880 10692 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 10962 9908 10968 9920
rect 10919 9880 10968 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14792 9880 15025 9908
rect 14792 9868 14798 9880
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15378 9908 15384 9920
rect 15059 9880 15384 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16482 9908 16488 9920
rect 16443 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22603 9911 22661 9917
rect 22603 9908 22615 9911
rect 22152 9880 22615 9908
rect 22152 9868 22158 9880
rect 22603 9877 22615 9880
rect 22649 9877 22661 9911
rect 22603 9871 22661 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 4706 9664 4712 9716
rect 4764 9704 4770 9716
rect 5813 9707 5871 9713
rect 5813 9704 5825 9707
rect 4764 9676 5825 9704
rect 4764 9664 4770 9676
rect 5813 9673 5825 9676
rect 5859 9673 5871 9707
rect 6454 9704 6460 9716
rect 6415 9676 6460 9704
rect 5813 9667 5871 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 8018 9704 8024 9716
rect 7979 9676 8024 9704
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 9858 9704 9864 9716
rect 9819 9676 9864 9704
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10134 9704 10140 9716
rect 10008 9676 10140 9704
rect 10008 9664 10014 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 11698 9704 11704 9716
rect 11659 9676 11704 9704
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12253 9707 12311 9713
rect 12253 9673 12265 9707
rect 12299 9704 12311 9707
rect 13354 9704 13360 9716
rect 12299 9676 13360 9704
rect 12299 9673 12311 9676
rect 12253 9667 12311 9673
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15712 9676 15761 9704
rect 15712 9664 15718 9676
rect 15749 9673 15761 9676
rect 15795 9673 15807 9707
rect 15749 9667 15807 9673
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 16117 9707 16175 9713
rect 16117 9704 16129 9707
rect 15896 9676 16129 9704
rect 15896 9664 15902 9676
rect 16117 9673 16129 9676
rect 16163 9673 16175 9707
rect 17310 9704 17316 9716
rect 16117 9667 16175 9673
rect 16316 9676 17316 9704
rect 1627 9639 1685 9645
rect 1627 9605 1639 9639
rect 1673 9636 1685 9639
rect 5166 9636 5172 9648
rect 1673 9608 5028 9636
rect 5127 9608 5172 9636
rect 1673 9605 1685 9608
rect 1627 9599 1685 9605
rect 4246 9568 4252 9580
rect 4207 9540 4252 9568
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 5000 9568 5028 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 9876 9636 9904 9664
rect 10505 9639 10563 9645
rect 10505 9636 10517 9639
rect 9876 9608 10517 9636
rect 10505 9605 10517 9608
rect 10551 9636 10563 9639
rect 10870 9636 10876 9648
rect 10551 9608 10876 9636
rect 10551 9605 10563 9608
rect 10505 9599 10563 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 11112 9608 11345 9636
rect 11112 9596 11118 9608
rect 11333 9605 11345 9608
rect 11379 9605 11391 9639
rect 11333 9599 11391 9605
rect 13538 9596 13544 9648
rect 13596 9636 13602 9648
rect 13596 9608 13814 9636
rect 13596 9596 13602 9608
rect 6822 9568 6828 9580
rect 5000 9540 6828 9568
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7466 9568 7472 9580
rect 7055 9540 7472 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8812 9540 8953 9568
rect 8812 9528 8818 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 13786 9568 13814 9608
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 16316 9636 16344 9676
rect 17310 9664 17316 9676
rect 17368 9704 17374 9716
rect 17405 9707 17463 9713
rect 17405 9704 17417 9707
rect 17368 9676 17417 9704
rect 17368 9664 17374 9676
rect 17405 9673 17417 9676
rect 17451 9673 17463 9707
rect 17405 9667 17463 9673
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 19245 9707 19303 9713
rect 19245 9704 19257 9707
rect 19116 9676 19257 9704
rect 19116 9664 19122 9676
rect 19245 9673 19257 9676
rect 19291 9673 19303 9707
rect 19245 9667 19303 9673
rect 20993 9707 21051 9713
rect 20993 9673 21005 9707
rect 21039 9704 21051 9707
rect 21082 9704 21088 9716
rect 21039 9676 21088 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 22462 9704 22468 9716
rect 22423 9676 22468 9704
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 15252 9608 16344 9636
rect 15252 9596 15258 9608
rect 19610 9596 19616 9648
rect 19668 9636 19674 9648
rect 20441 9639 20499 9645
rect 20441 9636 20453 9639
rect 19668 9608 20453 9636
rect 19668 9596 19674 9608
rect 20441 9605 20453 9608
rect 20487 9636 20499 9639
rect 21266 9636 21272 9648
rect 20487 9608 21272 9636
rect 20487 9605 20499 9608
rect 20441 9599 20499 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 21450 9596 21456 9648
rect 21508 9636 21514 9648
rect 22833 9639 22891 9645
rect 22833 9636 22845 9639
rect 21508 9608 22845 9636
rect 21508 9596 21514 9608
rect 22833 9605 22845 9608
rect 22879 9605 22891 9639
rect 22833 9599 22891 9605
rect 22922 9596 22928 9648
rect 22980 9636 22986 9648
rect 23799 9639 23857 9645
rect 23799 9636 23811 9639
rect 22980 9608 23811 9636
rect 22980 9596 22986 9608
rect 23799 9605 23811 9608
rect 23845 9605 23857 9639
rect 23799 9599 23857 9605
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13786 9540 13921 9568
rect 8941 9531 8999 9537
rect 13909 9537 13921 9540
rect 13955 9568 13967 9571
rect 17218 9568 17224 9580
rect 13955 9540 17224 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 18046 9568 18052 9580
rect 18007 9540 18052 9568
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20254 9568 20260 9580
rect 19935 9540 20260 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20254 9528 20260 9540
rect 20312 9568 20318 9580
rect 22094 9568 22100 9580
rect 20312 9540 22100 9568
rect 20312 9528 20318 9540
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 24118 9568 24124 9580
rect 24079 9540 24124 9568
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2222 9500 2228 9512
rect 2096 9472 2228 9500
rect 2096 9460 2102 9472
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2498 9500 2504 9512
rect 2459 9472 2504 9500
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 8849 9503 8907 9509
rect 2648 9472 6868 9500
rect 2648 9460 2654 9472
rect 2863 9435 2921 9441
rect 2863 9401 2875 9435
rect 2909 9432 2921 9435
rect 3789 9435 3847 9441
rect 3789 9432 3801 9435
rect 2909 9404 3801 9432
rect 2909 9401 2921 9404
rect 2863 9395 2921 9401
rect 3789 9401 3801 9404
rect 3835 9432 3847 9435
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 3835 9404 4077 9432
rect 3835 9401 3847 9404
rect 3789 9395 3847 9401
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 4065 9395 4123 9401
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 4570 9435 4628 9441
rect 4570 9432 4582 9435
rect 4203 9404 4582 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4570 9401 4582 9404
rect 4616 9432 4628 9435
rect 4798 9432 4804 9444
rect 4616 9404 4804 9432
rect 4616 9401 4628 9404
rect 4570 9395 4628 9401
rect 4798 9392 4804 9404
rect 4856 9432 4862 9444
rect 5445 9435 5503 9441
rect 5445 9432 5457 9435
rect 4856 9404 5457 9432
rect 4856 9392 4862 9404
rect 5445 9401 5457 9404
rect 5491 9432 5503 9435
rect 5534 9432 5540 9444
rect 5491 9404 5540 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 2958 9364 2964 9376
rect 2648 9336 2964 9364
rect 2648 9324 2654 9336
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 6840 9364 6868 9472
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 18969 9503 19027 9509
rect 8895 9472 9076 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 7156 9404 7201 9432
rect 7156 9392 7162 9404
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7653 9435 7711 9441
rect 7653 9432 7665 9435
rect 7340 9404 7665 9432
rect 7340 9392 7346 9404
rect 7653 9401 7665 9404
rect 7699 9432 7711 9435
rect 9048 9432 9076 9472
rect 18969 9469 18981 9503
rect 19015 9500 19027 9503
rect 23728 9503 23786 9509
rect 19015 9472 19748 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 9303 9435 9361 9441
rect 9303 9432 9315 9435
rect 7699 9404 8984 9432
rect 9048 9404 9315 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 7834 9364 7840 9376
rect 6840 9336 7840 9364
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8956 9364 8984 9404
rect 9303 9401 9315 9404
rect 9349 9432 9361 9435
rect 9950 9432 9956 9444
rect 9349 9404 9956 9432
rect 9349 9401 9361 9404
rect 9303 9395 9361 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 10778 9432 10784 9444
rect 10739 9404 10784 9432
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 10928 9404 10973 9432
rect 10928 9392 10934 9404
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13265 9435 13323 9441
rect 13265 9432 13277 9435
rect 12860 9404 13277 9432
rect 12860 9392 12866 9404
rect 13265 9401 13277 9404
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 13357 9435 13415 9441
rect 13357 9401 13369 9435
rect 13403 9432 13415 9435
rect 14826 9432 14832 9444
rect 13403 9404 13814 9432
rect 14787 9404 14832 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 13786 9376 13814 9404
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 15470 9432 15476 9444
rect 14976 9404 15021 9432
rect 15431 9404 15476 9432
rect 14976 9392 14982 9404
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 16482 9432 16488 9444
rect 16443 9404 16488 9432
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 17129 9435 17187 9441
rect 16632 9404 16677 9432
rect 16632 9392 16638 9404
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 18230 9432 18236 9444
rect 17175 9404 18236 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 18370 9435 18428 9441
rect 18370 9401 18382 9435
rect 18416 9401 18428 9435
rect 18370 9395 18428 9401
rect 11606 9364 11612 9376
rect 8956 9336 11612 9364
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12676 9336 12909 9364
rect 12676 9324 12682 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 13722 9324 13728 9376
rect 13780 9364 13814 9376
rect 14182 9364 14188 9376
rect 13780 9336 14188 9364
rect 13780 9324 13786 9336
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14550 9364 14556 9376
rect 14511 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17770 9364 17776 9376
rect 17368 9336 17776 9364
rect 17368 9324 17374 9336
rect 17770 9324 17776 9336
rect 17828 9364 17834 9376
rect 18385 9364 18413 9395
rect 19720 9373 19748 9472
rect 23728 9469 23740 9503
rect 23774 9500 23786 9503
rect 24136 9500 24164 9528
rect 23774 9472 24164 9500
rect 23774 9469 23786 9472
rect 23728 9463 23786 9469
rect 19981 9435 20039 9441
rect 19981 9401 19993 9435
rect 20027 9401 20039 9435
rect 21450 9432 21456 9444
rect 21411 9404 21456 9432
rect 19981 9395 20039 9401
rect 17828 9336 18413 9364
rect 19705 9367 19763 9373
rect 17828 9324 17834 9336
rect 19705 9333 19717 9367
rect 19751 9364 19763 9367
rect 19996 9364 20024 9395
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 22094 9432 22100 9444
rect 21600 9404 21645 9432
rect 22055 9404 22100 9432
rect 21600 9392 21606 9404
rect 22094 9392 22100 9404
rect 22152 9392 22158 9444
rect 21560 9364 21588 9392
rect 19751 9336 21588 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9160 2562 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 2556 9132 5917 9160
rect 2556 9120 2562 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 5905 9123 5963 9129
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7098 9160 7104 9172
rect 7055 9132 7104 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7098 9120 7104 9132
rect 7156 9160 7162 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7156 9132 7297 9160
rect 7156 9120 7162 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8812 9132 9045 9160
rect 8812 9120 8818 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10192 9132 10609 9160
rect 10192 9120 10198 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11563 9163 11621 9169
rect 11563 9160 11575 9163
rect 11480 9132 11575 9160
rect 11480 9120 11486 9132
rect 11563 9129 11575 9132
rect 11609 9160 11621 9163
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11609 9132 11897 9160
rect 11609 9129 11621 9132
rect 11563 9123 11621 9129
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 13817 9163 13875 9169
rect 13817 9160 13829 9163
rect 13780 9132 13829 9160
rect 13780 9120 13786 9132
rect 13817 9129 13829 9132
rect 13863 9129 13875 9163
rect 13817 9123 13875 9129
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 18104 9132 18245 9160
rect 18104 9120 18110 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19797 9163 19855 9169
rect 19797 9160 19809 9163
rect 19024 9132 19809 9160
rect 19024 9120 19030 9132
rect 19797 9129 19809 9132
rect 19843 9129 19855 9163
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 19797 9123 19855 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20717 9163 20775 9169
rect 20717 9129 20729 9163
rect 20763 9160 20775 9163
rect 20990 9160 20996 9172
rect 20763 9132 20996 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21600 9132 21925 9160
rect 21600 9120 21606 9132
rect 21913 9129 21925 9132
rect 21959 9129 21971 9163
rect 21913 9123 21971 9129
rect 4433 9095 4491 9101
rect 4433 9061 4445 9095
rect 4479 9092 4491 9095
rect 4706 9092 4712 9104
rect 4479 9064 4712 9092
rect 4479 9061 4491 9064
rect 4433 9055 4491 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 6410 9095 6468 9101
rect 6410 9092 6422 9095
rect 5592 9064 6422 9092
rect 5592 9052 5598 9064
rect 6410 9061 6422 9064
rect 6456 9092 6468 9095
rect 6638 9092 6644 9104
rect 6456 9064 6644 9092
rect 6456 9061 6468 9064
rect 6410 9055 6468 9061
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 9401 9095 9459 9101
rect 9401 9092 9413 9095
rect 6880 9064 9413 9092
rect 6880 9052 6886 9064
rect 9401 9061 9413 9064
rect 9447 9092 9459 9095
rect 9674 9092 9680 9104
rect 9447 9064 9680 9092
rect 9447 9061 9459 9064
rect 9401 9055 9459 9061
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13262 9101 13268 9104
rect 13218 9095 13268 9101
rect 13218 9092 13230 9095
rect 13044 9064 13230 9092
rect 13044 9052 13050 9064
rect 13218 9061 13230 9064
rect 13264 9061 13268 9095
rect 13218 9055 13268 9061
rect 13262 9052 13268 9055
rect 13320 9052 13326 9104
rect 14550 9052 14556 9104
rect 14608 9092 14614 9104
rect 14918 9092 14924 9104
rect 14608 9064 14924 9092
rect 14608 9052 14614 9064
rect 14918 9052 14924 9064
rect 14976 9092 14982 9104
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 14976 9064 15485 9092
rect 14976 9052 14982 9064
rect 15473 9061 15485 9064
rect 15519 9092 15531 9095
rect 17037 9095 17095 9101
rect 17037 9092 17049 9095
rect 15519 9064 17049 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 17037 9061 17049 9064
rect 17083 9061 17095 9095
rect 17037 9055 17095 9061
rect 19886 9052 19892 9104
rect 19944 9092 19950 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 19944 9064 21097 9092
rect 19944 9052 19950 9064
rect 21085 9061 21097 9064
rect 21131 9092 21143 9095
rect 21726 9092 21732 9104
rect 21131 9064 21732 9092
rect 21131 9061 21143 9064
rect 21085 9055 21143 9061
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 106 8984 112 9036
rect 164 9024 170 9036
rect 1464 9027 1522 9033
rect 1464 9024 1476 9027
rect 164 8996 1476 9024
rect 164 8984 170 8996
rect 1464 8993 1476 8996
rect 1510 9024 1522 9027
rect 1762 9024 1768 9036
rect 1510 8996 1768 9024
rect 1510 8993 1522 8996
rect 1464 8987 1522 8993
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 2869 9027 2927 9033
rect 2869 8993 2881 9027
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 2498 8916 2504 8968
rect 2556 8956 2562 8968
rect 2884 8956 2912 8987
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 3421 9027 3479 9033
rect 3421 9024 3433 9027
rect 3200 8996 3433 9024
rect 3200 8984 3206 8996
rect 3421 8993 3433 8996
rect 3467 8993 3479 9027
rect 6086 9024 6092 9036
rect 6047 8996 6092 9024
rect 3421 8987 3479 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8570 9024 8576 9036
rect 8531 8996 8576 9024
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11514 9024 11520 9036
rect 11471 8996 11520 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 17586 8984 17592 9036
rect 17644 9024 17650 9036
rect 18414 9024 18420 9036
rect 17644 8996 18420 9024
rect 17644 8984 17650 8996
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 18932 8996 18977 9024
rect 18932 8984 18938 8996
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 22500 9027 22558 9033
rect 22500 9024 22512 9027
rect 21876 8996 22512 9024
rect 21876 8984 21882 8996
rect 22500 8993 22512 8996
rect 22546 9024 22558 9027
rect 23106 9024 23112 9036
rect 22546 8996 23112 9024
rect 22546 8993 22558 8996
rect 22500 8987 22558 8993
rect 23106 8984 23112 8996
rect 23164 9024 23170 9036
rect 23512 9027 23570 9033
rect 23512 9024 23524 9027
rect 23164 8996 23524 9024
rect 23164 8984 23170 8996
rect 23512 8993 23524 8996
rect 23558 8993 23570 9027
rect 23512 8987 23570 8993
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2556 8928 3801 8956
rect 2556 8916 2562 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 3936 8928 4629 8956
rect 3936 8916 3942 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 7282 8956 7288 8968
rect 5307 8928 7288 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 1535 8891 1593 8897
rect 1535 8857 1547 8891
rect 1581 8888 1593 8891
rect 2958 8888 2964 8900
rect 1581 8860 2964 8888
rect 1581 8857 1593 8860
rect 1535 8851 1593 8857
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 3694 8848 3700 8900
rect 3752 8888 3758 8900
rect 5276 8888 5304 8919
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9398 8956 9404 8968
rect 8803 8928 9404 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 11054 8956 11060 8968
rect 9723 8928 11060 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12894 8956 12900 8968
rect 12855 8928 12900 8956
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15427 8928 16896 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 3752 8860 5304 8888
rect 3752 8848 3758 8860
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 15194 8888 15200 8900
rect 12032 8860 15200 8888
rect 12032 8848 12038 8860
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 15286 8848 15292 8900
rect 15344 8888 15350 8900
rect 15396 8888 15424 8919
rect 15930 8888 15936 8900
rect 15344 8860 15424 8888
rect 15891 8860 15936 8888
rect 15344 8848 15350 8860
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 16868 8888 16896 8928
rect 16942 8916 16948 8968
rect 17000 8956 17006 8968
rect 17218 8956 17224 8968
rect 17000 8928 17045 8956
rect 17179 8928 17224 8956
rect 17000 8916 17006 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17678 8916 17684 8968
rect 17736 8956 17742 8968
rect 17865 8959 17923 8965
rect 17865 8956 17877 8959
rect 17736 8928 17877 8956
rect 17736 8916 17742 8928
rect 17865 8925 17877 8928
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18966 8916 18972 8968
rect 19024 8956 19030 8968
rect 19153 8959 19211 8965
rect 19153 8956 19165 8959
rect 19024 8928 19165 8956
rect 19024 8916 19030 8928
rect 19153 8925 19165 8928
rect 19199 8956 19211 8959
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19199 8928 19441 8956
rect 19199 8925 19211 8928
rect 19153 8919 19211 8925
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 20254 8916 20260 8968
rect 20312 8956 20318 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20312 8928 21005 8956
rect 20312 8916 20318 8928
rect 20993 8925 21005 8928
rect 21039 8956 21051 8959
rect 22603 8959 22661 8965
rect 22603 8956 22615 8959
rect 21039 8928 22615 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 22603 8925 22615 8928
rect 22649 8925 22661 8959
rect 22603 8919 22661 8925
rect 16868 8860 18000 8888
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2038 8820 2044 8832
rect 1995 8792 2044 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 2314 8820 2320 8832
rect 2275 8792 2320 8820
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 4890 8780 4896 8832
rect 4948 8820 4954 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 4948 8792 5549 8820
rect 4948 8780 4954 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 7742 8820 7748 8832
rect 7703 8792 7748 8820
rect 5537 8783 5595 8789
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10008 8792 10885 8820
rect 10008 8780 10014 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 10873 8783 10931 8789
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 14826 8820 14832 8832
rect 14787 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16574 8820 16580 8832
rect 16531 8792 16580 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16574 8780 16580 8792
rect 16632 8820 16638 8832
rect 17678 8820 17684 8832
rect 16632 8792 17684 8820
rect 16632 8780 16638 8792
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 17972 8820 18000 8860
rect 18230 8848 18236 8900
rect 18288 8888 18294 8900
rect 21174 8888 21180 8900
rect 18288 8860 21180 8888
rect 18288 8848 18294 8860
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 21266 8848 21272 8900
rect 21324 8888 21330 8900
rect 21545 8891 21603 8897
rect 21545 8888 21557 8891
rect 21324 8860 21557 8888
rect 21324 8848 21330 8860
rect 21545 8857 21557 8860
rect 21591 8857 21603 8891
rect 21545 8851 21603 8857
rect 23615 8823 23673 8829
rect 23615 8820 23627 8823
rect 17972 8792 23627 8820
rect 23615 8789 23627 8792
rect 23661 8789 23673 8823
rect 23615 8783 23673 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2222 8616 2228 8628
rect 2183 8588 2228 8616
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3326 8616 3332 8628
rect 2915 8588 3332 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 4764 8588 5825 8616
rect 4764 8576 4770 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 5813 8579 5871 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 9858 8616 9864 8628
rect 9815 8588 9864 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 9858 8576 9864 8588
rect 9916 8616 9922 8628
rect 11054 8616 11060 8628
rect 9916 8588 10916 8616
rect 11015 8588 11060 8616
rect 9916 8576 9922 8588
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1857 8551 1915 8557
rect 1857 8548 1869 8551
rect 1636 8520 1869 8548
rect 1636 8508 1642 8520
rect 1857 8517 1869 8520
rect 1903 8548 1915 8551
rect 2593 8551 2651 8557
rect 2593 8548 2605 8551
rect 1903 8520 2605 8548
rect 1903 8517 1915 8520
rect 1857 8511 1915 8517
rect 2593 8517 2605 8520
rect 2639 8517 2651 8551
rect 7558 8548 7564 8560
rect 7471 8520 7564 8548
rect 2593 8511 2651 8517
rect 7558 8508 7564 8520
rect 7616 8548 7622 8560
rect 10686 8548 10692 8560
rect 7616 8520 10692 8548
rect 7616 8508 7622 8520
rect 10686 8508 10692 8520
rect 10744 8508 10750 8560
rect 10888 8548 10916 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14550 8616 14556 8628
rect 14323 8588 14556 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14550 8576 14556 8588
rect 14608 8616 14614 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 14608 8588 16129 8616
rect 14608 8576 14614 8588
rect 16117 8585 16129 8588
rect 16163 8616 16175 8619
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 16163 8588 16497 8616
rect 16163 8585 16175 8588
rect 16117 8579 16175 8585
rect 16485 8585 16497 8588
rect 16531 8585 16543 8619
rect 17770 8616 17776 8628
rect 17731 8588 17776 8616
rect 16485 8579 16543 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18414 8616 18420 8628
rect 18375 8588 18420 8616
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 19886 8616 19892 8628
rect 19847 8588 19892 8616
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 21726 8616 21732 8628
rect 21687 8588 21732 8616
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 23106 8616 23112 8628
rect 23067 8588 23112 8616
rect 23106 8576 23112 8588
rect 23164 8616 23170 8628
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 23164 8588 23857 8616
rect 23164 8576 23170 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 12897 8551 12955 8557
rect 12897 8548 12909 8551
rect 10888 8520 12909 8548
rect 12897 8517 12909 8520
rect 12943 8548 12955 8551
rect 12986 8548 12992 8560
rect 12943 8520 12992 8548
rect 12943 8517 12955 8520
rect 12897 8511 12955 8517
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 14642 8548 14648 8560
rect 13786 8520 14648 8548
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2038 8480 2044 8492
rect 1995 8452 2044 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2958 8440 2964 8492
rect 3016 8480 3022 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 3016 8452 3249 8480
rect 3016 8440 3022 8452
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3237 8443 3295 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8480 7067 8483
rect 7742 8480 7748 8492
rect 7055 8452 7748 8480
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 12618 8480 12624 8492
rect 8496 8452 12624 8480
rect 1728 8415 1786 8421
rect 1728 8381 1740 8415
rect 1774 8412 1786 8415
rect 2314 8412 2320 8424
rect 1774 8384 2320 8412
rect 1774 8381 1786 8384
rect 1728 8375 1786 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 8496 8421 8524 8452
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8480 13415 8483
rect 13786 8480 13814 8520
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 16807 8551 16865 8557
rect 16807 8517 16819 8551
rect 16853 8548 16865 8551
rect 21450 8548 21456 8560
rect 16853 8520 21456 8548
rect 16853 8517 16865 8520
rect 16807 8511 16865 8517
rect 21450 8508 21456 8520
rect 21508 8508 21514 8560
rect 13403 8452 13814 8480
rect 15013 8483 15071 8489
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 15197 8483 15255 8489
rect 15197 8480 15209 8483
rect 15059 8452 15209 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15197 8449 15209 8452
rect 15243 8480 15255 8483
rect 18046 8480 18052 8492
rect 15243 8452 18052 8480
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18966 8480 18972 8492
rect 18927 8452 18972 8480
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 21634 8480 21640 8492
rect 20855 8452 21640 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 8481 8415 8539 8421
rect 8481 8412 8493 8415
rect 8312 8384 8493 8412
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 1581 8347 1639 8353
rect 1581 8344 1593 8347
rect 1544 8316 1593 8344
rect 1544 8304 1550 8316
rect 1581 8313 1593 8316
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 1596 8276 1624 8307
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 3329 8347 3387 8353
rect 2740 8316 3261 8344
rect 2740 8304 2746 8316
rect 2869 8279 2927 8285
rect 2869 8276 2881 8279
rect 1596 8248 2881 8276
rect 2869 8245 2881 8248
rect 2915 8276 2927 8279
rect 2961 8279 3019 8285
rect 2961 8276 2973 8279
rect 2915 8248 2973 8276
rect 2915 8245 2927 8248
rect 2869 8239 2927 8245
rect 2961 8245 2973 8248
rect 3007 8245 3019 8279
rect 3233 8276 3261 8316
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 3418 8344 3424 8356
rect 3375 8316 3424 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 5255 8347 5313 8353
rect 5255 8313 5267 8347
rect 5301 8313 5313 8347
rect 5255 8307 5313 8313
rect 4246 8276 4252 8288
rect 3233 8248 4252 8276
rect 2961 8239 3019 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4798 8276 4804 8288
rect 4711 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8276 4862 8288
rect 5270 8276 5298 8307
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6641 8347 6699 8353
rect 5500 8316 6453 8344
rect 5500 8304 5506 8316
rect 5350 8276 5356 8288
rect 4856 8248 5356 8276
rect 4856 8236 4862 8248
rect 5350 8236 5356 8248
rect 5408 8276 5414 8288
rect 6089 8279 6147 8285
rect 6089 8276 6101 8279
rect 5408 8248 6101 8276
rect 5408 8236 5414 8248
rect 6089 8245 6101 8248
rect 6135 8245 6147 8279
rect 6425 8276 6453 8316
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6730 8344 6736 8356
rect 6687 8316 6736 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6730 8304 6736 8316
rect 6788 8344 6794 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 6788 8316 7113 8344
rect 6788 8304 6794 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 7101 8307 7159 8313
rect 8312 8285 8340 8384
rect 8481 8381 8493 8384
rect 8527 8381 8539 8415
rect 8481 8375 8539 8381
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8628 8384 8953 8412
rect 8628 8372 8634 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 16704 8415 16762 8421
rect 16704 8381 16716 8415
rect 16750 8381 16762 8415
rect 16704 8375 16762 8381
rect 9214 8344 9220 8356
rect 9175 8316 9220 8344
rect 9214 8304 9220 8316
rect 9272 8304 9278 8356
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10137 8347 10195 8353
rect 10137 8344 10149 8347
rect 10008 8316 10149 8344
rect 10008 8304 10014 8316
rect 10137 8313 10149 8316
rect 10183 8313 10195 8347
rect 10137 8307 10195 8313
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10284 8316 10329 8344
rect 10284 8304 10290 8316
rect 12986 8304 12992 8356
rect 13044 8344 13050 8356
rect 13678 8347 13736 8353
rect 13678 8344 13690 8347
rect 13044 8316 13690 8344
rect 13044 8304 13050 8316
rect 13678 8313 13690 8316
rect 13724 8313 13736 8347
rect 13678 8307 13736 8313
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 15289 8347 15347 8353
rect 15289 8344 15301 8347
rect 14240 8316 15301 8344
rect 14240 8304 14246 8316
rect 15289 8313 15301 8316
rect 15335 8344 15347 8347
rect 15378 8344 15384 8356
rect 15335 8316 15384 8344
rect 15335 8313 15347 8316
rect 15289 8307 15347 8313
rect 15378 8304 15384 8316
rect 15436 8304 15442 8356
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8344 15899 8347
rect 15930 8344 15936 8356
rect 15887 8316 15936 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 15930 8304 15936 8316
rect 15988 8304 15994 8356
rect 8297 8279 8355 8285
rect 8297 8276 8309 8279
rect 6425 8248 8309 8276
rect 6089 8239 6147 8245
rect 8297 8245 8309 8248
rect 8343 8245 8355 8279
rect 11514 8276 11520 8288
rect 11475 8248 11520 8276
rect 8297 8239 8355 8245
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 15654 8276 15660 8288
rect 13136 8248 15660 8276
rect 13136 8236 13142 8248
rect 15654 8236 15660 8248
rect 15712 8276 15718 8288
rect 16719 8276 16747 8375
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22316 8415 22374 8421
rect 22316 8412 22328 8415
rect 22060 8384 22328 8412
rect 22060 8372 22066 8384
rect 22316 8381 22328 8384
rect 22362 8412 22374 8415
rect 22741 8415 22799 8421
rect 22741 8412 22753 8415
rect 22362 8384 22753 8412
rect 22362 8381 22374 8384
rect 22316 8375 22374 8381
rect 22741 8381 22753 8384
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 18785 8347 18843 8353
rect 18785 8344 18797 8347
rect 17368 8316 18797 8344
rect 17368 8304 17374 8316
rect 18785 8313 18797 8316
rect 18831 8344 18843 8347
rect 19150 8344 19156 8356
rect 18831 8316 19156 8344
rect 18831 8313 18843 8316
rect 18785 8307 18843 8313
rect 19150 8304 19156 8316
rect 19208 8344 19214 8356
rect 19290 8347 19348 8353
rect 19290 8344 19302 8347
rect 19208 8316 19302 8344
rect 19208 8304 19214 8316
rect 19290 8313 19302 8316
rect 19336 8313 19348 8347
rect 19290 8307 19348 8313
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 20956 8316 21001 8344
rect 20956 8304 20962 8316
rect 21174 8304 21180 8356
rect 21232 8344 21238 8356
rect 21453 8347 21511 8353
rect 21453 8344 21465 8347
rect 21232 8316 21465 8344
rect 21232 8304 21238 8316
rect 21453 8313 21465 8316
rect 21499 8313 21511 8347
rect 21453 8307 21511 8313
rect 17129 8279 17187 8285
rect 17129 8276 17141 8279
rect 15712 8248 17141 8276
rect 15712 8236 15718 8248
rect 17129 8245 17141 8248
rect 17175 8245 17187 8279
rect 17129 8239 17187 8245
rect 20625 8279 20683 8285
rect 20625 8245 20637 8279
rect 20671 8276 20683 8279
rect 20916 8276 20944 8304
rect 20671 8248 20944 8276
rect 20671 8245 20683 8248
rect 20625 8239 20683 8245
rect 21634 8236 21640 8288
rect 21692 8276 21698 8288
rect 22094 8276 22100 8288
rect 21692 8248 22100 8276
rect 21692 8236 21698 8248
rect 22094 8236 22100 8248
rect 22152 8236 22158 8288
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 22419 8279 22477 8285
rect 22419 8276 22431 8279
rect 22244 8248 22431 8276
rect 22244 8236 22250 8248
rect 22419 8245 22431 8248
rect 22465 8245 22477 8279
rect 22419 8239 22477 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1728 8044 1961 8072
rect 1728 8032 1734 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3476 8044 3801 8072
rect 3476 8032 3482 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4614 8072 4620 8084
rect 4479 8044 4620 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 6086 8072 6092 8084
rect 6047 8044 6092 8072
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8251 8075 8309 8081
rect 8251 8072 8263 8075
rect 7800 8044 8263 8072
rect 7800 8032 7806 8044
rect 8251 8041 8263 8044
rect 8297 8041 8309 8075
rect 8570 8072 8576 8084
rect 8531 8044 8576 8072
rect 8251 8035 8309 8041
rect 8570 8032 8576 8044
rect 8628 8072 8634 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8628 8044 8953 8072
rect 8628 8032 8634 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 10134 8072 10140 8084
rect 10095 8044 10140 8072
rect 8941 8035 8999 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10244 8044 10609 8072
rect 106 7964 112 8016
rect 164 8004 170 8016
rect 3970 8004 3976 8016
rect 164 7976 3976 8004
rect 164 7964 170 7976
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 5163 8007 5221 8013
rect 5163 7973 5175 8007
rect 5209 8004 5221 8007
rect 5350 8004 5356 8016
rect 5209 7976 5356 8004
rect 5209 7973 5221 7976
rect 5163 7967 5221 7973
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 6730 8004 6736 8016
rect 5736 7976 6736 8004
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 5736 7945 5764 7976
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 10244 8004 10272 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 12069 8075 12127 8081
rect 12069 8072 12081 8075
rect 11112 8044 12081 8072
rect 11112 8032 11118 8044
rect 12069 8041 12081 8044
rect 12115 8041 12127 8075
rect 12069 8035 12127 8041
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12952 8044 13001 8072
rect 12952 8032 12958 8044
rect 12989 8041 13001 8044
rect 13035 8072 13047 8075
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13035 8044 13645 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 15286 8072 15292 8084
rect 15151 8044 15292 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15473 8075 15531 8081
rect 15473 8072 15485 8075
rect 15436 8044 15485 8072
rect 15436 8032 15442 8044
rect 15473 8041 15485 8044
rect 15519 8041 15531 8075
rect 15473 8035 15531 8041
rect 15887 8075 15945 8081
rect 15887 8041 15899 8075
rect 15933 8072 15945 8075
rect 16482 8072 16488 8084
rect 15933 8044 16488 8072
rect 15933 8041 15945 8044
rect 15887 8035 15945 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8072 16727 8075
rect 16942 8072 16948 8084
rect 16715 8044 16948 8072
rect 16715 8041 16727 8044
rect 16669 8035 16727 8041
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17678 8072 17684 8084
rect 17639 8044 17684 8072
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 21450 8032 21456 8084
rect 21508 8072 21514 8084
rect 22830 8072 22836 8084
rect 21508 8044 22836 8072
rect 21508 8032 21514 8044
rect 22830 8032 22836 8044
rect 22888 8032 22894 8084
rect 10410 8004 10416 8016
rect 9916 7976 10416 8004
rect 9916 7964 9922 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 17082 8007 17140 8013
rect 17082 8004 17094 8007
rect 14200 7976 17094 8004
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 3421 7939 3479 7945
rect 3421 7936 3433 7939
rect 2915 7908 3433 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 3421 7905 3433 7908
rect 3467 7905 3479 7939
rect 3421 7899 3479 7905
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2884 7868 2912 7899
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8180 7939 8238 7945
rect 8180 7936 8192 7939
rect 7892 7908 8192 7936
rect 7892 7896 7898 7908
rect 8180 7905 8192 7908
rect 8226 7936 8238 7939
rect 9030 7936 9036 7948
rect 8226 7908 9036 7936
rect 8226 7905 8238 7908
rect 8180 7899 8238 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 9456 7908 10241 7936
rect 9456 7896 9462 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 11974 7936 11980 7948
rect 11935 7908 11980 7936
rect 10229 7899 10287 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 12124 7908 12449 7936
rect 12124 7896 12130 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 12676 7908 13553 7936
rect 12676 7896 12682 7908
rect 13541 7905 13553 7908
rect 13587 7936 13599 7939
rect 13630 7936 13636 7948
rect 13587 7908 13636 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14090 7936 14096 7948
rect 14051 7908 14096 7936
rect 14090 7896 14096 7908
rect 14148 7896 14154 7948
rect 2556 7840 2912 7868
rect 3145 7871 3203 7877
rect 2556 7828 2562 7840
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 4798 7868 4804 7880
rect 3191 7840 4804 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6236 7840 6653 7868
rect 6236 7828 6242 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7006 7868 7012 7880
rect 6963 7840 7012 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 6932 7800 6960 7831
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 12084 7868 12112 7896
rect 8536 7840 12112 7868
rect 8536 7828 8542 7840
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 13044 7840 13369 7868
rect 13044 7828 13050 7840
rect 13357 7837 13369 7840
rect 13403 7868 13415 7871
rect 14200 7868 14228 7976
rect 17082 7973 17094 7976
rect 17128 8004 17140 8007
rect 17310 8004 17316 8016
rect 17128 7976 17316 8004
rect 17128 7973 17140 7976
rect 17082 7967 17140 7973
rect 17310 7964 17316 7976
rect 17368 7964 17374 8016
rect 17770 7964 17776 8016
rect 17828 8004 17834 8016
rect 21082 8004 21088 8016
rect 17828 7976 19012 8004
rect 21043 7976 21088 8004
rect 17828 7964 17834 7976
rect 18984 7948 19012 7976
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 21174 7964 21180 8016
rect 21232 8004 21238 8016
rect 21637 8007 21695 8013
rect 21637 8004 21649 8007
rect 21232 7976 21649 8004
rect 21232 7964 21238 7976
rect 21637 7973 21649 7976
rect 21683 7973 21695 8007
rect 21637 7967 21695 7973
rect 15816 7939 15874 7945
rect 15816 7905 15828 7939
rect 15862 7936 15874 7939
rect 16298 7936 16304 7948
rect 15862 7908 16304 7936
rect 15862 7905 15874 7908
rect 15816 7899 15874 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 18414 7896 18420 7948
rect 18472 7936 18478 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 18472 7908 18521 7936
rect 18472 7896 18478 7908
rect 18509 7905 18521 7908
rect 18555 7905 18567 7939
rect 18966 7936 18972 7948
rect 18879 7908 18972 7936
rect 18509 7899 18567 7905
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 16758 7868 16764 7880
rect 13403 7840 14228 7868
rect 16719 7840 16764 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21266 7868 21272 7880
rect 21039 7840 21272 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 3936 7772 6960 7800
rect 3936 7760 3942 7772
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 1762 7732 1768 7744
rect 1719 7704 1768 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 7926 7732 7932 7744
rect 7887 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11606 7732 11612 7744
rect 11195 7704 11612 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 14458 7692 14464 7744
rect 14516 7732 14522 7744
rect 22002 7732 22008 7744
rect 14516 7704 22008 7732
rect 14516 7692 14522 7704
rect 22002 7692 22008 7704
rect 22060 7692 22066 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2958 7488 2964 7540
rect 3016 7528 3022 7540
rect 3421 7531 3479 7537
rect 3421 7528 3433 7531
rect 3016 7500 3433 7528
rect 3016 7488 3022 7500
rect 3421 7497 3433 7500
rect 3467 7497 3479 7531
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3421 7491 3479 7497
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 4856 7500 5733 7528
rect 4856 7488 4862 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7650 7528 7656 7540
rect 6840 7500 7656 7528
rect 1670 7460 1676 7472
rect 1596 7432 1676 7460
rect 1596 7392 1624 7432
rect 1670 7420 1676 7432
rect 1728 7420 1734 7472
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 2777 7463 2835 7469
rect 2777 7460 2789 7463
rect 2740 7432 2789 7460
rect 2740 7420 2746 7432
rect 2777 7429 2789 7432
rect 2823 7460 2835 7463
rect 4154 7460 4160 7472
rect 2823 7432 4160 7460
rect 2823 7429 2835 7432
rect 2777 7423 2835 7429
rect 4154 7420 4160 7432
rect 4212 7460 4218 7472
rect 6840 7460 6868 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9723 7531 9781 7537
rect 9723 7528 9735 7531
rect 9640 7500 9735 7528
rect 9640 7488 9646 7500
rect 9723 7497 9735 7500
rect 9769 7497 9781 7531
rect 10042 7528 10048 7540
rect 10003 7500 10048 7528
rect 9723 7491 9781 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 11514 7528 11520 7540
rect 10244 7500 11520 7528
rect 4212 7432 6868 7460
rect 6963 7463 7021 7469
rect 4212 7420 4218 7432
rect 6963 7429 6975 7463
rect 7009 7460 7021 7463
rect 9950 7460 9956 7472
rect 7009 7432 9956 7460
rect 7009 7429 7021 7432
rect 6963 7423 7021 7429
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 1504 7364 1624 7392
rect 2041 7395 2099 7401
rect 1504 7333 1532 7364
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2130 7392 2136 7404
rect 2087 7364 2136 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3050 7392 3056 7404
rect 3007 7364 3056 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 4890 7392 4896 7404
rect 4851 7364 4896 7392
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6907 7364 7389 7392
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7293 1547 7327
rect 1489 7287 1547 7293
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1636 7296 1685 7324
rect 1636 7284 1642 7296
rect 1673 7293 1685 7296
rect 1719 7324 1731 7327
rect 1854 7324 1860 7336
rect 1719 7296 1860 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1912 7296 2329 7324
rect 1912 7284 1918 7296
rect 2317 7293 2329 7296
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 4249 7327 4307 7333
rect 4249 7293 4261 7327
rect 4295 7324 4307 7327
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4295 7296 4537 7324
rect 4295 7293 4307 7296
rect 4249 7287 4307 7293
rect 4525 7293 4537 7296
rect 4571 7293 4583 7327
rect 4525 7287 4583 7293
rect 4540 7256 4568 7287
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 6907 7333 6935 7364
rect 7377 7361 7389 7364
rect 7423 7392 7435 7395
rect 10244 7392 10272 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 14001 7531 14059 7537
rect 11756 7500 13814 7528
rect 11756 7488 11762 7500
rect 10410 7460 10416 7472
rect 10371 7432 10416 7460
rect 10410 7420 10416 7432
rect 10468 7420 10474 7472
rect 11241 7463 11299 7469
rect 11241 7429 11253 7463
rect 11287 7460 11299 7463
rect 11422 7460 11428 7472
rect 11287 7432 11428 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 11422 7420 11428 7432
rect 11480 7460 11486 7472
rect 13081 7463 13139 7469
rect 13081 7460 13093 7463
rect 11480 7432 13093 7460
rect 11480 7420 11486 7432
rect 13081 7429 13093 7432
rect 13127 7429 13139 7463
rect 13630 7460 13636 7472
rect 13591 7432 13636 7460
rect 13081 7423 13139 7429
rect 13630 7420 13636 7432
rect 13688 7420 13694 7472
rect 7423 7364 10272 7392
rect 10689 7395 10747 7401
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 10689 7361 10701 7395
rect 10735 7392 10747 7395
rect 11146 7392 11152 7404
rect 10735 7364 11152 7392
rect 10735 7361 10747 7364
rect 10689 7355 10747 7361
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 12066 7392 12072 7404
rect 11747 7364 12072 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12802 7392 12808 7404
rect 12575 7364 12808 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13786 7392 13814 7500
rect 14001 7497 14013 7531
rect 14047 7528 14059 7531
rect 14090 7528 14096 7540
rect 14047 7500 14096 7528
rect 14047 7497 14059 7500
rect 14001 7491 14059 7497
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 14415 7531 14473 7537
rect 14415 7497 14427 7531
rect 14461 7528 14473 7531
rect 14734 7528 14740 7540
rect 14461 7500 14740 7528
rect 14461 7497 14473 7500
rect 14415 7491 14473 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15197 7531 15255 7537
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15378 7528 15384 7540
rect 15243 7500 15384 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15378 7488 15384 7500
rect 15436 7528 15442 7540
rect 15562 7528 15568 7540
rect 15436 7500 15568 7528
rect 15436 7488 15442 7500
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 16991 7531 17049 7537
rect 16991 7528 17003 7531
rect 15804 7500 17003 7528
rect 15804 7488 15810 7500
rect 16991 7497 17003 7500
rect 17037 7497 17049 7531
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 16991 7491 17049 7497
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 18966 7528 18972 7540
rect 18927 7500 18972 7528
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19208 7500 19257 7528
rect 19208 7488 19214 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 20349 7531 20407 7537
rect 20349 7497 20361 7531
rect 20395 7528 20407 7531
rect 21082 7528 21088 7540
rect 20395 7500 21088 7528
rect 20395 7497 20407 7500
rect 20349 7491 20407 7497
rect 21082 7488 21088 7500
rect 21140 7528 21146 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 21140 7500 22385 7528
rect 21140 7488 21146 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 22373 7491 22431 7497
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 15933 7463 15991 7469
rect 15933 7460 15945 7463
rect 15528 7432 15945 7460
rect 15528 7420 15534 7432
rect 15933 7429 15945 7432
rect 15979 7460 15991 7463
rect 16022 7460 16028 7472
rect 15979 7432 16028 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 20898 7420 20904 7472
rect 20956 7460 20962 7472
rect 22097 7463 22155 7469
rect 22097 7460 22109 7463
rect 20956 7432 22109 7460
rect 20956 7420 20962 7432
rect 22097 7429 22109 7432
rect 22143 7429 22155 7463
rect 22097 7423 22155 7429
rect 18046 7392 18052 7404
rect 13786 7364 16931 7392
rect 18007 7364 18052 7392
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4672 7296 4813 7324
rect 4672 7284 4678 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 6892 7327 6950 7333
rect 6892 7293 6904 7327
rect 6938 7293 6950 7327
rect 6892 7287 6950 7293
rect 9652 7327 9710 7333
rect 9652 7293 9664 7327
rect 9698 7324 9710 7327
rect 10042 7324 10048 7336
rect 9698 7296 10048 7324
rect 9698 7293 9710 7296
rect 9652 7287 9710 7293
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 14344 7327 14402 7333
rect 14344 7293 14356 7327
rect 14390 7324 14402 7327
rect 14458 7324 14464 7336
rect 14390 7296 14464 7324
rect 14390 7293 14402 7296
rect 14344 7287 14402 7293
rect 14458 7284 14464 7296
rect 14516 7324 14522 7336
rect 16903 7333 16931 7364
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 19300 7364 19441 7392
rect 19300 7352 19306 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 19429 7355 19487 7361
rect 19765 7364 21005 7392
rect 14737 7327 14795 7333
rect 14737 7324 14749 7327
rect 14516 7296 14749 7324
rect 14516 7284 14522 7296
rect 14737 7293 14749 7296
rect 14783 7293 14795 7327
rect 14737 7287 14795 7293
rect 16888 7327 16946 7333
rect 16888 7293 16900 7327
rect 16934 7324 16946 7327
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 16934 7296 17693 7324
rect 16934 7293 16946 7296
rect 16888 7287 16946 7293
rect 17681 7293 17693 7296
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 4982 7256 4988 7268
rect 4540 7228 4988 7256
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5994 7256 6000 7268
rect 5040 7228 6000 7256
rect 5040 7216 5046 7228
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 7926 7256 7932 7268
rect 7887 7228 7932 7256
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8021 7259 8079 7265
rect 8021 7225 8033 7259
rect 8067 7225 8079 7259
rect 8021 7219 8079 7225
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8662 7256 8668 7268
rect 8619 7228 8668 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 5350 7188 5356 7200
rect 5311 7160 5356 7188
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 7745 7191 7803 7197
rect 7745 7157 7757 7191
rect 7791 7188 7803 7191
rect 8036 7188 8064 7219
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 12618 7256 12624 7268
rect 10836 7228 10881 7256
rect 12579 7228 12624 7256
rect 10836 7216 10842 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 15378 7256 15384 7268
rect 15339 7228 15384 7256
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 15473 7259 15531 7265
rect 15473 7225 15485 7259
rect 15519 7256 15531 7259
rect 15562 7256 15568 7268
rect 15519 7228 15568 7256
rect 15519 7225 15531 7228
rect 15473 7219 15531 7225
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19765 7265 19793 7364
rect 20993 7361 21005 7364
rect 21039 7392 21051 7395
rect 21039 7364 21541 7392
rect 21039 7361 21051 7364
rect 20993 7355 21051 7361
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 20640 7296 21189 7324
rect 19750 7259 19808 7265
rect 19750 7256 19762 7259
rect 19208 7228 19762 7256
rect 19208 7216 19214 7228
rect 19750 7225 19762 7228
rect 19796 7225 19808 7259
rect 19750 7219 19808 7225
rect 20640 7200 20668 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 21513 7265 21541 7364
rect 21498 7259 21556 7265
rect 21498 7225 21510 7259
rect 21544 7225 21556 7259
rect 21498 7219 21556 7225
rect 8202 7188 8208 7200
rect 7791 7160 8208 7188
rect 7791 7157 7803 7160
rect 7745 7151 7803 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 8941 7191 8999 7197
rect 8941 7157 8953 7191
rect 8987 7188 8999 7191
rect 9030 7188 9036 7200
rect 8987 7160 9036 7188
rect 8987 7157 8999 7160
rect 8941 7151 8999 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 11974 7188 11980 7200
rect 11887 7160 11980 7188
rect 11974 7148 11980 7160
rect 12032 7188 12038 7200
rect 12434 7188 12440 7200
rect 12032 7160 12440 7188
rect 12032 7148 12038 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 16298 7188 16304 7200
rect 16259 7160 16304 7188
rect 16298 7148 16304 7160
rect 16356 7148 16362 7200
rect 16758 7188 16764 7200
rect 16719 7160 16764 7188
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 18414 7148 18420 7200
rect 18472 7188 18478 7200
rect 18509 7191 18567 7197
rect 18509 7188 18521 7191
rect 18472 7160 18521 7188
rect 18472 7148 18478 7160
rect 18509 7157 18521 7160
rect 18555 7157 18567 7191
rect 20622 7188 20628 7200
rect 20583 7160 20628 7188
rect 18509 7151 18567 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 1673 6987 1731 6993
rect 1673 6984 1685 6987
rect 1544 6956 1685 6984
rect 1544 6944 1550 6956
rect 1673 6953 1685 6956
rect 1719 6953 1731 6987
rect 2498 6984 2504 6996
rect 2459 6956 2504 6984
rect 1673 6947 1731 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 5859 6987 5917 6993
rect 5859 6953 5871 6987
rect 5905 6984 5917 6987
rect 6914 6984 6920 6996
rect 5905 6956 6920 6984
rect 5905 6953 5917 6956
rect 5859 6947 5917 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 8202 6984 8208 6996
rect 8163 6956 8208 6984
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10597 6987 10655 6993
rect 9916 6956 10041 6984
rect 9916 6944 9922 6956
rect 1397 6919 1455 6925
rect 1397 6885 1409 6919
rect 1443 6916 1455 6919
rect 1946 6916 1952 6928
rect 1443 6888 1952 6916
rect 1443 6885 1455 6888
rect 1397 6879 1455 6885
rect 1946 6876 1952 6888
rect 2004 6876 2010 6928
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 7647 6919 7705 6925
rect 2832 6888 6960 6916
rect 2832 6876 2838 6888
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 3028 6851 3086 6857
rect 3028 6817 3040 6851
rect 3074 6848 3086 6851
rect 3786 6848 3792 6860
rect 3074 6820 3792 6848
rect 3074 6817 3086 6820
rect 3028 6811 3086 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4246 6848 4252 6860
rect 4207 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4632 6857 4660 6888
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5788 6851 5846 6857
rect 5788 6848 5800 6851
rect 5592 6820 5800 6848
rect 5592 6808 5598 6820
rect 5788 6817 5800 6820
rect 5834 6848 5846 6851
rect 5902 6848 5908 6860
rect 5834 6820 5908 6848
rect 5834 6817 5846 6820
rect 5788 6811 5846 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6932 6857 6960 6888
rect 7647 6885 7659 6919
rect 7693 6916 7705 6919
rect 7834 6916 7840 6928
rect 7693 6888 7840 6916
rect 7693 6885 7705 6888
rect 7647 6879 7705 6885
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 10013 6925 10041 6956
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 10778 6984 10784 6996
rect 10643 6956 10784 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 10778 6944 10784 6956
rect 10836 6984 10842 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10836 6956 10885 6984
rect 10836 6944 10842 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 16945 6987 17003 6993
rect 16945 6984 16957 6987
rect 16816 6956 16957 6984
rect 16816 6944 16822 6956
rect 16945 6953 16957 6956
rect 16991 6953 17003 6987
rect 16945 6947 17003 6953
rect 19242 6944 19248 6996
rect 19300 6984 19306 6996
rect 19521 6987 19579 6993
rect 19521 6984 19533 6987
rect 19300 6956 19533 6984
rect 19300 6944 19306 6956
rect 19521 6953 19533 6956
rect 19567 6953 19579 6987
rect 19521 6947 19579 6953
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 21266 6984 21272 6996
rect 20763 6956 21272 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 9998 6919 10056 6925
rect 9998 6885 10010 6919
rect 10044 6885 10056 6919
rect 11606 6916 11612 6928
rect 11567 6888 11612 6916
rect 9998 6879 10056 6885
rect 11606 6876 11612 6888
rect 11664 6916 11670 6928
rect 12437 6919 12495 6925
rect 12437 6916 12449 6919
rect 11664 6888 12449 6916
rect 11664 6876 11670 6888
rect 12437 6885 12449 6888
rect 12483 6916 12495 6919
rect 12618 6916 12624 6928
rect 12483 6888 12624 6916
rect 12483 6885 12495 6888
rect 12437 6879 12495 6885
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 13538 6916 13544 6928
rect 13499 6888 13544 6916
rect 13538 6876 13544 6888
rect 13596 6876 13602 6928
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 15473 6919 15531 6925
rect 13872 6888 13917 6916
rect 13872 6876 13878 6888
rect 15473 6885 15485 6919
rect 15519 6916 15531 6919
rect 15562 6916 15568 6928
rect 15519 6888 15568 6916
rect 15519 6885 15531 6888
rect 15473 6879 15531 6885
rect 15562 6876 15568 6888
rect 15620 6876 15626 6928
rect 16022 6916 16028 6928
rect 15983 6888 16028 6916
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 20990 6876 20996 6928
rect 21048 6916 21054 6928
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 21048 6888 21097 6916
rect 21048 6876 21054 6888
rect 21085 6885 21097 6888
rect 21131 6916 21143 6919
rect 21726 6916 21732 6928
rect 21131 6888 21732 6916
rect 21131 6885 21143 6888
rect 21085 6879 21143 6885
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7190 6848 7196 6860
rect 6963 6820 7196 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 7190 6808 7196 6820
rect 7248 6848 7254 6860
rect 8570 6848 8576 6860
rect 7248 6820 8576 6848
rect 7248 6808 7254 6820
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9272 6820 9689 6848
rect 9272 6808 9278 6820
rect 9677 6817 9689 6820
rect 9723 6848 9735 6851
rect 9858 6848 9864 6860
rect 9723 6820 9864 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4396 6752 4813 6780
rect 4396 6740 4402 6752
rect 4801 6749 4813 6752
rect 4847 6780 4859 6783
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4847 6752 5089 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 7374 6780 7380 6792
rect 7331 6752 7380 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11974 6780 11980 6792
rect 11563 6752 11980 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 13556 6780 13584 6876
rect 17126 6848 17132 6860
rect 17087 6820 17132 6848
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17276 6820 17417 6848
rect 17276 6808 17282 6820
rect 17405 6817 17417 6820
rect 17451 6848 17463 6851
rect 17770 6848 17776 6860
rect 17451 6820 17776 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 18598 6848 18604 6860
rect 18559 6820 18604 6848
rect 18598 6808 18604 6820
rect 18656 6808 18662 6860
rect 18966 6848 18972 6860
rect 18927 6820 18972 6848
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 20622 6848 20628 6860
rect 19291 6820 20628 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 21692 6820 21737 6848
rect 21692 6808 21698 6820
rect 13722 6780 13728 6792
rect 13556 6752 13728 6780
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6780 15439 6783
rect 16390 6780 16396 6792
rect 15427 6752 16396 6780
rect 15427 6749 15439 6752
rect 15381 6743 15439 6749
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6780 21051 6783
rect 21358 6780 21364 6792
rect 21039 6752 21364 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21358 6740 21364 6752
rect 21416 6780 21422 6792
rect 22186 6780 22192 6792
rect 21416 6752 22192 6780
rect 21416 6740 21422 6752
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 3099 6715 3157 6721
rect 3099 6681 3111 6715
rect 3145 6712 3157 6715
rect 8757 6715 8815 6721
rect 8757 6712 8769 6715
rect 3145 6684 8769 6712
rect 3145 6681 3157 6684
rect 3099 6675 3157 6681
rect 8757 6681 8769 6684
rect 8803 6712 8815 6715
rect 8846 6712 8852 6724
rect 8803 6684 8852 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 12066 6712 12072 6724
rect 12027 6684 12072 6712
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 14277 6715 14335 6721
rect 14277 6681 14289 6715
rect 14323 6712 14335 6715
rect 15654 6712 15660 6724
rect 14323 6684 15660 6712
rect 14323 6681 14335 6684
rect 14277 6675 14335 6681
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 11204 6616 11253 6644
rect 11204 6604 11210 6616
rect 11241 6613 11253 6616
rect 11287 6613 11299 6647
rect 12802 6644 12808 6656
rect 12763 6616 12808 6644
rect 11241 6607 11299 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 15105 6647 15163 6653
rect 15105 6613 15117 6647
rect 15151 6644 15163 6647
rect 15378 6644 15384 6656
rect 15151 6616 15384 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 15378 6604 15384 6616
rect 15436 6644 15442 6656
rect 15838 6644 15844 6656
rect 15436 6616 15844 6644
rect 15436 6604 15442 6616
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2685 6443 2743 6449
rect 2685 6409 2697 6443
rect 2731 6440 2743 6443
rect 3142 6440 3148 6452
rect 2731 6412 3148 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2976 6245 3004 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 3786 6400 3792 6412
rect 3844 6440 3850 6452
rect 3844 6412 7598 6440
rect 3844 6400 3850 6412
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 5592 6344 5733 6372
rect 5592 6332 5598 6344
rect 5721 6341 5733 6344
rect 5767 6372 5779 6375
rect 7466 6372 7472 6384
rect 5767 6344 7472 6372
rect 5767 6341 5779 6344
rect 5721 6335 5779 6341
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7570 6304 7598 6412
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8260 6412 8585 6440
rect 8260 6400 8266 6412
rect 8573 6409 8585 6412
rect 8619 6440 8631 6443
rect 8938 6440 8944 6452
rect 8619 6412 8944 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10778 6440 10784 6452
rect 10459 6412 10784 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 11606 6440 11612 6452
rect 11567 6412 11612 6440
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13872 6412 13921 6440
rect 13872 6400 13878 6412
rect 13909 6409 13921 6412
rect 13955 6440 13967 6443
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13955 6412 14197 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14185 6403 14243 6409
rect 17126 6400 17132 6452
rect 17184 6440 17190 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17184 6412 17417 6440
rect 17184 6400 17190 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 19058 6400 19064 6452
rect 19116 6440 19122 6452
rect 19613 6443 19671 6449
rect 19613 6440 19625 6443
rect 19116 6412 19625 6440
rect 19116 6400 19122 6412
rect 19613 6409 19625 6412
rect 19659 6409 19671 6443
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 19613 6403 19671 6409
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21358 6440 21364 6452
rect 21319 6412 21364 6440
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8662 6372 8668 6384
rect 8168 6344 8668 6372
rect 8168 6332 8174 6344
rect 8662 6332 8668 6344
rect 8720 6372 8726 6384
rect 11149 6375 11207 6381
rect 11149 6372 11161 6375
rect 8720 6344 11161 6372
rect 8720 6332 8726 6344
rect 11149 6341 11161 6344
rect 11195 6372 11207 6375
rect 12066 6372 12072 6384
rect 11195 6344 12072 6372
rect 11195 6341 11207 6344
rect 11149 6335 11207 6341
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 16853 6375 16911 6381
rect 16853 6341 16865 6375
rect 16899 6372 16911 6375
rect 17218 6372 17224 6384
rect 16899 6344 17224 6372
rect 16899 6341 16911 6344
rect 16853 6335 16911 6341
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 17310 6332 17316 6384
rect 17368 6372 17374 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17368 6344 17693 6372
rect 17368 6332 17374 6344
rect 17681 6341 17693 6344
rect 17727 6372 17739 6375
rect 17773 6375 17831 6381
rect 17773 6372 17785 6375
rect 17727 6344 17785 6372
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 17773 6341 17785 6344
rect 17819 6341 17831 6375
rect 17773 6335 17831 6341
rect 18969 6375 19027 6381
rect 18969 6341 18981 6375
rect 19015 6372 19027 6375
rect 19978 6372 19984 6384
rect 19015 6344 19984 6372
rect 19015 6341 19027 6344
rect 18969 6335 19027 6341
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 8294 6304 8300 6316
rect 7570 6276 8300 6304
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8846 6304 8852 6316
rect 8807 6276 8852 6304
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6304 9551 6307
rect 11422 6304 11428 6316
rect 9539 6276 11428 6304
rect 9539 6273 9551 6276
rect 9493 6267 9551 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6304 17003 6307
rect 19518 6304 19524 6316
rect 16991 6276 19524 6304
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 19518 6264 19524 6276
rect 19576 6304 19582 6316
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19576 6276 19901 6304
rect 19576 6264 19582 6276
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6304 20591 6307
rect 21174 6304 21180 6316
rect 20579 6276 21180 6304
rect 20579 6273 20591 6276
rect 20533 6267 20591 6273
rect 21174 6264 21180 6276
rect 21232 6264 21238 6316
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6236 6699 6239
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6687 6208 7113 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 7101 6199 7159 6205
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3252 6100 3280 6199
rect 3510 6168 3516 6180
rect 3471 6140 3516 6168
rect 3510 6128 3516 6140
rect 3568 6128 3574 6180
rect 4662 6171 4720 6177
rect 4662 6168 4674 6171
rect 4172 6140 4674 6168
rect 4172 6112 4200 6140
rect 4662 6137 4674 6140
rect 4708 6168 4720 6171
rect 5350 6168 5356 6180
rect 4708 6140 5356 6168
rect 4708 6137 4720 6140
rect 4662 6131 4720 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 7116 6168 7144 6199
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7248 6208 7297 6236
rect 7248 6196 7254 6208
rect 7285 6205 7297 6208
rect 7331 6236 7343 6239
rect 7742 6236 7748 6248
rect 7331 6208 7748 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 12986 6236 12992 6248
rect 12947 6208 12992 6236
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 14734 6236 14740 6248
rect 14695 6208 14740 6236
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 18046 6236 18052 6248
rect 18007 6208 18052 6236
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 19245 6239 19303 6245
rect 19245 6236 19257 6239
rect 18656 6208 19257 6236
rect 18656 6196 18662 6208
rect 19245 6205 19257 6208
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 8018 6168 8024 6180
rect 7116 6140 8024 6168
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 8996 6140 9041 6168
rect 8996 6128 9002 6140
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10597 6171 10655 6177
rect 10597 6168 10609 6171
rect 10100 6140 10609 6168
rect 10100 6128 10106 6140
rect 10597 6137 10609 6140
rect 10643 6137 10655 6171
rect 10597 6131 10655 6137
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 10778 6168 10784 6180
rect 10735 6140 10784 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 13354 6177 13360 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 11486 6140 12817 6168
rect 4154 6100 4160 6112
rect 2832 6072 3280 6100
rect 4115 6072 4160 6100
rect 2832 6060 2838 6072
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 7834 6100 7840 6112
rect 7795 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 11486 6100 11514 6140
rect 12805 6137 12817 6140
rect 12851 6168 12863 6171
rect 13310 6171 13360 6177
rect 13310 6168 13322 6171
rect 12851 6140 13322 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 13310 6137 13322 6140
rect 13356 6137 13360 6171
rect 13310 6131 13360 6137
rect 13354 6128 13360 6131
rect 13412 6168 13418 6180
rect 14553 6171 14611 6177
rect 14553 6168 14565 6171
rect 13412 6140 14565 6168
rect 13412 6128 13418 6140
rect 14553 6137 14565 6140
rect 14599 6168 14611 6171
rect 15058 6171 15116 6177
rect 15058 6168 15070 6171
rect 14599 6140 15070 6168
rect 14599 6137 14611 6140
rect 14553 6131 14611 6137
rect 15058 6137 15070 6140
rect 15104 6137 15116 6171
rect 15058 6131 15116 6137
rect 17681 6171 17739 6177
rect 17681 6137 17693 6171
rect 17727 6168 17739 6171
rect 18370 6171 18428 6177
rect 18370 6168 18382 6171
rect 17727 6140 18382 6168
rect 17727 6137 17739 6140
rect 17681 6131 17739 6137
rect 18370 6137 18382 6140
rect 18416 6137 18428 6171
rect 18370 6131 18428 6137
rect 19978 6128 19984 6180
rect 20036 6168 20042 6180
rect 20036 6140 20081 6168
rect 20036 6128 20042 6140
rect 11974 6100 11980 6112
rect 9824 6072 11514 6100
rect 11935 6072 11980 6100
rect 9824 6060 9830 6072
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15620 6072 15669 6100
rect 15620 6060 15626 6072
rect 15657 6069 15669 6072
rect 15703 6100 15715 6103
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15703 6072 15945 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 15933 6063 15991 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2774 5896 2780 5908
rect 2735 5868 2780 5896
rect 2774 5856 2780 5868
rect 2832 5896 2838 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 2832 5868 3801 5896
rect 2832 5856 2838 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 3789 5859 3847 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 7374 5896 7380 5908
rect 7335 5868 7380 5896
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 9858 5896 9864 5908
rect 9819 5868 9864 5896
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 12207 5899 12265 5905
rect 12207 5896 12219 5899
rect 10928 5868 12219 5896
rect 10928 5856 10934 5868
rect 12207 5865 12219 5868
rect 12253 5865 12265 5899
rect 12207 5859 12265 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 14090 5896 14096 5908
rect 12676 5868 14096 5896
rect 12676 5856 12682 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 18104 5868 18153 5896
rect 18104 5856 18110 5868
rect 18141 5865 18153 5868
rect 18187 5896 18199 5899
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 18187 5868 18521 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19797 5899 19855 5905
rect 19797 5896 19809 5899
rect 19576 5868 19809 5896
rect 19576 5856 19582 5868
rect 19797 5865 19809 5868
rect 19843 5865 19855 5899
rect 19797 5859 19855 5865
rect 4154 5788 4160 5840
rect 4212 5828 4218 5840
rect 4846 5831 4904 5837
rect 4846 5828 4858 5831
rect 4212 5800 4858 5828
rect 4212 5788 4218 5800
rect 4846 5797 4858 5800
rect 4892 5797 4904 5831
rect 4846 5791 4904 5797
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 6362 5828 6368 5840
rect 5316 5800 6368 5828
rect 5316 5788 5322 5800
rect 6362 5788 6368 5800
rect 6420 5828 6426 5840
rect 6457 5831 6515 5837
rect 6457 5828 6469 5831
rect 6420 5800 6469 5828
rect 6420 5788 6426 5800
rect 6457 5797 6469 5800
rect 6503 5797 6515 5831
rect 8202 5828 8208 5840
rect 8163 5800 8208 5828
rect 6457 5791 6515 5797
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 10686 5828 10692 5840
rect 10647 5800 10692 5828
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 13770 5831 13828 5837
rect 13770 5828 13782 5831
rect 13412 5800 13782 5828
rect 13412 5788 13418 5800
rect 13770 5797 13782 5800
rect 13816 5797 13828 5831
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 13770 5791 13828 5797
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 17034 5828 17040 5840
rect 16995 5800 17040 5828
rect 17034 5788 17040 5800
rect 17092 5788 17098 5840
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 12069 5763 12127 5769
rect 3568 5732 4154 5760
rect 3568 5720 3574 5732
rect 4126 5692 4154 5732
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12158 5760 12164 5772
rect 12115 5732 12164 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 18380 5732 18429 5760
rect 18380 5720 18386 5732
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18966 5760 18972 5772
rect 18927 5732 18972 5760
rect 18417 5723 18475 5729
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 21174 5720 21180 5772
rect 21232 5760 21238 5772
rect 23544 5763 23602 5769
rect 23544 5760 23556 5763
rect 21232 5732 23556 5760
rect 21232 5720 21238 5732
rect 23544 5729 23556 5732
rect 23590 5760 23602 5763
rect 23842 5760 23848 5772
rect 23590 5732 23848 5760
rect 23590 5729 23602 5732
rect 23544 5723 23602 5729
rect 23842 5720 23848 5732
rect 23900 5720 23906 5772
rect 4522 5692 4528 5704
rect 4126 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6454 5692 6460 5704
rect 6411 5664 6460 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6638 5692 6644 5704
rect 6599 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 11422 5692 11428 5704
rect 10643 5664 11428 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 6656 5624 6684 5652
rect 8404 5624 8432 5655
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 13446 5692 13452 5704
rect 13407 5664 13452 5692
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 16942 5692 16948 5704
rect 16903 5664 16948 5692
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 11149 5627 11207 5633
rect 11149 5624 11161 5627
rect 6656 5596 11161 5624
rect 11149 5593 11161 5596
rect 11195 5624 11207 5627
rect 11238 5624 11244 5636
rect 11195 5596 11244 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 15396 5624 15424 5652
rect 15930 5624 15936 5636
rect 15396 5596 15936 5624
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 17236 5624 17264 5655
rect 15988 5596 17264 5624
rect 15988 5584 15994 5596
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 10100 5528 10333 5556
rect 10100 5516 10106 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 10321 5519 10379 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 23615 5559 23673 5565
rect 23615 5525 23627 5559
rect 23661 5556 23673 5559
rect 24210 5556 24216 5568
rect 23661 5528 24216 5556
rect 23661 5525 23673 5528
rect 23615 5519 23673 5525
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4522 5352 4528 5364
rect 4295 5324 4528 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7834 5352 7840 5364
rect 7747 5324 7840 5352
rect 7834 5312 7840 5324
rect 7892 5352 7898 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 7892 5324 9689 5352
rect 7892 5312 7898 5324
rect 5721 5287 5779 5293
rect 5721 5253 5733 5287
rect 5767 5284 5779 5287
rect 6638 5284 6644 5296
rect 5767 5256 6644 5284
rect 5767 5253 5779 5256
rect 5721 5247 5779 5253
rect 6638 5244 6644 5256
rect 6696 5244 6702 5296
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 5031 5188 5181 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5169 5185 5181 5188
rect 5215 5216 5227 5219
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 5215 5188 6837 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7484 5120 7941 5148
rect 5261 5083 5319 5089
rect 5261 5049 5273 5083
rect 5307 5080 5319 5083
rect 5442 5080 5448 5092
rect 5307 5052 5448 5080
rect 5307 5049 5319 5052
rect 5261 5043 5319 5049
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 7484 5024 7512 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 8266 5089 8294 5324
rect 9677 5321 9689 5324
rect 9723 5352 9735 5355
rect 9766 5352 9772 5364
rect 9723 5324 9772 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10686 5352 10692 5364
rect 10647 5324 10692 5352
rect 10686 5312 10692 5324
rect 10744 5352 10750 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10744 5324 10977 5352
rect 10744 5312 10750 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 11422 5352 11428 5364
rect 11383 5324 11428 5352
rect 10965 5315 11023 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13412 5324 13461 5352
rect 13412 5312 13418 5324
rect 13449 5321 13461 5324
rect 13495 5352 13507 5355
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13495 5324 13829 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 13817 5315 13875 5321
rect 9784 5216 9812 5312
rect 12986 5216 12992 5228
rect 9784 5188 10180 5216
rect 12947 5188 12992 5216
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9355 5120 9781 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9769 5117 9781 5120
rect 9815 5148 9827 5151
rect 9950 5148 9956 5160
rect 9815 5120 9956 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10152 5089 10180 5188
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 12434 5148 12440 5160
rect 12395 5120 12440 5148
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12676 5120 12909 5148
rect 12676 5108 12682 5120
rect 12897 5117 12909 5120
rect 12943 5148 12955 5151
rect 13538 5148 13544 5160
rect 12943 5120 13544 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 8251 5083 8309 5089
rect 8251 5049 8263 5083
rect 8297 5049 8309 5083
rect 8251 5043 8309 5049
rect 10131 5083 10189 5089
rect 10131 5049 10143 5083
rect 10177 5049 10189 5083
rect 13832 5080 13860 5315
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 14424 5324 15209 5352
rect 14424 5312 14430 5324
rect 15197 5321 15209 5324
rect 15243 5352 15255 5355
rect 15470 5352 15476 5364
rect 15243 5324 15476 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 15620 5324 16865 5352
rect 15620 5312 15626 5324
rect 16853 5321 16865 5324
rect 16899 5352 16911 5355
rect 17034 5352 17040 5364
rect 16899 5324 17040 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18380 5324 18429 5352
rect 18380 5312 18386 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 22370 5352 22376 5364
rect 19208 5324 22376 5352
rect 19208 5312 19214 5324
rect 22370 5312 22376 5324
rect 22428 5312 22434 5364
rect 23842 5352 23848 5364
rect 23803 5324 23848 5352
rect 23842 5312 23848 5324
rect 23900 5312 23906 5364
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 15654 5284 15660 5296
rect 14332 5256 15660 5284
rect 14332 5244 14338 5256
rect 15654 5244 15660 5256
rect 15712 5284 15718 5296
rect 15712 5256 16160 5284
rect 15712 5244 15718 5256
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5216 15899 5219
rect 16022 5216 16028 5228
rect 15887 5188 16028 5216
rect 15887 5185 15899 5188
rect 15841 5179 15899 5185
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16132 5225 16160 5256
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 17000 5188 17325 5216
rect 17000 5176 17006 5188
rect 17313 5185 17325 5188
rect 17359 5216 17371 5219
rect 18831 5219 18889 5225
rect 18831 5216 18843 5219
rect 17359 5188 18843 5216
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 18831 5185 18843 5188
rect 18877 5185 18889 5219
rect 18831 5179 18889 5185
rect 13998 5148 14004 5160
rect 13959 5120 14004 5148
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 14921 5151 14979 5157
rect 14921 5117 14933 5151
rect 14967 5148 14979 5151
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 14967 5120 15577 5148
rect 14967 5117 14979 5120
rect 14921 5111 14979 5117
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 18744 5151 18802 5157
rect 18744 5117 18756 5151
rect 18790 5148 18802 5151
rect 19150 5148 19156 5160
rect 18790 5120 19156 5148
rect 18790 5117 18802 5120
rect 18744 5111 18802 5117
rect 14322 5083 14380 5089
rect 14322 5080 14334 5083
rect 13832 5052 14334 5080
rect 10131 5043 10189 5049
rect 14322 5049 14334 5052
rect 14368 5049 14380 5083
rect 14322 5043 14380 5049
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 4154 5012 4160 5024
rect 2372 4984 4160 5012
rect 2372 4972 2378 4984
rect 4154 4972 4160 4984
rect 4212 5012 4218 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4212 4984 4537 5012
rect 4212 4972 4218 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 7466 5012 7472 5024
rect 7427 4984 7472 5012
rect 4525 4975 4583 4981
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 15580 5012 15608 5111
rect 19150 5108 19156 5120
rect 19208 5108 19214 5160
rect 24210 5108 24216 5160
rect 24268 5148 24274 5160
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 24268 5120 24593 5148
rect 24268 5108 24274 5120
rect 24581 5117 24593 5120
rect 24627 5148 24639 5151
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24627 5120 25145 5148
rect 24627 5117 24639 5120
rect 24581 5111 24639 5117
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 15933 5083 15991 5089
rect 15933 5049 15945 5083
rect 15979 5049 15991 5083
rect 15933 5043 15991 5049
rect 15948 5012 15976 5043
rect 19150 5012 19156 5024
rect 15580 4984 15976 5012
rect 19111 4984 19156 5012
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 24765 5015 24823 5021
rect 24765 4981 24777 5015
rect 24811 5012 24823 5015
rect 27338 5012 27344 5024
rect 24811 4984 27344 5012
rect 24811 4981 24823 4984
rect 24765 4975 24823 4981
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 5442 4808 5448 4820
rect 5215 4780 5448 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8202 4808 8208 4820
rect 8159 4780 8208 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8202 4768 8208 4780
rect 8260 4808 8266 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8260 4780 8401 4808
rect 8260 4768 8266 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8720 4780 8769 4808
rect 8720 4768 8726 4780
rect 8757 4777 8769 4780
rect 8803 4777 8815 4811
rect 8757 4771 8815 4777
rect 12207 4811 12265 4817
rect 12207 4777 12219 4811
rect 12253 4808 12265 4811
rect 12802 4808 12808 4820
rect 12253 4780 12808 4808
rect 12253 4777 12265 4780
rect 12207 4771 12265 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13170 4808 13176 4820
rect 13035 4780 13176 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13170 4768 13176 4780
rect 13228 4808 13234 4820
rect 13446 4808 13452 4820
rect 13228 4780 13452 4808
rect 13228 4768 13234 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13998 4808 14004 4820
rect 13832 4780 14004 4808
rect 7555 4743 7613 4749
rect 7555 4709 7567 4743
rect 7601 4740 7613 4743
rect 7834 4740 7840 4752
rect 7601 4712 7840 4740
rect 7601 4709 7613 4712
rect 7555 4703 7613 4709
rect 7834 4700 7840 4712
rect 7892 4740 7898 4752
rect 8018 4740 8024 4752
rect 7892 4712 8024 4740
rect 7892 4700 7898 4712
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 8846 4700 8852 4752
rect 8904 4740 8910 4752
rect 9490 4740 9496 4752
rect 8904 4712 9496 4740
rect 8904 4700 8910 4712
rect 9490 4700 9496 4712
rect 9548 4740 9554 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9548 4712 9873 4740
rect 9548 4700 9554 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 11422 4740 11428 4752
rect 10459 4712 11428 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 11422 4700 11428 4712
rect 11480 4700 11486 4752
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 13832 4749 13860 4780
rect 13998 4768 14004 4780
rect 14056 4808 14062 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 14056 4780 14105 4808
rect 14056 4768 14062 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15378 4808 15384 4820
rect 15151 4780 15384 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 16080 4780 16313 4808
rect 16080 4768 16086 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 16301 4771 16359 4777
rect 16390 4768 16396 4820
rect 16448 4808 16454 4820
rect 16991 4811 17049 4817
rect 16991 4808 17003 4811
rect 16448 4780 17003 4808
rect 16448 4768 16454 4780
rect 16991 4777 17003 4780
rect 17037 4777 17049 4811
rect 16991 4771 17049 4777
rect 18509 4811 18567 4817
rect 18509 4777 18521 4811
rect 18555 4808 18567 4811
rect 18966 4808 18972 4820
rect 18555 4780 18972 4808
rect 18555 4777 18567 4780
rect 18509 4771 18567 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 12529 4743 12587 4749
rect 12529 4740 12541 4743
rect 12492 4712 12541 4740
rect 12492 4700 12498 4712
rect 12529 4709 12541 4712
rect 12575 4709 12587 4743
rect 12529 4703 12587 4709
rect 13817 4743 13875 4749
rect 13817 4709 13829 4743
rect 13863 4709 13875 4743
rect 13817 4703 13875 4709
rect 15473 4743 15531 4749
rect 15473 4709 15485 4743
rect 15519 4740 15531 4743
rect 15562 4740 15568 4752
rect 15519 4712 15568 4740
rect 15519 4709 15531 4712
rect 15473 4703 15531 4709
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 4706 4681 4712 4684
rect 4684 4675 4712 4681
rect 4684 4672 4696 4675
rect 2924 4644 4696 4672
rect 2924 4632 2930 4644
rect 4684 4641 4696 4644
rect 4684 4635 4712 4641
rect 4706 4632 4712 4635
rect 4764 4632 4770 4684
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 5905 4635 5963 4641
rect 5920 4604 5948 4635
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 12158 4681 12164 4684
rect 12136 4675 12164 4681
rect 12136 4672 12148 4675
rect 12071 4644 12148 4672
rect 12136 4641 12148 4644
rect 12216 4672 12222 4684
rect 13078 4672 13084 4684
rect 12216 4644 13084 4672
rect 12136 4635 12164 4641
rect 12158 4632 12164 4635
rect 12216 4632 12222 4644
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4641 13415 4675
rect 13538 4672 13544 4684
rect 13499 4644 13544 4672
rect 13357 4635 13415 4641
rect 5994 4604 6000 4616
rect 5920 4576 6000 4604
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 7190 4604 7196 4616
rect 6411 4576 7196 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 10686 4604 10692 4616
rect 9815 4576 10692 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 13372 4604 13400 4635
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 16850 4672 16856 4684
rect 16811 4644 16856 4672
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 15378 4604 15384 4616
rect 13372 4576 13492 4604
rect 15339 4576 15384 4604
rect 4755 4539 4813 4545
rect 4755 4505 4767 4539
rect 4801 4536 4813 4539
rect 6454 4536 6460 4548
rect 4801 4508 6460 4536
rect 4801 4505 4813 4508
rect 4755 4499 4813 4505
rect 6454 4496 6460 4508
rect 6512 4536 6518 4548
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 6512 4508 6653 4536
rect 6512 4496 6518 4508
rect 6641 4505 6653 4508
rect 6687 4505 6699 4539
rect 6641 4499 6699 4505
rect 13464 4480 13492 4576
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 15672 4536 15700 4567
rect 13780 4508 15700 4536
rect 13780 4496 13786 4508
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 13262 4468 13268 4480
rect 6052 4440 13268 4468
rect 6052 4428 6058 4440
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 18598 4468 18604 4480
rect 13504 4440 18604 4468
rect 13504 4428 13510 4440
rect 18598 4428 18604 4440
rect 18656 4428 18662 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 6086 4264 6092 4276
rect 5999 4236 6092 4264
rect 6086 4224 6092 4236
rect 6144 4264 6150 4276
rect 6546 4264 6552 4276
rect 6144 4236 6552 4264
rect 6144 4224 6150 4236
rect 6546 4224 6552 4236
rect 6604 4264 6610 4276
rect 7834 4264 7840 4276
rect 6604 4236 7840 4264
rect 6604 4224 6610 4236
rect 7834 4224 7840 4236
rect 7892 4264 7898 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 7892 4236 9137 4264
rect 7892 4224 7898 4236
rect 9125 4233 9137 4236
rect 9171 4264 9183 4267
rect 9309 4267 9367 4273
rect 9309 4264 9321 4267
rect 9171 4236 9321 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9309 4233 9321 4236
rect 9355 4233 9367 4267
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 9309 4227 9367 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11238 4264 11244 4276
rect 11164 4236 11244 4264
rect 4706 4196 4712 4208
rect 4619 4168 4712 4196
rect 4706 4156 4712 4168
rect 4764 4196 4770 4208
rect 5534 4196 5540 4208
rect 4764 4168 5540 4196
rect 4764 4156 4770 4168
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 5721 4199 5779 4205
rect 5721 4165 5733 4199
rect 5767 4196 5779 4199
rect 5994 4196 6000 4208
rect 5767 4168 6000 4196
rect 5767 4165 5779 4168
rect 5721 4159 5779 4165
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 7745 4199 7803 4205
rect 7745 4165 7757 4199
rect 7791 4196 7803 4199
rect 8018 4196 8024 4208
rect 7791 4168 8024 4196
rect 7791 4165 7803 4168
rect 7745 4159 7803 4165
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 8662 4156 8668 4208
rect 8720 4196 8726 4208
rect 8757 4199 8815 4205
rect 8757 4196 8769 4199
rect 8720 4168 8769 4196
rect 8720 4156 8726 4168
rect 8757 4165 8769 4168
rect 8803 4165 8815 4199
rect 8757 4159 8815 4165
rect 9784 4100 10594 4128
rect 6984 4063 7042 4069
rect 6984 4029 6996 4063
rect 7030 4060 7042 4063
rect 7374 4060 7380 4072
rect 7030 4032 7380 4060
rect 7030 4029 7042 4032
rect 6984 4023 7042 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 9490 4060 9496 4072
rect 9232 4032 9496 4060
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 8202 3992 8208 4004
rect 7239 3964 8208 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 9232 3992 9260 4032
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9784 4069 9812 4100
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9631 4032 9781 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9769 4023 9827 4029
rect 9876 4032 10149 4060
rect 8352 3964 9260 3992
rect 9309 3995 9367 4001
rect 8352 3952 8358 3964
rect 9309 3961 9321 3995
rect 9355 3992 9367 3995
rect 9876 3992 9904 4032
rect 10137 4029 10149 4032
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 9355 3964 9904 3992
rect 10566 3992 10594 4100
rect 11164 4060 11192 4236
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 12158 4264 12164 4276
rect 12119 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12897 4267 12955 4273
rect 12897 4264 12909 4267
rect 12299 4236 12909 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12897 4233 12909 4236
rect 12943 4264 12955 4267
rect 13446 4264 13452 4276
rect 12943 4236 13452 4264
rect 12943 4233 12955 4236
rect 12897 4227 12955 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 14369 4267 14427 4273
rect 14369 4264 14381 4267
rect 13596 4236 14381 4264
rect 13596 4224 13602 4236
rect 14369 4233 14381 4236
rect 14415 4233 14427 4267
rect 14369 4227 14427 4233
rect 14691 4267 14749 4273
rect 14691 4233 14703 4267
rect 14737 4264 14749 4267
rect 14826 4264 14832 4276
rect 14737 4236 14832 4264
rect 14737 4233 14749 4236
rect 14691 4227 14749 4233
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15703 4267 15761 4273
rect 15703 4264 15715 4267
rect 15528 4236 15715 4264
rect 15528 4224 15534 4236
rect 15703 4233 15715 4236
rect 15749 4233 15761 4267
rect 15703 4227 15761 4233
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 16715 4267 16773 4273
rect 16715 4264 16727 4267
rect 15896 4236 16727 4264
rect 15896 4224 15902 4236
rect 16715 4233 16727 4236
rect 16761 4233 16773 4267
rect 16715 4227 16773 4233
rect 14550 4156 14556 4208
rect 14608 4196 14614 4208
rect 15381 4199 15439 4205
rect 14608 4168 15148 4196
rect 14608 4156 14614 4168
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 14734 4128 14740 4140
rect 13771 4100 14740 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 11368 4063 11426 4069
rect 11368 4060 11380 4063
rect 11164 4032 11380 4060
rect 11368 4029 11380 4032
rect 11414 4029 11426 4063
rect 11368 4023 11426 4029
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 11572 4032 13001 4060
rect 11572 4020 11578 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 12989 4023 13047 4029
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14588 4063 14646 4069
rect 14588 4060 14600 4063
rect 14516 4032 14600 4060
rect 14516 4020 14522 4032
rect 14588 4029 14600 4032
rect 14634 4060 14646 4063
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14634 4032 15025 4060
rect 14634 4029 14646 4032
rect 14588 4023 14646 4029
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15120 4060 15148 4168
rect 15381 4165 15393 4199
rect 15427 4196 15439 4199
rect 15562 4196 15568 4208
rect 15427 4168 15568 4196
rect 15427 4165 15439 4168
rect 15381 4159 15439 4165
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 16114 4128 16120 4140
rect 16075 4100 16120 4128
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20714 4128 20720 4140
rect 19208 4100 20720 4128
rect 19208 4088 19214 4100
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 15632 4063 15690 4069
rect 15632 4060 15644 4063
rect 15120 4032 15644 4060
rect 15013 4023 15071 4029
rect 15632 4029 15644 4032
rect 15678 4060 15690 4063
rect 16132 4060 16160 4088
rect 15678 4032 16160 4060
rect 16644 4063 16702 4069
rect 15678 4029 15690 4032
rect 15632 4023 15690 4029
rect 16644 4029 16656 4063
rect 16690 4060 16702 4063
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 16690 4032 17509 4060
rect 16690 4029 16702 4032
rect 16644 4023 16702 4029
rect 17497 4029 17509 4032
rect 17543 4060 17555 4063
rect 19058 4060 19064 4072
rect 17543 4032 19064 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 19058 4020 19064 4032
rect 19116 4060 19122 4072
rect 22002 4060 22008 4072
rect 19116 4032 22008 4060
rect 19116 4020 19122 4032
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 12253 3995 12311 4001
rect 12253 3992 12265 3995
rect 10566 3964 12265 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 12253 3961 12265 3964
rect 12299 3961 12311 3995
rect 12253 3955 12311 3961
rect 14093 3995 14151 4001
rect 14093 3961 14105 3995
rect 14139 3992 14151 3995
rect 17310 3992 17316 4004
rect 14139 3964 17316 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 9950 3924 9956 3936
rect 9911 3896 9956 3924
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 11471 3927 11529 3933
rect 11471 3893 11483 3927
rect 11517 3924 11529 3927
rect 12618 3924 12624 3936
rect 11517 3896 12624 3924
rect 11517 3893 11529 3896
rect 11471 3887 11529 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 16850 3924 16856 3936
rect 16763 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3924 16914 3936
rect 17037 3927 17095 3933
rect 17037 3924 17049 3927
rect 16908 3896 17049 3924
rect 16908 3884 16914 3896
rect 17037 3893 17049 3896
rect 17083 3893 17095 3927
rect 17037 3887 17095 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7466 3720 7472 3732
rect 7427 3692 7472 3720
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8260 3692 8769 3720
rect 8260 3680 8266 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 8757 3683 8815 3689
rect 10367 3723 10425 3729
rect 10367 3689 10379 3723
rect 10413 3720 10425 3723
rect 10686 3720 10692 3732
rect 10413 3692 10692 3720
rect 10413 3689 10425 3692
rect 10367 3683 10425 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 13412 3692 13814 3720
rect 13412 3680 13418 3692
rect 8294 3612 8300 3664
rect 8352 3652 8358 3664
rect 8389 3655 8447 3661
rect 8389 3652 8401 3655
rect 8352 3624 8401 3652
rect 8352 3612 8358 3624
rect 8389 3621 8401 3624
rect 8435 3621 8447 3655
rect 8389 3615 8447 3621
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 9861 3655 9919 3661
rect 9861 3652 9873 3655
rect 9548 3624 9873 3652
rect 9548 3612 9554 3624
rect 9861 3621 9873 3624
rect 9907 3621 9919 3655
rect 9861 3615 9919 3621
rect 12989 3655 13047 3661
rect 12989 3621 13001 3655
rect 13035 3652 13047 3655
rect 13446 3652 13452 3664
rect 13035 3624 13452 3652
rect 13035 3621 13047 3624
rect 12989 3615 13047 3621
rect 13446 3612 13452 3624
rect 13504 3652 13510 3664
rect 13786 3652 13814 3692
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 15436 3692 15485 3720
rect 15436 3680 15442 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 19889 3723 19947 3729
rect 19889 3689 19901 3723
rect 19935 3720 19947 3723
rect 19978 3720 19984 3732
rect 19935 3692 19984 3720
rect 19935 3689 19947 3692
rect 19889 3683 19947 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 18414 3652 18420 3664
rect 13504 3624 13584 3652
rect 13786 3624 18420 3652
rect 13504 3612 13510 3624
rect 7650 3584 7656 3596
rect 7611 3556 7656 3584
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7800 3556 7849 3584
rect 7800 3544 7806 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 7837 3547 7895 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 13354 3584 13360 3596
rect 13315 3556 13360 3584
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 13556 3593 13584 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3584 13599 3587
rect 13906 3584 13912 3596
rect 13587 3556 13912 3584
rect 13587 3553 13599 3556
rect 13541 3547 13599 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 19702 3584 19708 3596
rect 16908 3556 19708 3584
rect 16908 3544 16914 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 10134 3380 10140 3392
rect 10095 3352 10140 3380
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 11422 3380 11428 3392
rect 11383 3352 11428 3380
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 6546 3176 6552 3188
rect 6507 3148 6552 3176
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7239 3179 7297 3185
rect 7239 3145 7251 3179
rect 7285 3176 7297 3179
rect 7926 3176 7932 3188
rect 7285 3148 7932 3176
rect 7285 3145 7297 3148
rect 7239 3139 7297 3145
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 10551 3179 10609 3185
rect 10551 3145 10563 3179
rect 10597 3176 10609 3179
rect 11146 3176 11152 3188
rect 10597 3148 11152 3176
rect 10597 3145 10609 3148
rect 10551 3139 10609 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12575 3179 12633 3185
rect 12575 3176 12587 3179
rect 12032 3148 12587 3176
rect 12032 3136 12038 3148
rect 12575 3145 12587 3148
rect 12621 3145 12633 3179
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 12575 3139 12633 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14274 3176 14280 3188
rect 14235 3148 14280 3176
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 19334 3176 19340 3188
rect 19295 3148 19340 3176
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19702 3176 19708 3188
rect 19663 3148 19708 3176
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 11333 3111 11391 3117
rect 11333 3108 11345 3111
rect 11296 3080 11345 3108
rect 11296 3068 11302 3080
rect 11333 3077 11345 3080
rect 11379 3108 11391 3111
rect 13587 3111 13645 3117
rect 13587 3108 13599 3111
rect 11379 3080 13599 3108
rect 11379 3077 11391 3080
rect 11333 3071 11391 3077
rect 13587 3077 13599 3080
rect 13633 3077 13645 3111
rect 13587 3071 13645 3077
rect 20073 3111 20131 3117
rect 20073 3077 20085 3111
rect 20119 3108 20131 3111
rect 22002 3108 22008 3120
rect 20119 3080 22008 3108
rect 20119 3077 20131 3080
rect 20073 3071 20131 3077
rect 22002 3068 22008 3080
rect 22060 3068 22066 3120
rect 24765 3111 24823 3117
rect 24765 3077 24777 3111
rect 24811 3108 24823 3111
rect 27614 3108 27620 3120
rect 24811 3080 27620 3108
rect 24811 3077 24823 3080
rect 24765 3071 24823 3077
rect 27614 3068 27620 3080
rect 27672 3068 27678 3120
rect 7650 3000 7656 3052
rect 7708 3040 7714 3052
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 7708 3012 7941 3040
rect 7708 3000 7714 3012
rect 7929 3009 7941 3012
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10321 3043 10379 3049
rect 10321 3040 10333 3043
rect 10192 3012 10333 3040
rect 10192 3000 10198 3012
rect 10321 3009 10333 3012
rect 10367 3040 10379 3043
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 10367 3012 13093 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 13081 3009 13093 3012
rect 13127 3009 13139 3043
rect 13722 3040 13728 3052
rect 13081 3003 13139 3009
rect 13372 3012 13728 3040
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 7136 2975 7194 2981
rect 7136 2972 7148 2975
rect 4028 2944 7148 2972
rect 4028 2932 4034 2944
rect 7136 2941 7148 2944
rect 7182 2972 7194 2975
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7182 2944 7573 2972
rect 7182 2941 7194 2944
rect 7136 2935 7194 2941
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 8205 2975 8263 2981
rect 8205 2941 8217 2975
rect 8251 2972 8263 2975
rect 8846 2972 8852 2984
rect 8251 2944 8852 2972
rect 8251 2941 8263 2944
rect 8205 2935 8263 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 10480 2975 10538 2981
rect 10480 2941 10492 2975
rect 10526 2972 10538 2975
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 10526 2944 10977 2972
rect 10526 2941 10538 2944
rect 10480 2935 10538 2941
rect 10965 2941 10977 2944
rect 11011 2972 11023 2975
rect 11698 2972 11704 2984
rect 11011 2944 11704 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 12360 2904 12388 2935
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12584 2944 12909 2972
rect 12584 2932 12590 2944
rect 12897 2941 12909 2944
rect 12943 2972 12955 2975
rect 13372 2972 13400 3012
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 12943 2944 13400 2972
rect 13516 2975 13574 2981
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13516 2941 13528 2975
rect 13562 2972 13574 2975
rect 14274 2972 14280 2984
rect 13562 2944 14280 2972
rect 13562 2941 13574 2944
rect 13516 2935 13574 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 18944 2975 19002 2981
rect 18944 2941 18956 2975
rect 18990 2972 19002 2975
rect 19334 2972 19340 2984
rect 18990 2944 19340 2972
rect 18990 2941 19002 2944
rect 18944 2935 19002 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 12544 2904 12572 2932
rect 12360 2876 12572 2904
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 19904 2904 19932 2935
rect 24026 2932 24032 2984
rect 24084 2972 24090 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24084 2944 24593 2972
rect 24084 2932 24090 2944
rect 24581 2941 24593 2944
rect 24627 2972 24639 2975
rect 25133 2975 25191 2981
rect 25133 2972 25145 2975
rect 24627 2944 25145 2972
rect 24627 2941 24639 2944
rect 24581 2935 24639 2941
rect 25133 2941 25145 2944
rect 25179 2941 25191 2975
rect 25133 2935 25191 2941
rect 20441 2907 20499 2913
rect 20441 2904 20453 2907
rect 12676 2876 20453 2904
rect 12676 2864 12682 2876
rect 20441 2873 20453 2876
rect 20487 2873 20499 2907
rect 20441 2867 20499 2873
rect 8386 2836 8392 2848
rect 8347 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 18138 2836 18144 2848
rect 13127 2808 18144 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 19015 2839 19073 2845
rect 19015 2805 19027 2839
rect 19061 2836 19073 2839
rect 19150 2836 19156 2848
rect 19061 2808 19156 2836
rect 19061 2805 19073 2808
rect 19015 2799 19073 2805
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 4387 2635 4445 2641
rect 4387 2601 4399 2635
rect 4433 2632 4445 2635
rect 6178 2632 6184 2644
rect 4433 2604 6184 2632
rect 4433 2601 4445 2604
rect 4387 2595 4445 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10367 2635 10425 2641
rect 10367 2632 10379 2635
rect 10100 2604 10379 2632
rect 10100 2592 10106 2604
rect 10367 2601 10379 2604
rect 10413 2601 10425 2635
rect 10367 2595 10425 2601
rect 12759 2635 12817 2641
rect 12759 2601 12771 2635
rect 12805 2632 12817 2635
rect 12894 2632 12900 2644
rect 12805 2604 12900 2632
rect 12805 2601 12817 2604
rect 12759 2595 12817 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 25222 2632 25228 2644
rect 25183 2604 25228 2632
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 4706 2496 4712 2508
rect 4362 2468 4712 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7576 2496 7604 2592
rect 11330 2524 11336 2576
rect 11388 2564 11394 2576
rect 11388 2536 13814 2564
rect 11388 2524 11394 2536
rect 6963 2468 7604 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 7892 2468 8585 2496
rect 7892 2456 7898 2468
rect 8573 2465 8585 2468
rect 8619 2496 8631 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8619 2468 9137 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9306 2456 9312 2508
rect 9364 2496 9370 2508
rect 10264 2499 10322 2505
rect 10264 2496 10276 2499
rect 9364 2468 10276 2496
rect 9364 2456 9370 2468
rect 10264 2465 10276 2468
rect 10310 2496 10322 2499
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10310 2468 10701 2496
rect 10310 2465 10322 2468
rect 10264 2459 10322 2465
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 12688 2499 12746 2505
rect 12688 2465 12700 2499
rect 12734 2496 12746 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12734 2468 13093 2496
rect 12734 2465 12746 2468
rect 12688 2459 12746 2465
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13786 2496 13814 2536
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 13786 2468 15945 2496
rect 13081 2459 13139 2465
rect 15933 2465 15945 2468
rect 15979 2496 15991 2499
rect 16485 2499 16543 2505
rect 16485 2496 16497 2499
rect 15979 2468 16497 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 16485 2465 16497 2468
rect 16531 2465 16543 2499
rect 19150 2496 19156 2508
rect 19111 2468 19156 2496
rect 16485 2459 16543 2465
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 12703 2428 12731 2459
rect 19150 2456 19156 2468
rect 19208 2496 19214 2508
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 19208 2468 19717 2496
rect 19208 2456 19214 2468
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 21361 2499 21419 2505
rect 21361 2465 21373 2499
rect 21407 2496 21419 2499
rect 21450 2496 21456 2508
rect 21407 2468 21456 2496
rect 21407 2465 21419 2468
rect 21361 2459 21419 2465
rect 21450 2456 21456 2468
rect 21508 2496 21514 2508
rect 21913 2499 21971 2505
rect 21913 2496 21925 2499
rect 21508 2468 21925 2496
rect 21508 2456 21514 2468
rect 21913 2465 21925 2468
rect 21959 2465 21971 2499
rect 21913 2459 21971 2465
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 25240 2496 25268 2592
rect 24627 2468 25268 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 6328 2400 12731 2428
rect 6328 2388 6334 2400
rect 8757 2363 8815 2369
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 10042 2360 10048 2372
rect 8803 2332 10048 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 16850 2320 16856 2372
rect 16908 2360 16914 2372
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 16908 2332 19349 2360
rect 16908 2320 16914 2332
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 27614 2360 27620 2372
rect 24811 2332 27620 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 27614 2320 27620 2332
rect 27672 2320 27678 2372
rect 4706 2292 4712 2304
rect 4667 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2292 16175 2295
rect 17770 2292 17776 2304
rect 16163 2264 17776 2292
rect 16163 2261 16175 2264
rect 16117 2255 16175 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 21545 2295 21603 2301
rect 21545 2261 21557 2295
rect 21591 2292 21603 2295
rect 23014 2292 23020 2304
rect 21591 2264 23020 2292
rect 21591 2261 21603 2264
rect 21545 2255 21603 2261
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 658 76 664 128
rect 716 116 722 128
rect 1302 116 1308 128
rect 716 88 1308 116
rect 716 76 722 88
rect 1302 76 1308 88
rect 1360 76 1366 128
<< via1 >>
rect 4436 27072 4488 27124
rect 5448 27072 5500 27124
rect 18972 26868 19024 26920
rect 23388 26868 23440 26920
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 10600 25304 10652 25356
rect 11152 25304 11204 25356
rect 14004 25304 14056 25356
rect 14740 25304 14792 25356
rect 10048 25100 10100 25152
rect 10784 25100 10836 25152
rect 12808 25143 12860 25152
rect 12808 25109 12817 25143
rect 12817 25109 12851 25143
rect 12851 25109 12860 25143
rect 12808 25100 12860 25109
rect 14096 25100 14148 25152
rect 14832 25100 14884 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 16396 24896 16448 24948
rect 10600 24871 10652 24880
rect 10600 24837 10609 24871
rect 10609 24837 10643 24871
rect 10643 24837 10652 24871
rect 10600 24828 10652 24837
rect 11796 24828 11848 24880
rect 11336 24760 11388 24812
rect 12808 24760 12860 24812
rect 8300 24692 8352 24744
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 11704 24692 11756 24744
rect 14004 24692 14056 24744
rect 14556 24692 14608 24744
rect 11152 24667 11204 24676
rect 11152 24633 11161 24667
rect 11161 24633 11195 24667
rect 11195 24633 11204 24667
rect 11152 24624 11204 24633
rect 12164 24624 12216 24676
rect 9036 24556 9088 24608
rect 9312 24556 9364 24608
rect 11704 24556 11756 24608
rect 12624 24556 12676 24608
rect 14464 24624 14516 24676
rect 15844 24624 15896 24676
rect 13728 24556 13780 24608
rect 14740 24556 14792 24608
rect 15936 24556 15988 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 11704 24352 11756 24404
rect 4712 24284 4764 24336
rect 6736 24284 6788 24336
rect 15384 24352 15436 24404
rect 17408 24352 17460 24404
rect 19432 24352 19484 24404
rect 27712 24352 27764 24404
rect 12624 24327 12676 24336
rect 12624 24293 12633 24327
rect 12633 24293 12667 24327
rect 12667 24293 12676 24327
rect 12624 24284 12676 24293
rect 13452 24284 13504 24336
rect 13912 24284 13964 24336
rect 6184 24216 6236 24268
rect 7564 24259 7616 24268
rect 7564 24225 7608 24259
rect 7608 24225 7616 24259
rect 7564 24216 7616 24225
rect 9404 24216 9456 24268
rect 10416 24259 10468 24268
rect 10416 24225 10425 24259
rect 10425 24225 10459 24259
rect 10459 24225 10468 24259
rect 10416 24216 10468 24225
rect 14004 24216 14056 24268
rect 15568 24216 15620 24268
rect 16580 24216 16632 24268
rect 17684 24216 17736 24268
rect 23112 24216 23164 24268
rect 25136 24216 25188 24268
rect 112 24080 164 24132
rect 13084 24123 13136 24132
rect 13084 24089 13093 24123
rect 13093 24089 13127 24123
rect 13127 24089 13136 24123
rect 13084 24080 13136 24089
rect 27620 24148 27672 24200
rect 6920 24012 6972 24064
rect 7840 24012 7892 24064
rect 9220 24012 9272 24064
rect 10876 24012 10928 24064
rect 12256 24055 12308 24064
rect 12256 24021 12265 24055
rect 12265 24021 12299 24055
rect 12299 24021 12308 24055
rect 12256 24012 12308 24021
rect 21916 24012 21968 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 6460 23808 6512 23860
rect 8392 23808 8444 23860
rect 9404 23808 9456 23860
rect 10140 23808 10192 23860
rect 10416 23808 10468 23860
rect 12348 23808 12400 23860
rect 16580 23851 16632 23860
rect 16580 23817 16589 23851
rect 16589 23817 16623 23851
rect 16623 23817 16632 23851
rect 16580 23808 16632 23817
rect 18236 23851 18288 23860
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 22376 23808 22428 23860
rect 24952 23808 25004 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 7564 23783 7616 23792
rect 7564 23749 7573 23783
rect 7573 23749 7607 23783
rect 7607 23749 7616 23783
rect 7564 23740 7616 23749
rect 13084 23783 13136 23792
rect 13084 23749 13093 23783
rect 13093 23749 13127 23783
rect 13127 23749 13136 23783
rect 13084 23740 13136 23749
rect 14004 23740 14056 23792
rect 14648 23740 14700 23792
rect 15384 23740 15436 23792
rect 12256 23672 12308 23724
rect 14096 23715 14148 23724
rect 14096 23681 14105 23715
rect 14105 23681 14139 23715
rect 14139 23681 14148 23715
rect 14096 23672 14148 23681
rect 14464 23715 14516 23724
rect 14464 23681 14473 23715
rect 14473 23681 14507 23715
rect 14507 23681 14516 23715
rect 14464 23672 14516 23681
rect 1124 23604 1176 23656
rect 5540 23604 5592 23656
rect 3792 23536 3844 23588
rect 5356 23536 5408 23588
rect 10140 23604 10192 23656
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 10968 23604 11020 23656
rect 19524 23740 19576 23792
rect 11152 23536 11204 23588
rect 11520 23579 11572 23588
rect 11520 23545 11529 23579
rect 11529 23545 11563 23579
rect 11563 23545 11572 23579
rect 11520 23536 11572 23545
rect 13544 23579 13596 23588
rect 4344 23468 4396 23520
rect 4896 23468 4948 23520
rect 6184 23511 6236 23520
rect 6184 23477 6193 23511
rect 6193 23477 6227 23511
rect 6227 23477 6236 23511
rect 6184 23468 6236 23477
rect 9128 23468 9180 23520
rect 12072 23468 12124 23520
rect 12256 23511 12308 23520
rect 12256 23477 12265 23511
rect 12265 23477 12299 23511
rect 12299 23477 12308 23511
rect 13544 23545 13553 23579
rect 13553 23545 13587 23579
rect 13587 23545 13596 23579
rect 13544 23536 13596 23545
rect 12256 23468 12308 23477
rect 13176 23468 13228 23520
rect 14280 23536 14332 23588
rect 17500 23536 17552 23588
rect 15660 23511 15712 23520
rect 15660 23477 15669 23511
rect 15669 23477 15703 23511
rect 15703 23477 15712 23511
rect 15660 23468 15712 23477
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 19064 23468 19116 23520
rect 27436 23740 27488 23792
rect 23112 23715 23164 23724
rect 23112 23681 23121 23715
rect 23121 23681 23155 23715
rect 23155 23681 23164 23715
rect 23112 23672 23164 23681
rect 25044 23672 25096 23724
rect 22928 23468 22980 23520
rect 23848 23468 23900 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5540 23264 5592 23316
rect 9128 23264 9180 23316
rect 10140 23264 10192 23316
rect 12072 23264 12124 23316
rect 12624 23264 12676 23316
rect 13176 23264 13228 23316
rect 4252 23239 4304 23248
rect 4252 23205 4261 23239
rect 4261 23205 4295 23239
rect 4295 23205 4304 23239
rect 4252 23196 4304 23205
rect 11704 23196 11756 23248
rect 13544 23196 13596 23248
rect 14096 23264 14148 23316
rect 14832 23196 14884 23248
rect 15936 23264 15988 23316
rect 17224 23264 17276 23316
rect 21456 23264 21508 23316
rect 15752 23196 15804 23248
rect 5172 23128 5224 23180
rect 6644 23128 6696 23180
rect 8024 23171 8076 23180
rect 8024 23137 8033 23171
rect 8033 23137 8067 23171
rect 8067 23137 8076 23171
rect 8024 23128 8076 23137
rect 8208 23171 8260 23180
rect 8208 23137 8217 23171
rect 8217 23137 8251 23171
rect 8251 23137 8260 23171
rect 8208 23128 8260 23137
rect 10232 23171 10284 23180
rect 10232 23137 10241 23171
rect 10241 23137 10275 23171
rect 10275 23137 10284 23171
rect 10232 23128 10284 23137
rect 11060 23128 11112 23180
rect 11520 23128 11572 23180
rect 12992 23171 13044 23180
rect 12992 23137 13001 23171
rect 13001 23137 13035 23171
rect 13035 23137 13044 23171
rect 12992 23128 13044 23137
rect 17408 23171 17460 23180
rect 17408 23137 17417 23171
rect 17417 23137 17451 23171
rect 17451 23137 17460 23171
rect 17408 23128 17460 23137
rect 17500 23128 17552 23180
rect 18972 23128 19024 23180
rect 3792 23060 3844 23112
rect 4528 23060 4580 23112
rect 8576 23060 8628 23112
rect 11980 23060 12032 23112
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14464 23060 14516 23112
rect 15476 23060 15528 23112
rect 17776 23103 17828 23112
rect 17776 23069 17785 23103
rect 17785 23069 17819 23103
rect 17819 23069 17828 23103
rect 17776 23060 17828 23069
rect 9956 22992 10008 23044
rect 2688 22967 2740 22976
rect 2688 22933 2697 22967
rect 2697 22933 2731 22967
rect 2731 22933 2740 22967
rect 2688 22924 2740 22933
rect 7380 22924 7432 22976
rect 7748 22924 7800 22976
rect 8208 22924 8260 22976
rect 11060 22967 11112 22976
rect 11060 22933 11069 22967
rect 11069 22933 11103 22967
rect 11103 22933 11112 22967
rect 11060 22924 11112 22933
rect 13084 22924 13136 22976
rect 14004 22924 14056 22976
rect 14556 22992 14608 23044
rect 20352 22992 20404 23044
rect 15292 22924 15344 22976
rect 16764 22924 16816 22976
rect 19892 22967 19944 22976
rect 19892 22933 19901 22967
rect 19901 22933 19935 22967
rect 19935 22933 19944 22967
rect 19892 22924 19944 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 4252 22720 4304 22772
rect 4344 22763 4396 22772
rect 4344 22729 4353 22763
rect 4353 22729 4387 22763
rect 4387 22729 4396 22763
rect 4344 22720 4396 22729
rect 4528 22720 4580 22772
rect 11980 22763 12032 22772
rect 11980 22729 11989 22763
rect 11989 22729 12023 22763
rect 12023 22729 12032 22763
rect 11980 22720 12032 22729
rect 13544 22720 13596 22772
rect 15752 22763 15804 22772
rect 112 22652 164 22704
rect 2688 22627 2740 22636
rect 2688 22593 2697 22627
rect 2697 22593 2731 22627
rect 2731 22593 2740 22627
rect 2688 22584 2740 22593
rect 6184 22584 6236 22636
rect 6644 22584 6696 22636
rect 7380 22584 7432 22636
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 10140 22584 10192 22636
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 4160 22448 4212 22500
rect 4344 22448 4396 22500
rect 5172 22491 5224 22500
rect 1492 22380 1544 22432
rect 5172 22457 5181 22491
rect 5181 22457 5215 22491
rect 5215 22457 5224 22491
rect 5172 22448 5224 22457
rect 4988 22380 5040 22432
rect 7564 22491 7616 22500
rect 6828 22380 6880 22432
rect 7564 22457 7573 22491
rect 7573 22457 7607 22491
rect 7607 22457 7616 22491
rect 7564 22448 7616 22457
rect 10232 22516 10284 22568
rect 15752 22729 15761 22763
rect 15761 22729 15795 22763
rect 15795 22729 15804 22763
rect 15752 22720 15804 22729
rect 17500 22720 17552 22772
rect 18972 22763 19024 22772
rect 18972 22729 18981 22763
rect 18981 22729 19015 22763
rect 19015 22729 19024 22763
rect 18972 22720 19024 22729
rect 15292 22584 15344 22636
rect 19432 22584 19484 22636
rect 19892 22627 19944 22636
rect 19892 22593 19901 22627
rect 19901 22593 19935 22627
rect 19935 22593 19944 22627
rect 19892 22584 19944 22593
rect 20260 22627 20312 22636
rect 20260 22593 20269 22627
rect 20269 22593 20303 22627
rect 20303 22593 20312 22627
rect 20260 22584 20312 22593
rect 16672 22516 16724 22568
rect 8760 22448 8812 22500
rect 10876 22448 10928 22500
rect 8024 22380 8076 22432
rect 9772 22380 9824 22432
rect 11704 22423 11756 22432
rect 11704 22389 11713 22423
rect 11713 22389 11747 22423
rect 11747 22389 11756 22423
rect 11704 22380 11756 22389
rect 13820 22380 13872 22432
rect 15476 22491 15528 22500
rect 15476 22457 15485 22491
rect 15485 22457 15519 22491
rect 15519 22457 15528 22491
rect 15476 22448 15528 22457
rect 16856 22448 16908 22500
rect 26424 22720 26476 22772
rect 24768 22695 24820 22704
rect 24768 22661 24777 22695
rect 24777 22661 24811 22695
rect 24811 22661 24820 22695
rect 24768 22652 24820 22661
rect 22008 22516 22060 22568
rect 20076 22448 20128 22500
rect 16212 22380 16264 22432
rect 17500 22380 17552 22432
rect 18328 22380 18380 22432
rect 20996 22380 21048 22432
rect 22652 22380 22704 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2688 22219 2740 22228
rect 2688 22185 2697 22219
rect 2697 22185 2731 22219
rect 2731 22185 2740 22219
rect 2688 22176 2740 22185
rect 4988 22219 5040 22228
rect 4988 22185 4997 22219
rect 4997 22185 5031 22219
rect 5031 22185 5040 22219
rect 4988 22176 5040 22185
rect 6828 22219 6880 22228
rect 6828 22185 6837 22219
rect 6837 22185 6871 22219
rect 6871 22185 6880 22219
rect 6828 22176 6880 22185
rect 9036 22219 9088 22228
rect 9036 22185 9045 22219
rect 9045 22185 9079 22219
rect 9079 22185 9088 22219
rect 9036 22176 9088 22185
rect 4160 22108 4212 22160
rect 6460 22108 6512 22160
rect 8668 22108 8720 22160
rect 2688 22083 2740 22092
rect 2688 22049 2697 22083
rect 2697 22049 2731 22083
rect 2731 22049 2740 22083
rect 2688 22040 2740 22049
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 5172 22040 5224 22092
rect 7564 22040 7616 22092
rect 8852 22040 8904 22092
rect 9220 22108 9272 22160
rect 10876 22176 10928 22228
rect 12256 22176 12308 22228
rect 13728 22176 13780 22228
rect 14832 22176 14884 22228
rect 15844 22176 15896 22228
rect 11704 22108 11756 22160
rect 13084 22108 13136 22160
rect 15936 22108 15988 22160
rect 17960 22151 18012 22160
rect 17960 22117 17969 22151
rect 17969 22117 18003 22151
rect 18003 22117 18012 22151
rect 17960 22108 18012 22117
rect 15384 22040 15436 22092
rect 16672 22040 16724 22092
rect 17776 22040 17828 22092
rect 19984 22176 20036 22228
rect 22008 22176 22060 22228
rect 20996 22151 21048 22160
rect 20996 22117 21005 22151
rect 21005 22117 21039 22151
rect 21039 22117 21048 22151
rect 20996 22108 21048 22117
rect 22284 22108 22336 22160
rect 20352 22040 20404 22092
rect 2504 21836 2556 21888
rect 3608 21836 3660 21888
rect 6000 21972 6052 22024
rect 7932 21972 7984 22024
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 10692 21972 10744 22024
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 15476 21972 15528 22024
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 21180 21972 21232 22024
rect 10876 21904 10928 21956
rect 11980 21904 12032 21956
rect 5540 21836 5592 21888
rect 7748 21836 7800 21888
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 11060 21836 11112 21888
rect 13084 21836 13136 21888
rect 14464 21904 14516 21956
rect 14280 21836 14332 21888
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2872 21632 2924 21684
rect 4160 21675 4212 21684
rect 4160 21641 4169 21675
rect 4169 21641 4203 21675
rect 4203 21641 4212 21675
rect 8852 21675 8904 21684
rect 4160 21632 4212 21641
rect 8852 21641 8861 21675
rect 8861 21641 8895 21675
rect 8895 21641 8904 21675
rect 8852 21632 8904 21641
rect 12716 21632 12768 21684
rect 7656 21564 7708 21616
rect 3608 21539 3660 21548
rect 2872 21471 2924 21480
rect 2872 21437 2881 21471
rect 2881 21437 2915 21471
rect 2915 21437 2924 21471
rect 2872 21428 2924 21437
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 6000 21496 6052 21548
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 11244 21496 11296 21548
rect 4988 21428 5040 21480
rect 5540 21360 5592 21412
rect 5724 21360 5776 21412
rect 7748 21428 7800 21480
rect 8760 21428 8812 21480
rect 2228 21292 2280 21344
rect 2688 21292 2740 21344
rect 4988 21335 5040 21344
rect 4988 21301 4997 21335
rect 4997 21301 5031 21335
rect 5031 21301 5040 21335
rect 4988 21292 5040 21301
rect 6460 21292 6512 21344
rect 8852 21360 8904 21412
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 13544 21564 13596 21616
rect 15384 21564 15436 21616
rect 17776 21632 17828 21684
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 22284 21675 22336 21684
rect 20076 21632 20128 21641
rect 22284 21641 22293 21675
rect 22293 21641 22327 21675
rect 22327 21641 22336 21675
rect 22284 21632 22336 21641
rect 22652 21675 22704 21684
rect 22652 21641 22661 21675
rect 22661 21641 22695 21675
rect 22695 21641 22704 21675
rect 22652 21632 22704 21641
rect 19064 21564 19116 21616
rect 20352 21607 20404 21616
rect 20352 21573 20361 21607
rect 20361 21573 20395 21607
rect 20395 21573 20404 21607
rect 20352 21564 20404 21573
rect 14004 21539 14056 21548
rect 14004 21505 14013 21539
rect 14013 21505 14047 21539
rect 14047 21505 14056 21539
rect 14004 21496 14056 21505
rect 15844 21496 15896 21548
rect 16488 21496 16540 21548
rect 10692 21360 10744 21412
rect 15200 21428 15252 21480
rect 15936 21428 15988 21480
rect 17040 21428 17092 21480
rect 18696 21496 18748 21548
rect 19248 21496 19300 21548
rect 21364 21471 21416 21480
rect 11244 21360 11296 21412
rect 13636 21403 13688 21412
rect 13636 21369 13645 21403
rect 13645 21369 13679 21403
rect 13679 21369 13688 21403
rect 13636 21360 13688 21369
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 12256 21292 12308 21344
rect 13820 21360 13872 21412
rect 17960 21360 18012 21412
rect 16672 21335 16724 21344
rect 16672 21301 16681 21335
rect 16681 21301 16715 21335
rect 16715 21301 16724 21335
rect 16672 21292 16724 21301
rect 18420 21292 18472 21344
rect 19340 21292 19392 21344
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 21272 21292 21324 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2228 21131 2280 21140
rect 2228 21097 2237 21131
rect 2237 21097 2271 21131
rect 2271 21097 2280 21131
rect 7932 21131 7984 21140
rect 2228 21088 2280 21097
rect 1952 21063 2004 21072
rect 1952 21029 1961 21063
rect 1961 21029 1995 21063
rect 1995 21029 2004 21063
rect 1952 21020 2004 21029
rect 2412 20995 2464 21004
rect 2412 20961 2421 20995
rect 2421 20961 2455 20995
rect 2455 20961 2464 20995
rect 2412 20952 2464 20961
rect 2504 20995 2556 21004
rect 2504 20961 2513 20995
rect 2513 20961 2547 20995
rect 2547 20961 2556 20995
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 8852 21088 8904 21140
rect 9220 21088 9272 21140
rect 2504 20952 2556 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 7012 21063 7064 21072
rect 7012 21029 7021 21063
rect 7021 21029 7055 21063
rect 7055 21029 7064 21063
rect 7012 21020 7064 21029
rect 7564 21063 7616 21072
rect 7564 21029 7573 21063
rect 7573 21029 7607 21063
rect 7607 21029 7616 21063
rect 7564 21020 7616 21029
rect 4068 20952 4120 20961
rect 2688 20816 2740 20868
rect 3884 20884 3936 20936
rect 5724 20952 5776 21004
rect 6000 20952 6052 21004
rect 8576 20952 8628 21004
rect 11336 21088 11388 21140
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 13452 21020 13504 21072
rect 13636 21088 13688 21140
rect 15292 21088 15344 21140
rect 15844 21131 15896 21140
rect 15844 21097 15853 21131
rect 15853 21097 15887 21131
rect 15887 21097 15896 21131
rect 15844 21088 15896 21097
rect 20076 21088 20128 21140
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 16488 21020 16540 21072
rect 16672 21020 16724 21072
rect 17132 21020 17184 21072
rect 18604 21020 18656 21072
rect 11152 20952 11204 21004
rect 11336 20952 11388 21004
rect 13820 20995 13872 21004
rect 13820 20961 13829 20995
rect 13829 20961 13863 20995
rect 13863 20961 13872 20995
rect 15384 20995 15436 21004
rect 13820 20952 13872 20961
rect 15384 20961 15402 20995
rect 15402 20961 15436 20995
rect 15384 20952 15436 20961
rect 15752 20952 15804 21004
rect 21272 20952 21324 21004
rect 22468 20995 22520 21004
rect 7656 20884 7708 20936
rect 9404 20884 9456 20936
rect 4160 20859 4212 20868
rect 4160 20825 4169 20859
rect 4169 20825 4203 20859
rect 4203 20825 4212 20859
rect 4160 20816 4212 20825
rect 9220 20816 9272 20868
rect 2136 20748 2188 20800
rect 5540 20748 5592 20800
rect 6276 20791 6328 20800
rect 6276 20757 6285 20791
rect 6285 20757 6319 20791
rect 6319 20757 6328 20791
rect 6276 20748 6328 20757
rect 7380 20748 7432 20800
rect 10140 20884 10192 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 13176 20884 13228 20936
rect 16764 20884 16816 20936
rect 16580 20816 16632 20868
rect 17868 20884 17920 20936
rect 18788 20884 18840 20936
rect 19432 20884 19484 20936
rect 22468 20961 22477 20995
rect 22477 20961 22511 20995
rect 22511 20961 22520 20995
rect 22468 20952 22520 20961
rect 24676 20952 24728 21004
rect 21456 20884 21508 20936
rect 17040 20816 17092 20868
rect 22744 20816 22796 20868
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 20352 20748 20404 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 480 20544 532 20596
rect 1768 20340 1820 20392
rect 2412 20544 2464 20596
rect 4160 20544 4212 20596
rect 7012 20544 7064 20596
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 9864 20544 9916 20596
rect 15384 20587 15436 20596
rect 6276 20408 6328 20460
rect 1400 20272 1452 20324
rect 1952 20272 2004 20324
rect 2228 20340 2280 20392
rect 3700 20383 3752 20392
rect 3700 20349 3709 20383
rect 3709 20349 3743 20383
rect 3743 20349 3752 20383
rect 3884 20383 3936 20392
rect 3700 20340 3752 20349
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 5172 20383 5224 20392
rect 5172 20349 5181 20383
rect 5181 20349 5215 20383
rect 5215 20349 5224 20383
rect 5172 20340 5224 20349
rect 5540 20340 5592 20392
rect 8668 20340 8720 20392
rect 4160 20272 4212 20324
rect 4252 20272 4304 20324
rect 6460 20272 6512 20324
rect 8852 20272 8904 20324
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 17868 20587 17920 20596
rect 17868 20553 17877 20587
rect 17877 20553 17911 20587
rect 17911 20553 17920 20587
rect 17868 20544 17920 20553
rect 18604 20544 18656 20596
rect 19432 20544 19484 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 10784 20476 10836 20528
rect 11152 20476 11204 20528
rect 13268 20476 13320 20528
rect 14004 20476 14056 20528
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 16120 20476 16172 20528
rect 14372 20408 14424 20460
rect 14464 20408 14516 20460
rect 17592 20476 17644 20528
rect 18512 20476 18564 20528
rect 16580 20451 16632 20460
rect 16580 20417 16589 20451
rect 16589 20417 16623 20451
rect 16623 20417 16632 20451
rect 16580 20408 16632 20417
rect 18420 20408 18472 20460
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 21272 20451 21324 20460
rect 21272 20417 21281 20451
rect 21281 20417 21315 20451
rect 21315 20417 21324 20451
rect 21272 20408 21324 20417
rect 22836 20408 22888 20460
rect 2412 20204 2464 20256
rect 4068 20204 4120 20256
rect 6000 20204 6052 20256
rect 6276 20247 6328 20256
rect 6276 20213 6285 20247
rect 6285 20213 6319 20247
rect 6319 20213 6328 20247
rect 6276 20204 6328 20213
rect 12256 20247 12308 20256
rect 12256 20213 12265 20247
rect 12265 20213 12299 20247
rect 12299 20213 12308 20247
rect 12256 20204 12308 20213
rect 13452 20204 13504 20256
rect 22008 20340 22060 20392
rect 18696 20315 18748 20324
rect 18696 20281 18705 20315
rect 18705 20281 18739 20315
rect 18739 20281 18748 20315
rect 18696 20272 18748 20281
rect 20352 20315 20404 20324
rect 20352 20281 20361 20315
rect 20361 20281 20395 20315
rect 20395 20281 20404 20315
rect 20352 20272 20404 20281
rect 21272 20272 21324 20324
rect 22468 20272 22520 20324
rect 16396 20204 16448 20256
rect 21824 20247 21876 20256
rect 21824 20213 21833 20247
rect 21833 20213 21867 20247
rect 21867 20213 21876 20247
rect 21824 20204 21876 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1952 20000 2004 20052
rect 1492 19864 1544 19916
rect 2136 20000 2188 20052
rect 7104 20000 7156 20052
rect 8852 20043 8904 20052
rect 8852 20009 8861 20043
rect 8861 20009 8895 20043
rect 8895 20009 8904 20043
rect 8852 20000 8904 20009
rect 9404 20043 9456 20052
rect 9404 20009 9413 20043
rect 9413 20009 9447 20043
rect 9447 20009 9456 20043
rect 9404 20000 9456 20009
rect 10784 20043 10836 20052
rect 10784 20009 10793 20043
rect 10793 20009 10827 20043
rect 10827 20009 10836 20043
rect 10784 20000 10836 20009
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 13636 20000 13688 20052
rect 14372 20043 14424 20052
rect 14372 20009 14381 20043
rect 14381 20009 14415 20043
rect 14415 20009 14424 20043
rect 14372 20000 14424 20009
rect 15660 20000 15712 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 16764 20043 16816 20052
rect 16764 20009 16773 20043
rect 16773 20009 16807 20043
rect 16807 20009 16816 20043
rect 16764 20000 16816 20009
rect 18604 20043 18656 20052
rect 18604 20009 18613 20043
rect 18613 20009 18647 20043
rect 18647 20009 18656 20043
rect 18604 20000 18656 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 20352 20000 20404 20052
rect 3884 19932 3936 19984
rect 6460 19932 6512 19984
rect 9772 19932 9824 19984
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2412 19864 2464 19873
rect 2228 19796 2280 19848
rect 3792 19864 3844 19916
rect 4068 19907 4120 19916
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 4344 19907 4396 19916
rect 4344 19873 4353 19907
rect 4353 19873 4387 19907
rect 4387 19873 4396 19907
rect 4344 19864 4396 19873
rect 2044 19728 2096 19780
rect 2780 19728 2832 19780
rect 3700 19728 3752 19780
rect 6092 19796 6144 19848
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 10048 19796 10100 19848
rect 10968 19932 11020 19984
rect 12256 19932 12308 19984
rect 13452 19932 13504 19984
rect 16304 19932 16356 19984
rect 17408 19975 17460 19984
rect 17408 19941 17417 19975
rect 17417 19941 17451 19975
rect 17451 19941 17460 19975
rect 17408 19932 17460 19941
rect 21088 19975 21140 19984
rect 14280 19864 14332 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16212 19864 16264 19916
rect 19248 19864 19300 19916
rect 21088 19941 21097 19975
rect 21097 19941 21131 19975
rect 21131 19941 21140 19975
rect 21088 19932 21140 19941
rect 22008 19975 22060 19984
rect 22008 19941 22017 19975
rect 22017 19941 22051 19975
rect 22051 19941 22060 19975
rect 22008 19932 22060 19941
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 22468 19907 22520 19916
rect 22468 19873 22477 19907
rect 22477 19873 22511 19907
rect 22511 19873 22520 19907
rect 22468 19864 22520 19873
rect 22836 19864 22888 19916
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 20996 19839 21048 19848
rect 1952 19660 2004 19712
rect 2596 19660 2648 19712
rect 4160 19660 4212 19712
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 7196 19660 7248 19712
rect 7656 19660 7708 19712
rect 18972 19728 19024 19780
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 21824 19728 21876 19780
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 13176 19660 13228 19712
rect 18420 19660 18472 19712
rect 21364 19660 21416 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1768 19499 1820 19508
rect 1768 19465 1777 19499
rect 1777 19465 1811 19499
rect 1811 19465 1820 19499
rect 1768 19456 1820 19465
rect 2412 19388 2464 19440
rect 2780 19388 2832 19440
rect 3976 19456 4028 19508
rect 4252 19456 4304 19508
rect 6092 19456 6144 19508
rect 9772 19499 9824 19508
rect 6460 19431 6512 19440
rect 6460 19397 6469 19431
rect 6469 19397 6503 19431
rect 6503 19397 6512 19431
rect 6460 19388 6512 19397
rect 7104 19363 7156 19372
rect 7104 19329 7113 19363
rect 7113 19329 7147 19363
rect 7147 19329 7156 19363
rect 7104 19320 7156 19329
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 17316 19456 17368 19508
rect 17408 19456 17460 19508
rect 17868 19456 17920 19508
rect 20628 19456 20680 19508
rect 21088 19456 21140 19508
rect 8576 19388 8628 19440
rect 14464 19388 14516 19440
rect 15844 19388 15896 19440
rect 18788 19388 18840 19440
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4344 19252 4396 19304
rect 5448 19295 5500 19304
rect 5448 19261 5457 19295
rect 5457 19261 5491 19295
rect 5491 19261 5500 19295
rect 5448 19252 5500 19261
rect 4160 19184 4212 19236
rect 4988 19184 5040 19236
rect 5540 19184 5592 19236
rect 6368 19252 6420 19304
rect 6276 19116 6328 19168
rect 7196 19227 7248 19236
rect 7196 19193 7205 19227
rect 7205 19193 7239 19227
rect 7239 19193 7248 19227
rect 7196 19184 7248 19193
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 13176 19363 13228 19372
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12164 19252 12216 19304
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 15660 19320 15712 19372
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 19248 19320 19300 19372
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 21272 19320 21324 19372
rect 14832 19295 14884 19304
rect 10968 19116 11020 19168
rect 12072 19116 12124 19168
rect 12256 19116 12308 19168
rect 14832 19261 14841 19295
rect 14841 19261 14875 19295
rect 14875 19261 14884 19295
rect 14832 19252 14884 19261
rect 15108 19184 15160 19236
rect 12532 19116 12584 19168
rect 13912 19116 13964 19168
rect 14280 19116 14332 19168
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 19248 19159 19300 19168
rect 16304 19116 16356 19125
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 19432 19116 19484 19168
rect 21272 19227 21324 19236
rect 21272 19193 21281 19227
rect 21281 19193 21315 19227
rect 21315 19193 21324 19227
rect 21272 19184 21324 19193
rect 22376 19184 22428 19236
rect 22836 19227 22888 19236
rect 22836 19193 22845 19227
rect 22845 19193 22879 19227
rect 22879 19193 22888 19227
rect 22836 19184 22888 19193
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 22468 19159 22520 19168
rect 22468 19125 22477 19159
rect 22477 19125 22511 19159
rect 22511 19125 22520 19159
rect 22468 19116 22520 19125
rect 23664 19159 23716 19168
rect 23664 19125 23673 19159
rect 23673 19125 23707 19159
rect 23707 19125 23716 19159
rect 23664 19116 23716 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 112 18912 164 18964
rect 6368 18955 6420 18964
rect 6368 18921 6377 18955
rect 6377 18921 6411 18955
rect 6411 18921 6420 18955
rect 6368 18912 6420 18921
rect 7656 18912 7708 18964
rect 7932 18912 7984 18964
rect 8484 18912 8536 18964
rect 9220 18912 9272 18964
rect 10048 18912 10100 18964
rect 12164 18912 12216 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 2412 18819 2464 18828
rect 2412 18785 2421 18819
rect 2421 18785 2455 18819
rect 2455 18785 2464 18819
rect 2412 18776 2464 18785
rect 2596 18844 2648 18896
rect 4252 18844 4304 18896
rect 7196 18844 7248 18896
rect 7840 18844 7892 18896
rect 12072 18844 12124 18896
rect 12532 18887 12584 18896
rect 12532 18853 12541 18887
rect 12541 18853 12575 18887
rect 12575 18853 12584 18887
rect 12532 18844 12584 18853
rect 13176 18887 13228 18896
rect 13176 18853 13185 18887
rect 13185 18853 13219 18887
rect 13219 18853 13228 18887
rect 13176 18844 13228 18853
rect 14096 18844 14148 18896
rect 18512 18912 18564 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 20628 18955 20680 18964
rect 15844 18887 15896 18896
rect 15844 18853 15853 18887
rect 15853 18853 15887 18887
rect 15887 18853 15896 18887
rect 15844 18844 15896 18853
rect 17408 18887 17460 18896
rect 17408 18853 17417 18887
rect 17417 18853 17451 18887
rect 17451 18853 17460 18887
rect 17408 18844 17460 18853
rect 19248 18844 19300 18896
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 20996 18912 21048 18964
rect 23664 18912 23716 18964
rect 21088 18887 21140 18896
rect 21088 18853 21097 18887
rect 21097 18853 21131 18887
rect 21131 18853 21140 18887
rect 21088 18844 21140 18853
rect 21180 18844 21232 18896
rect 2688 18819 2740 18828
rect 2688 18785 2697 18819
rect 2697 18785 2731 18819
rect 2731 18785 2740 18819
rect 2688 18776 2740 18785
rect 3700 18819 3752 18828
rect 3700 18785 3709 18819
rect 3709 18785 3743 18819
rect 3743 18785 3752 18819
rect 3700 18776 3752 18785
rect 4896 18776 4948 18828
rect 6092 18776 6144 18828
rect 9772 18819 9824 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 3332 18708 3384 18760
rect 5448 18708 5500 18760
rect 7012 18751 7064 18760
rect 2228 18640 2280 18692
rect 2688 18640 2740 18692
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 7472 18708 7524 18760
rect 9772 18785 9781 18819
rect 9781 18785 9815 18819
rect 9815 18785 9824 18819
rect 9772 18776 9824 18785
rect 9404 18708 9456 18760
rect 9496 18708 9548 18760
rect 22376 18776 22428 18828
rect 22836 18776 22888 18828
rect 24676 18776 24728 18828
rect 11612 18708 11664 18760
rect 13912 18708 13964 18760
rect 14832 18708 14884 18760
rect 15108 18751 15160 18760
rect 15108 18717 15117 18751
rect 15117 18717 15151 18751
rect 15151 18717 15160 18751
rect 15108 18708 15160 18717
rect 16212 18751 16264 18760
rect 7656 18640 7708 18692
rect 7932 18640 7984 18692
rect 9772 18640 9824 18692
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 1492 18572 1544 18624
rect 2136 18572 2188 18624
rect 3240 18572 3292 18624
rect 4988 18572 5040 18624
rect 5448 18572 5500 18624
rect 7012 18572 7064 18624
rect 8852 18572 8904 18624
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 9588 18572 9640 18624
rect 11244 18572 11296 18624
rect 12164 18615 12216 18624
rect 12164 18581 12173 18615
rect 12173 18581 12207 18615
rect 12207 18581 12216 18615
rect 12164 18572 12216 18581
rect 16856 18640 16908 18692
rect 18880 18640 18932 18692
rect 20628 18708 20680 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 17500 18572 17552 18624
rect 18328 18572 18380 18624
rect 22560 18572 22612 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2596 18411 2648 18420
rect 2596 18377 2605 18411
rect 2605 18377 2639 18411
rect 2639 18377 2648 18411
rect 2596 18368 2648 18377
rect 3332 18368 3384 18420
rect 3976 18368 4028 18420
rect 5356 18368 5408 18420
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 9404 18411 9456 18420
rect 9404 18377 9413 18411
rect 9413 18377 9447 18411
rect 9447 18377 9456 18411
rect 9404 18368 9456 18377
rect 11612 18411 11664 18420
rect 11612 18377 11621 18411
rect 11621 18377 11655 18411
rect 11655 18377 11664 18411
rect 11612 18368 11664 18377
rect 13176 18368 13228 18420
rect 13912 18411 13964 18420
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 13912 18368 13964 18377
rect 14832 18368 14884 18420
rect 15844 18368 15896 18420
rect 16856 18368 16908 18420
rect 17408 18368 17460 18420
rect 21272 18368 21324 18420
rect 24676 18368 24728 18420
rect 2044 18343 2096 18352
rect 2044 18309 2053 18343
rect 2053 18309 2087 18343
rect 2087 18309 2096 18343
rect 2044 18300 2096 18309
rect 3884 18300 3936 18352
rect 9036 18300 9088 18352
rect 16028 18343 16080 18352
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 8852 18232 8904 18284
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 16028 18309 16037 18343
rect 16037 18309 16071 18343
rect 16071 18309 16080 18343
rect 16028 18300 16080 18309
rect 18972 18300 19024 18352
rect 22376 18300 22428 18352
rect 10048 18232 10100 18241
rect 12256 18232 12308 18284
rect 20076 18232 20128 18284
rect 20904 18232 20956 18284
rect 22008 18232 22060 18284
rect 3884 18096 3936 18148
rect 4160 18139 4212 18148
rect 4160 18105 4169 18139
rect 4169 18105 4203 18139
rect 4203 18105 4212 18139
rect 4160 18096 4212 18105
rect 5264 18096 5316 18148
rect 3240 18028 3292 18080
rect 4252 18028 4304 18080
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 5540 18071 5592 18080
rect 5540 18037 5549 18071
rect 5549 18037 5583 18071
rect 5583 18037 5592 18071
rect 5540 18028 5592 18037
rect 6092 18071 6144 18080
rect 6092 18037 6101 18071
rect 6101 18037 6135 18071
rect 6135 18037 6144 18071
rect 6092 18028 6144 18037
rect 6368 18028 6420 18080
rect 6920 18164 6972 18216
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 15108 18207 15160 18216
rect 7932 18096 7984 18148
rect 9128 18139 9180 18148
rect 7104 18071 7156 18080
rect 7104 18037 7113 18071
rect 7113 18037 7147 18071
rect 7147 18037 7156 18071
rect 7104 18028 7156 18037
rect 9128 18105 9137 18139
rect 9137 18105 9171 18139
rect 9171 18105 9180 18139
rect 9128 18096 9180 18105
rect 9864 18096 9916 18148
rect 10140 18139 10192 18148
rect 10140 18105 10149 18139
rect 10149 18105 10183 18139
rect 10183 18105 10192 18139
rect 10140 18096 10192 18105
rect 10692 18139 10744 18148
rect 10692 18105 10701 18139
rect 10701 18105 10735 18139
rect 10735 18105 10744 18139
rect 10692 18096 10744 18105
rect 12164 18096 12216 18148
rect 13912 18096 13964 18148
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 14832 18096 14884 18148
rect 15844 18096 15896 18148
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 12072 18028 12124 18080
rect 13452 18028 13504 18080
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 18052 18164 18104 18216
rect 19340 18164 19392 18216
rect 19432 18096 19484 18148
rect 23572 18164 23624 18216
rect 24124 18164 24176 18216
rect 17500 18028 17552 18080
rect 19248 18028 19300 18080
rect 19340 18028 19392 18080
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 21272 18139 21324 18148
rect 21272 18105 21281 18139
rect 21281 18105 21315 18139
rect 21315 18105 21324 18139
rect 21272 18096 21324 18105
rect 22100 18096 22152 18148
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 22376 18028 22428 18080
rect 22836 18071 22888 18080
rect 22836 18037 22845 18071
rect 22845 18037 22879 18071
rect 22879 18037 22888 18071
rect 22836 18028 22888 18037
rect 23204 18028 23256 18080
rect 24584 18028 24636 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3884 17824 3936 17876
rect 4160 17824 4212 17876
rect 5356 17824 5408 17876
rect 6000 17867 6052 17876
rect 6000 17833 6009 17867
rect 6009 17833 6043 17867
rect 6043 17833 6052 17867
rect 6000 17824 6052 17833
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 10048 17824 10100 17876
rect 12164 17867 12216 17876
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 12624 17824 12676 17876
rect 13084 17824 13136 17876
rect 2504 17756 2556 17808
rect 4252 17756 4304 17808
rect 4436 17799 4488 17808
rect 4436 17765 4439 17799
rect 4439 17765 4473 17799
rect 4473 17765 4488 17799
rect 4436 17756 4488 17765
rect 1676 17688 1728 17740
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 9588 17756 9640 17808
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 12256 17756 12308 17808
rect 13452 17799 13504 17808
rect 13452 17765 13461 17799
rect 13461 17765 13495 17799
rect 13495 17765 13504 17799
rect 13452 17756 13504 17765
rect 13912 17756 13964 17808
rect 14096 17756 14148 17808
rect 2044 17620 2096 17672
rect 6276 17688 6328 17740
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 6368 17620 6420 17672
rect 8024 17620 8076 17672
rect 9496 17688 9548 17740
rect 9312 17620 9364 17672
rect 10876 17620 10928 17672
rect 11520 17620 11572 17672
rect 19432 17824 19484 17876
rect 20628 17867 20680 17876
rect 20628 17833 20637 17867
rect 20637 17833 20671 17867
rect 20671 17833 20680 17867
rect 20628 17824 20680 17833
rect 21088 17867 21140 17876
rect 21088 17833 21097 17867
rect 21097 17833 21131 17867
rect 21131 17833 21140 17867
rect 21088 17824 21140 17833
rect 16028 17799 16080 17808
rect 16028 17765 16037 17799
rect 16037 17765 16071 17799
rect 16071 17765 16080 17799
rect 16028 17756 16080 17765
rect 18880 17799 18932 17808
rect 18880 17765 18889 17799
rect 18889 17765 18923 17799
rect 18923 17765 18932 17799
rect 18880 17756 18932 17765
rect 20076 17799 20128 17808
rect 17408 17731 17460 17740
rect 17408 17697 17417 17731
rect 17417 17697 17451 17731
rect 17451 17697 17460 17731
rect 17408 17688 17460 17697
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 18972 17731 19024 17740
rect 18972 17697 18981 17731
rect 18981 17697 19015 17731
rect 19015 17697 19024 17731
rect 18972 17688 19024 17697
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 1952 17552 2004 17604
rect 4252 17552 4304 17604
rect 2044 17484 2096 17536
rect 4068 17484 4120 17536
rect 5080 17484 5132 17536
rect 15108 17552 15160 17604
rect 18144 17620 18196 17672
rect 20076 17765 20085 17799
rect 20085 17765 20119 17799
rect 20119 17765 20128 17799
rect 20076 17756 20128 17765
rect 21824 17756 21876 17808
rect 22836 17688 22888 17740
rect 24124 17688 24176 17740
rect 20076 17620 20128 17672
rect 21916 17620 21968 17672
rect 16212 17552 16264 17604
rect 17316 17595 17368 17604
rect 17316 17561 17325 17595
rect 17325 17561 17359 17595
rect 17359 17561 17368 17595
rect 23204 17620 23256 17672
rect 17316 17552 17368 17561
rect 22100 17595 22152 17604
rect 22100 17561 22109 17595
rect 22109 17561 22143 17595
rect 22143 17561 22152 17595
rect 22100 17552 22152 17561
rect 22744 17552 22796 17604
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 8944 17484 8996 17536
rect 10784 17484 10836 17536
rect 13544 17484 13596 17536
rect 14832 17484 14884 17536
rect 15936 17484 15988 17536
rect 22008 17484 22060 17536
rect 23296 17484 23348 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 5448 17280 5500 17332
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8208 17280 8260 17332
rect 11520 17323 11572 17332
rect 1400 17212 1452 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 3976 17144 4028 17196
rect 5356 17144 5408 17196
rect 8576 17144 8628 17196
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 13912 17280 13964 17332
rect 16028 17280 16080 17332
rect 17408 17323 17460 17332
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 18328 17323 18380 17332
rect 18328 17289 18337 17323
rect 18337 17289 18371 17323
rect 18371 17289 18380 17323
rect 18328 17280 18380 17289
rect 18972 17280 19024 17332
rect 22192 17280 22244 17332
rect 13176 17212 13228 17264
rect 13268 17212 13320 17264
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9956 17144 10008 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 14004 17144 14056 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2044 17076 2096 17128
rect 5080 17076 5132 17128
rect 7748 17076 7800 17128
rect 14740 17119 14792 17128
rect 14740 17085 14749 17119
rect 14749 17085 14783 17119
rect 14783 17085 14792 17119
rect 14740 17076 14792 17085
rect 14832 17076 14884 17128
rect 17868 17212 17920 17264
rect 17960 17212 18012 17264
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 24124 17212 24176 17264
rect 16580 17187 16632 17196
rect 16580 17153 16589 17187
rect 16589 17153 16623 17187
rect 16623 17153 16632 17187
rect 16580 17144 16632 17153
rect 24032 17144 24084 17196
rect 22284 17076 22336 17128
rect 23756 17119 23808 17128
rect 23756 17085 23774 17119
rect 23774 17085 23808 17119
rect 23756 17076 23808 17085
rect 5448 17008 5500 17060
rect 2688 16940 2740 16992
rect 3608 16940 3660 16992
rect 4436 16940 4488 16992
rect 6276 16983 6328 16992
rect 6276 16949 6285 16983
rect 6285 16949 6319 16983
rect 6319 16949 6328 16983
rect 6276 16940 6328 16949
rect 7012 16940 7064 16992
rect 7472 17008 7524 17060
rect 8944 17051 8996 17060
rect 8944 17017 8953 17051
rect 8953 17017 8987 17051
rect 8987 17017 8996 17051
rect 8944 17008 8996 17017
rect 12624 17051 12676 17060
rect 9864 16940 9916 16992
rect 12624 17017 12633 17051
rect 12633 17017 12667 17051
rect 12667 17017 12676 17051
rect 12624 17008 12676 17017
rect 14924 17008 14976 17060
rect 16212 17051 16264 17060
rect 16212 17017 16221 17051
rect 16221 17017 16255 17051
rect 16255 17017 16264 17051
rect 16212 17008 16264 17017
rect 16304 17051 16356 17060
rect 16304 17017 16313 17051
rect 16313 17017 16347 17051
rect 16347 17017 16356 17051
rect 16304 17008 16356 17017
rect 20720 17008 20772 17060
rect 20996 17051 21048 17060
rect 20996 17017 21005 17051
rect 21005 17017 21039 17051
rect 21039 17017 21048 17051
rect 20996 17008 21048 17017
rect 21640 17008 21692 17060
rect 12164 16940 12216 16992
rect 12808 16940 12860 16992
rect 14004 16983 14056 16992
rect 14004 16949 14013 16983
rect 14013 16949 14047 16983
rect 14047 16949 14056 16983
rect 14004 16940 14056 16949
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 19248 16983 19300 16992
rect 19248 16949 19257 16983
rect 19257 16949 19291 16983
rect 19291 16949 19300 16983
rect 19248 16940 19300 16949
rect 20444 16940 20496 16992
rect 20536 16940 20588 16992
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 22836 16940 22888 16992
rect 23204 16940 23256 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 4436 16779 4488 16788
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 4620 16736 4672 16788
rect 5540 16736 5592 16788
rect 7748 16779 7800 16788
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 9312 16736 9364 16788
rect 9956 16736 10008 16788
rect 14832 16736 14884 16788
rect 5264 16668 5316 16720
rect 1952 16575 2004 16584
rect 1952 16541 1961 16575
rect 1961 16541 1995 16575
rect 1995 16541 2004 16575
rect 1952 16532 2004 16541
rect 2504 16532 2556 16584
rect 2872 16600 2924 16652
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 4252 16600 4304 16652
rect 9496 16668 9548 16720
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 10048 16668 10100 16720
rect 13452 16668 13504 16720
rect 14924 16668 14976 16720
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 6092 16600 6144 16652
rect 6828 16600 6880 16652
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 8392 16600 8444 16652
rect 11060 16600 11112 16652
rect 12072 16643 12124 16652
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 16304 16736 16356 16788
rect 17868 16736 17920 16788
rect 20996 16736 21048 16788
rect 21916 16779 21968 16788
rect 21916 16745 21925 16779
rect 21925 16745 21959 16779
rect 21959 16745 21968 16779
rect 21916 16736 21968 16745
rect 24032 16736 24084 16788
rect 16120 16668 16172 16720
rect 20076 16668 20128 16720
rect 20444 16668 20496 16720
rect 20812 16668 20864 16720
rect 21824 16668 21876 16720
rect 22560 16711 22612 16720
rect 22560 16677 22569 16711
rect 22569 16677 22603 16711
rect 22603 16677 22612 16711
rect 22560 16668 22612 16677
rect 22652 16711 22704 16720
rect 22652 16677 22661 16711
rect 22661 16677 22695 16711
rect 22695 16677 22704 16711
rect 22652 16668 22704 16677
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 24216 16643 24268 16652
rect 24216 16609 24225 16643
rect 24225 16609 24259 16643
rect 24259 16609 24268 16643
rect 24216 16600 24268 16609
rect 3884 16575 3936 16584
rect 3884 16541 3893 16575
rect 3893 16541 3927 16575
rect 3927 16541 3936 16575
rect 3884 16532 3936 16541
rect 6644 16575 6696 16584
rect 6644 16541 6653 16575
rect 6653 16541 6687 16575
rect 6687 16541 6696 16575
rect 6644 16532 6696 16541
rect 10876 16532 10928 16584
rect 4068 16464 4120 16516
rect 4712 16464 4764 16516
rect 7748 16464 7800 16516
rect 8300 16464 8352 16516
rect 8484 16464 8536 16516
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 19524 16532 19576 16584
rect 20444 16532 20496 16584
rect 13268 16464 13320 16516
rect 2964 16396 3016 16448
rect 3056 16396 3108 16448
rect 7012 16396 7064 16448
rect 7656 16396 7708 16448
rect 8760 16396 8812 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 20720 16439 20772 16448
rect 20720 16405 20729 16439
rect 20729 16405 20763 16439
rect 20763 16405 20772 16439
rect 20720 16396 20772 16405
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 22100 16532 22152 16584
rect 22744 16532 22796 16584
rect 24124 16464 24176 16516
rect 20996 16396 21048 16448
rect 23204 16396 23256 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1952 16192 2004 16244
rect 2872 16192 2924 16244
rect 4436 16192 4488 16244
rect 6000 16167 6052 16176
rect 6000 16133 6009 16167
rect 6009 16133 6043 16167
rect 6043 16133 6052 16167
rect 8208 16192 8260 16244
rect 9864 16192 9916 16244
rect 12072 16235 12124 16244
rect 12072 16201 12081 16235
rect 12081 16201 12115 16235
rect 12115 16201 12124 16235
rect 12072 16192 12124 16201
rect 12624 16235 12676 16244
rect 12624 16201 12633 16235
rect 12633 16201 12667 16235
rect 12667 16201 12676 16235
rect 12624 16192 12676 16201
rect 13176 16192 13228 16244
rect 14096 16192 14148 16244
rect 6000 16124 6052 16133
rect 8760 16124 8812 16176
rect 12808 16124 12860 16176
rect 15292 16192 15344 16244
rect 16120 16235 16172 16244
rect 16120 16201 16129 16235
rect 16129 16201 16163 16235
rect 16163 16201 16172 16235
rect 16120 16192 16172 16201
rect 17224 16235 17276 16244
rect 17224 16201 17233 16235
rect 17233 16201 17267 16235
rect 17267 16201 17276 16235
rect 17224 16192 17276 16201
rect 20536 16235 20588 16244
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 20720 16192 20772 16244
rect 16488 16167 16540 16176
rect 16488 16133 16497 16167
rect 16497 16133 16531 16167
rect 16531 16133 16540 16167
rect 16488 16124 16540 16133
rect 1676 16056 1728 16108
rect 8944 16056 8996 16108
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 9956 16056 10008 16108
rect 13452 16056 13504 16108
rect 15384 16056 15436 16108
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 7932 15988 7984 16040
rect 8484 15988 8536 16040
rect 14924 15988 14976 16040
rect 3516 15920 3568 15972
rect 4620 15963 4672 15972
rect 4620 15929 4629 15963
rect 4629 15929 4663 15963
rect 4663 15929 4672 15963
rect 4620 15920 4672 15929
rect 4712 15963 4764 15972
rect 4712 15929 4721 15963
rect 4721 15929 4755 15963
rect 4755 15929 4764 15963
rect 5264 15963 5316 15972
rect 4712 15920 4764 15929
rect 5264 15929 5273 15963
rect 5273 15929 5307 15963
rect 5307 15929 5316 15963
rect 5264 15920 5316 15929
rect 112 15852 164 15904
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 6000 15852 6052 15904
rect 7012 15852 7064 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 8760 15963 8812 15972
rect 8760 15929 8769 15963
rect 8769 15929 8803 15963
rect 8803 15929 8812 15963
rect 10232 15963 10284 15972
rect 8760 15920 8812 15929
rect 9312 15852 9364 15904
rect 10232 15929 10241 15963
rect 10241 15929 10275 15963
rect 10275 15929 10284 15963
rect 10232 15920 10284 15929
rect 10876 15963 10928 15972
rect 9772 15852 9824 15904
rect 10876 15929 10885 15963
rect 10885 15929 10919 15963
rect 10919 15929 10928 15963
rect 10876 15920 10928 15929
rect 13360 15963 13412 15972
rect 13360 15929 13369 15963
rect 13369 15929 13403 15963
rect 13403 15929 13412 15963
rect 13360 15920 13412 15929
rect 13452 15963 13504 15972
rect 13452 15929 13461 15963
rect 13461 15929 13495 15963
rect 13495 15929 13504 15963
rect 13452 15920 13504 15929
rect 14740 15920 14792 15972
rect 15292 15920 15344 15972
rect 17960 16124 18012 16176
rect 20812 16167 20864 16176
rect 20812 16133 20821 16167
rect 20821 16133 20855 16167
rect 20855 16133 20864 16167
rect 20812 16124 20864 16133
rect 21088 16124 21140 16176
rect 17868 16056 17920 16108
rect 18420 15988 18472 16040
rect 19984 16056 20036 16108
rect 21916 16056 21968 16108
rect 22560 16124 22612 16176
rect 24216 16124 24268 16176
rect 22652 16056 22704 16108
rect 22928 16056 22980 16108
rect 23112 16056 23164 16108
rect 22836 15988 22888 16040
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 22100 15963 22152 15972
rect 19248 15852 19300 15904
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 22100 15920 22152 15929
rect 22560 15920 22612 15972
rect 21272 15852 21324 15861
rect 22192 15852 22244 15904
rect 22376 15852 22428 15904
rect 22652 15852 22704 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 7012 15648 7064 15700
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 13452 15648 13504 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 14004 15648 14056 15700
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 3148 15623 3200 15632
rect 3148 15589 3157 15623
rect 3157 15589 3191 15623
rect 3191 15589 3200 15623
rect 3148 15580 3200 15589
rect 7932 15623 7984 15632
rect 7932 15589 7941 15623
rect 7941 15589 7975 15623
rect 7975 15589 7984 15623
rect 7932 15580 7984 15589
rect 9496 15623 9548 15632
rect 9496 15589 9505 15623
rect 9505 15589 9539 15623
rect 9539 15589 9548 15623
rect 9496 15580 9548 15589
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 21272 15648 21324 15700
rect 22008 15691 22060 15700
rect 22008 15657 22017 15691
rect 22017 15657 22051 15691
rect 22051 15657 22060 15691
rect 22008 15648 22060 15657
rect 22192 15648 22244 15700
rect 15752 15623 15804 15632
rect 2228 15512 2280 15564
rect 3700 15512 3752 15564
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 5080 15512 5132 15564
rect 6000 15512 6052 15564
rect 8392 15512 8444 15564
rect 8484 15512 8536 15564
rect 11152 15512 11204 15564
rect 12256 15512 12308 15564
rect 15752 15589 15761 15623
rect 15761 15589 15795 15623
rect 15795 15589 15804 15623
rect 15752 15580 15804 15589
rect 19524 15580 19576 15632
rect 20996 15580 21048 15632
rect 21088 15623 21140 15632
rect 21088 15589 21097 15623
rect 21097 15589 21131 15623
rect 21131 15589 21140 15623
rect 22560 15623 22612 15632
rect 21088 15580 21140 15589
rect 22560 15589 22569 15623
rect 22569 15589 22603 15623
rect 22603 15589 22612 15623
rect 22560 15580 22612 15589
rect 23020 15648 23072 15700
rect 24124 15691 24176 15700
rect 24124 15657 24133 15691
rect 24133 15657 24167 15691
rect 24167 15657 24176 15691
rect 24124 15648 24176 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 23204 15580 23256 15632
rect 14372 15512 14424 15564
rect 2872 15444 2924 15496
rect 2964 15444 3016 15496
rect 4620 15444 4672 15496
rect 8116 15444 8168 15496
rect 10048 15487 10100 15496
rect 9496 15376 9548 15428
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 17868 15512 17920 15564
rect 24676 15512 24728 15564
rect 10876 15376 10928 15428
rect 16212 15419 16264 15428
rect 16212 15385 16221 15419
rect 16221 15385 16255 15419
rect 16255 15385 16264 15419
rect 16212 15376 16264 15385
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 2688 15351 2740 15360
rect 2688 15317 2697 15351
rect 2697 15317 2731 15351
rect 2731 15317 2740 15351
rect 2688 15308 2740 15317
rect 3424 15351 3476 15360
rect 3424 15317 3433 15351
rect 3433 15317 3467 15351
rect 3467 15317 3476 15351
rect 3424 15308 3476 15317
rect 4252 15308 4304 15360
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 8852 15308 8904 15360
rect 9312 15308 9364 15360
rect 9404 15308 9456 15360
rect 10140 15308 10192 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 11244 15308 11296 15360
rect 12532 15308 12584 15360
rect 17132 15308 17184 15360
rect 18144 15444 18196 15496
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 21824 15444 21876 15496
rect 17960 15376 18012 15428
rect 19064 15376 19116 15428
rect 20720 15376 20772 15428
rect 22100 15376 22152 15428
rect 18512 15351 18564 15360
rect 18512 15317 18521 15351
rect 18521 15317 18555 15351
rect 18555 15317 18564 15351
rect 18512 15308 18564 15317
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 20904 15308 20956 15360
rect 22744 15444 22796 15496
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1860 15104 1912 15156
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 3884 15104 3936 15156
rect 8116 15147 8168 15156
rect 8116 15113 8125 15147
rect 8125 15113 8159 15147
rect 8159 15113 8168 15147
rect 8116 15104 8168 15113
rect 9864 15104 9916 15156
rect 12256 15147 12308 15156
rect 12256 15113 12265 15147
rect 12265 15113 12299 15147
rect 12299 15113 12308 15147
rect 12256 15104 12308 15113
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 14372 15104 14424 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 17868 15104 17920 15156
rect 18420 15104 18472 15156
rect 19340 15104 19392 15156
rect 21088 15104 21140 15156
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 23204 15147 23256 15156
rect 23204 15113 23213 15147
rect 23213 15113 23247 15147
rect 23247 15113 23256 15147
rect 23204 15104 23256 15113
rect 2688 15036 2740 15088
rect 3148 15079 3200 15088
rect 3148 15045 3172 15079
rect 3172 15045 3200 15079
rect 3148 15036 3200 15045
rect 3792 15036 3844 15088
rect 4160 14968 4212 15020
rect 2320 14900 2372 14952
rect 2412 14900 2464 14952
rect 3424 14900 3476 14952
rect 10784 15036 10836 15088
rect 15660 15036 15712 15088
rect 21732 15036 21784 15088
rect 8300 14968 8352 15020
rect 10048 14968 10100 15020
rect 11152 14968 11204 15020
rect 12624 14968 12676 15020
rect 5172 14943 5224 14952
rect 5172 14909 5181 14943
rect 5181 14909 5215 14943
rect 5215 14909 5224 14943
rect 5172 14900 5224 14909
rect 5448 14900 5500 14952
rect 6000 14900 6052 14952
rect 2044 14832 2096 14884
rect 2780 14832 2832 14884
rect 2872 14832 2924 14884
rect 13084 14900 13136 14952
rect 14740 14968 14792 15020
rect 17592 14968 17644 15020
rect 19892 14968 19944 15020
rect 20536 14968 20588 15020
rect 21088 14968 21140 15020
rect 18420 14943 18472 14952
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 18512 14900 18564 14952
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 22376 15036 22428 15088
rect 22560 14968 22612 15020
rect 23572 14900 23624 14952
rect 9128 14875 9180 14884
rect 9128 14841 9137 14875
rect 9137 14841 9171 14875
rect 9171 14841 9180 14875
rect 9128 14832 9180 14841
rect 9220 14875 9272 14884
rect 9220 14841 9229 14875
rect 9229 14841 9263 14875
rect 9263 14841 9272 14875
rect 9220 14832 9272 14841
rect 9956 14832 10008 14884
rect 3884 14764 3936 14816
rect 4252 14764 4304 14816
rect 7012 14764 7064 14816
rect 8484 14764 8536 14816
rect 10784 14875 10836 14884
rect 10784 14841 10793 14875
rect 10793 14841 10827 14875
rect 10827 14841 10836 14875
rect 10784 14832 10836 14841
rect 12532 14832 12584 14884
rect 14372 14832 14424 14884
rect 15660 14875 15712 14884
rect 15660 14841 15669 14875
rect 15669 14841 15703 14875
rect 15703 14841 15712 14875
rect 15660 14832 15712 14841
rect 15752 14875 15804 14884
rect 15752 14841 15761 14875
rect 15761 14841 15795 14875
rect 15795 14841 15804 14875
rect 15752 14832 15804 14841
rect 18696 14832 18748 14884
rect 20904 14875 20956 14884
rect 20904 14841 20913 14875
rect 20913 14841 20947 14875
rect 20947 14841 20956 14875
rect 20904 14832 20956 14841
rect 21088 14832 21140 14884
rect 21640 14832 21692 14884
rect 11060 14764 11112 14816
rect 12808 14764 12860 14816
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 21180 14764 21232 14816
rect 23940 14764 23992 14816
rect 24676 14764 24728 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2596 14560 2648 14612
rect 4988 14560 5040 14612
rect 5172 14603 5224 14612
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 7012 14492 7064 14544
rect 8484 14535 8536 14544
rect 8484 14501 8493 14535
rect 8493 14501 8527 14535
rect 8527 14501 8536 14535
rect 8484 14492 8536 14501
rect 9128 14560 9180 14612
rect 9404 14492 9456 14544
rect 9772 14492 9824 14544
rect 10876 14560 10928 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11980 14560 12032 14612
rect 16948 14603 17000 14612
rect 10692 14492 10744 14544
rect 11796 14535 11848 14544
rect 11796 14501 11805 14535
rect 11805 14501 11839 14535
rect 11839 14501 11848 14535
rect 11796 14492 11848 14501
rect 2136 14424 2188 14476
rect 3516 14467 3568 14476
rect 3516 14433 3525 14467
rect 3525 14433 3559 14467
rect 3559 14433 3568 14467
rect 3516 14424 3568 14433
rect 4620 14424 4672 14476
rect 5448 14424 5500 14476
rect 6000 14424 6052 14476
rect 6644 14424 6696 14476
rect 8668 14467 8720 14476
rect 8668 14433 8686 14467
rect 8686 14433 8720 14467
rect 8668 14424 8720 14433
rect 9036 14424 9088 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 13912 14492 13964 14544
rect 15476 14535 15528 14544
rect 15476 14501 15485 14535
rect 15485 14501 15519 14535
rect 15519 14501 15528 14535
rect 15476 14492 15528 14501
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 18696 14603 18748 14612
rect 18696 14569 18705 14603
rect 18705 14569 18739 14603
rect 18739 14569 18748 14603
rect 18696 14560 18748 14569
rect 20904 14560 20956 14612
rect 17500 14492 17552 14544
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 21640 14535 21692 14544
rect 21640 14501 21649 14535
rect 21649 14501 21683 14535
rect 21683 14501 21692 14535
rect 21640 14492 21692 14501
rect 21732 14492 21784 14544
rect 12624 14424 12676 14476
rect 13452 14467 13504 14476
rect 4160 14356 4212 14408
rect 5356 14356 5408 14408
rect 7196 14356 7248 14408
rect 7656 14356 7708 14408
rect 9496 14356 9548 14408
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 22744 14424 22796 14476
rect 24124 14424 24176 14476
rect 13544 14356 13596 14408
rect 15384 14399 15436 14408
rect 15384 14365 15393 14399
rect 15393 14365 15427 14399
rect 15427 14365 15436 14399
rect 15384 14356 15436 14365
rect 16764 14356 16816 14408
rect 20720 14356 20772 14408
rect 2228 14288 2280 14340
rect 2320 14288 2372 14340
rect 3148 14288 3200 14340
rect 4528 14288 4580 14340
rect 9220 14288 9272 14340
rect 17684 14288 17736 14340
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4252 14263 4304 14272
rect 4252 14229 4276 14263
rect 4276 14229 4304 14263
rect 4252 14220 4304 14229
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 8944 14220 8996 14272
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 19708 14263 19760 14272
rect 19708 14229 19717 14263
rect 19717 14229 19751 14263
rect 19751 14229 19760 14263
rect 19708 14220 19760 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1952 13812 2004 13864
rect 2688 14016 2740 14068
rect 3884 14016 3936 14068
rect 6552 14016 6604 14068
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 9772 14016 9824 14068
rect 11980 14059 12032 14068
rect 11980 14025 11989 14059
rect 11989 14025 12023 14059
rect 12023 14025 12032 14059
rect 11980 14016 12032 14025
rect 6000 13991 6052 14000
rect 6000 13957 6009 13991
rect 6009 13957 6043 13991
rect 6043 13957 6052 13991
rect 6000 13948 6052 13957
rect 6736 13948 6788 14000
rect 7104 13948 7156 14000
rect 12808 13948 12860 14000
rect 13728 13948 13780 14000
rect 3608 13880 3660 13932
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 4436 13880 4488 13932
rect 5356 13880 5408 13932
rect 7932 13880 7984 13932
rect 8852 13880 8904 13932
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 16948 14016 17000 14068
rect 17408 14016 17460 14068
rect 17868 14016 17920 14068
rect 18420 14016 18472 14068
rect 20536 14059 20588 14068
rect 20536 14025 20545 14059
rect 20545 14025 20579 14059
rect 20579 14025 20588 14059
rect 20536 14016 20588 14025
rect 21088 14016 21140 14068
rect 23848 14016 23900 14068
rect 24952 14059 25004 14068
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 17132 13948 17184 14000
rect 19432 13948 19484 14000
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 8392 13812 8444 13864
rect 13544 13812 13596 13864
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 17316 13880 17368 13932
rect 19708 13880 19760 13932
rect 17868 13812 17920 13864
rect 18512 13812 18564 13864
rect 18880 13812 18932 13864
rect 21180 13855 21232 13864
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 21180 13812 21232 13821
rect 2412 13744 2464 13796
rect 3056 13787 3108 13796
rect 3056 13753 3065 13787
rect 3065 13753 3099 13787
rect 3099 13753 3108 13787
rect 3056 13744 3108 13753
rect 3792 13787 3844 13796
rect 3792 13753 3801 13787
rect 3801 13753 3835 13787
rect 3835 13753 3844 13787
rect 3792 13744 3844 13753
rect 6000 13744 6052 13796
rect 9220 13787 9272 13796
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 9220 13744 9272 13753
rect 10692 13787 10744 13796
rect 10692 13753 10701 13787
rect 10701 13753 10735 13787
rect 10735 13753 10744 13787
rect 10692 13744 10744 13753
rect 10784 13787 10836 13796
rect 10784 13753 10793 13787
rect 10793 13753 10827 13787
rect 10827 13753 10836 13787
rect 10784 13744 10836 13753
rect 11428 13744 11480 13796
rect 12808 13744 12860 13796
rect 2780 13676 2832 13728
rect 3516 13676 3568 13728
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 4528 13676 4580 13685
rect 6184 13676 6236 13728
rect 7012 13676 7064 13728
rect 7840 13676 7892 13728
rect 8300 13676 8352 13728
rect 13360 13676 13412 13728
rect 15476 13744 15528 13796
rect 15200 13676 15252 13728
rect 16028 13744 16080 13796
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 19156 13676 19208 13728
rect 19524 13744 19576 13796
rect 20536 13676 20588 13728
rect 21180 13676 21232 13728
rect 21456 13855 21508 13864
rect 21456 13821 21465 13855
rect 21465 13821 21499 13855
rect 21499 13821 21508 13855
rect 21456 13812 21508 13821
rect 21916 13855 21968 13864
rect 21916 13821 21925 13855
rect 21925 13821 21959 13855
rect 21959 13821 21968 13855
rect 21916 13812 21968 13821
rect 23020 13812 23072 13864
rect 24676 13855 24728 13864
rect 24676 13821 24720 13855
rect 24720 13821 24728 13855
rect 24676 13812 24728 13821
rect 22744 13787 22796 13796
rect 22744 13753 22753 13787
rect 22753 13753 22787 13787
rect 22787 13753 22796 13787
rect 22744 13744 22796 13753
rect 24124 13719 24176 13728
rect 24124 13685 24133 13719
rect 24133 13685 24167 13719
rect 24167 13685 24176 13719
rect 24124 13676 24176 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13472 1728 13524
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 2136 13472 2188 13524
rect 3608 13472 3660 13524
rect 9404 13515 9456 13524
rect 5264 13404 5316 13456
rect 6184 13404 6236 13456
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 7748 13404 7800 13456
rect 10784 13472 10836 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13452 13472 13504 13524
rect 15292 13472 15344 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 20812 13472 20864 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 2136 13336 2188 13388
rect 3056 13336 3108 13388
rect 3332 13336 3384 13388
rect 3700 13336 3752 13388
rect 4160 13336 4212 13388
rect 7104 13336 7156 13388
rect 9680 13336 9732 13388
rect 11244 13404 11296 13456
rect 13360 13447 13412 13456
rect 13360 13413 13369 13447
rect 13369 13413 13403 13447
rect 13403 13413 13412 13447
rect 13360 13404 13412 13413
rect 14372 13404 14424 13456
rect 15384 13404 15436 13456
rect 16212 13404 16264 13456
rect 16948 13404 17000 13456
rect 19156 13404 19208 13456
rect 10692 13336 10744 13388
rect 22744 13404 22796 13456
rect 20904 13379 20956 13388
rect 3424 13268 3476 13320
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 6000 13268 6052 13320
rect 2412 13200 2464 13252
rect 4528 13200 4580 13252
rect 4620 13200 4672 13252
rect 5356 13200 5408 13252
rect 8484 13268 8536 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13636 13268 13688 13320
rect 14280 13268 14332 13320
rect 16764 13268 16816 13320
rect 17040 13268 17092 13320
rect 17132 13200 17184 13252
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 21180 13336 21232 13388
rect 21916 13336 21968 13388
rect 22192 13336 22244 13388
rect 22652 13336 22704 13388
rect 23020 13379 23072 13388
rect 23020 13345 23029 13379
rect 23029 13345 23063 13379
rect 23063 13345 23072 13379
rect 23020 13336 23072 13345
rect 24216 13336 24268 13388
rect 24676 13336 24728 13388
rect 21088 13200 21140 13252
rect 21180 13200 21232 13252
rect 22468 13200 22520 13252
rect 2320 13132 2372 13184
rect 3516 13132 3568 13184
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 4988 13132 5040 13184
rect 5172 13132 5224 13184
rect 8116 13132 8168 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 9220 13132 9272 13184
rect 17684 13132 17736 13184
rect 18512 13132 18564 13184
rect 20536 13132 20588 13184
rect 21272 13132 21324 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2688 12928 2740 12980
rect 4436 12928 4488 12980
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 6184 12928 6236 12980
rect 7104 12928 7156 12980
rect 7748 12971 7800 12980
rect 7748 12937 7757 12971
rect 7757 12937 7791 12971
rect 7791 12937 7800 12971
rect 7748 12928 7800 12937
rect 8944 12928 8996 12980
rect 11612 12928 11664 12980
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 15384 12928 15436 12980
rect 16028 12928 16080 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 23020 12928 23072 12980
rect 2320 12860 2372 12912
rect 3792 12860 3844 12912
rect 4620 12860 4672 12912
rect 6552 12903 6604 12912
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 6552 12869 6561 12903
rect 6561 12869 6595 12903
rect 6595 12869 6604 12903
rect 6552 12860 6604 12869
rect 10692 12903 10744 12912
rect 10692 12869 10701 12903
rect 10701 12869 10735 12903
rect 10735 12869 10744 12903
rect 10692 12860 10744 12869
rect 10784 12860 10836 12912
rect 11244 12860 11296 12912
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 3148 12724 3200 12776
rect 5264 12792 5316 12844
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9772 12792 9824 12844
rect 4988 12724 5040 12776
rect 5448 12724 5500 12776
rect 6368 12724 6420 12776
rect 7472 12724 7524 12776
rect 3332 12656 3384 12708
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2228 12588 2280 12640
rect 7656 12656 7708 12708
rect 8024 12699 8076 12708
rect 8024 12665 8033 12699
rect 8033 12665 8067 12699
rect 8067 12665 8076 12699
rect 8024 12656 8076 12665
rect 8392 12656 8444 12708
rect 10140 12699 10192 12708
rect 6920 12588 6972 12640
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 7564 12588 7616 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 10140 12665 10149 12699
rect 10149 12665 10183 12699
rect 10183 12665 10192 12699
rect 10140 12656 10192 12665
rect 10600 12656 10652 12708
rect 11428 12724 11480 12776
rect 12164 12724 12216 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 15936 12792 15988 12844
rect 17040 12792 17092 12844
rect 18052 12860 18104 12912
rect 22468 12860 22520 12912
rect 18604 12792 18656 12844
rect 21364 12792 21416 12844
rect 21548 12835 21600 12844
rect 21548 12801 21557 12835
rect 21557 12801 21591 12835
rect 21591 12801 21600 12835
rect 21548 12792 21600 12801
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 10968 12588 11020 12640
rect 12900 12588 12952 12640
rect 13452 12588 13504 12640
rect 14464 12656 14516 12708
rect 18512 12767 18564 12776
rect 18512 12733 18521 12767
rect 18521 12733 18555 12767
rect 18555 12733 18564 12767
rect 18512 12724 18564 12733
rect 20812 12724 20864 12776
rect 16396 12656 16448 12708
rect 21180 12699 21232 12708
rect 21180 12665 21189 12699
rect 21189 12665 21223 12699
rect 21223 12665 21232 12699
rect 21180 12656 21232 12665
rect 21272 12699 21324 12708
rect 21272 12665 21281 12699
rect 21281 12665 21315 12699
rect 21315 12665 21324 12699
rect 21272 12656 21324 12665
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 16580 12631 16632 12640
rect 16580 12597 16589 12631
rect 16589 12597 16623 12631
rect 16623 12597 16632 12631
rect 16580 12588 16632 12597
rect 19156 12631 19208 12640
rect 19156 12597 19165 12631
rect 19165 12597 19199 12631
rect 19199 12597 19208 12631
rect 19156 12588 19208 12597
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20720 12588 20772 12640
rect 22192 12588 22244 12640
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 24216 12588 24268 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 4436 12384 4488 12436
rect 4620 12427 4672 12436
rect 4620 12393 4629 12427
rect 4629 12393 4663 12427
rect 4663 12393 4672 12427
rect 4620 12384 4672 12393
rect 8392 12384 8444 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 8852 12384 8904 12436
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 19156 12384 19208 12436
rect 20720 12384 20772 12436
rect 21180 12384 21232 12436
rect 23664 12384 23716 12436
rect 5356 12316 5408 12368
rect 7104 12316 7156 12368
rect 7564 12316 7616 12368
rect 7656 12316 7708 12368
rect 10140 12316 10192 12368
rect 10876 12359 10928 12368
rect 10876 12325 10885 12359
rect 10885 12325 10919 12359
rect 10919 12325 10928 12359
rect 10876 12316 10928 12325
rect 11428 12359 11480 12368
rect 11428 12325 11437 12359
rect 11437 12325 11471 12359
rect 11471 12325 11480 12359
rect 11428 12316 11480 12325
rect 11796 12316 11848 12368
rect 16580 12316 16632 12368
rect 17132 12316 17184 12368
rect 20260 12316 20312 12368
rect 20628 12316 20680 12368
rect 2044 12248 2096 12300
rect 4068 12248 4120 12300
rect 6000 12248 6052 12300
rect 9864 12248 9916 12300
rect 14372 12248 14424 12300
rect 17776 12291 17828 12300
rect 17776 12257 17785 12291
rect 17785 12257 17819 12291
rect 17819 12257 17828 12291
rect 17776 12248 17828 12257
rect 20812 12248 20864 12300
rect 22468 12291 22520 12300
rect 22468 12257 22512 12291
rect 22512 12257 22520 12291
rect 22468 12248 22520 12257
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 4344 12180 4396 12232
rect 6460 12180 6512 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 12348 12223 12400 12232
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 13360 12223 13412 12232
rect 2412 12112 2464 12164
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 2320 12044 2372 12096
rect 2964 12044 3016 12096
rect 3332 12044 3384 12096
rect 7840 12112 7892 12164
rect 10692 12112 10744 12164
rect 11428 12112 11480 12164
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 16672 12180 16724 12232
rect 18236 12180 18288 12232
rect 21272 12112 21324 12164
rect 21548 12155 21600 12164
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 6368 12044 6420 12096
rect 8116 12044 8168 12096
rect 9956 12044 10008 12096
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 15384 12044 15436 12096
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 18972 12044 19024 12096
rect 19064 12044 19116 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1952 11883 2004 11892
rect 1952 11849 1961 11883
rect 1961 11849 1995 11883
rect 1995 11849 2004 11883
rect 1952 11840 2004 11849
rect 2044 11840 2096 11892
rect 3976 11840 4028 11892
rect 2228 11815 2280 11824
rect 2228 11781 2252 11815
rect 2252 11781 2280 11815
rect 2228 11772 2280 11781
rect 2320 11704 2372 11756
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 6368 11840 6420 11892
rect 6920 11840 6972 11892
rect 9864 11840 9916 11892
rect 10876 11840 10928 11892
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 12440 11840 12492 11892
rect 12808 11883 12860 11892
rect 12808 11849 12817 11883
rect 12817 11849 12851 11883
rect 12851 11849 12860 11883
rect 12808 11840 12860 11849
rect 1952 11636 2004 11688
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 5540 11636 5592 11688
rect 10692 11704 10744 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 13728 11772 13780 11824
rect 15476 11840 15528 11892
rect 16580 11840 16632 11892
rect 19340 11840 19392 11892
rect 14648 11772 14700 11824
rect 14280 11704 14332 11756
rect 16028 11704 16080 11756
rect 16396 11747 16448 11756
rect 16396 11713 16405 11747
rect 16405 11713 16439 11747
rect 16439 11713 16448 11747
rect 16396 11704 16448 11713
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 2780 11611 2832 11620
rect 2780 11577 2789 11611
rect 2789 11577 2823 11611
rect 2823 11577 2832 11611
rect 2780 11568 2832 11577
rect 6092 11568 6144 11620
rect 6368 11568 6420 11620
rect 7104 11568 7156 11620
rect 9128 11636 9180 11688
rect 10508 11636 10560 11688
rect 20536 11840 20588 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 20076 11679 20128 11688
rect 20076 11645 20085 11679
rect 20085 11645 20119 11679
rect 20119 11645 20128 11679
rect 20076 11636 20128 11645
rect 20812 11636 20864 11688
rect 21088 11636 21140 11688
rect 24584 11679 24636 11688
rect 24584 11645 24593 11679
rect 24593 11645 24627 11679
rect 24627 11645 24636 11679
rect 24584 11636 24636 11645
rect 9496 11568 9548 11620
rect 9864 11568 9916 11620
rect 12808 11568 12860 11620
rect 13360 11568 13412 11620
rect 14372 11568 14424 11620
rect 14832 11611 14884 11620
rect 14832 11577 14864 11611
rect 14864 11577 14884 11611
rect 14832 11568 14884 11577
rect 14924 11611 14976 11620
rect 14924 11577 14933 11611
rect 14933 11577 14967 11611
rect 14967 11577 14976 11611
rect 14924 11568 14976 11577
rect 18236 11611 18288 11620
rect 18236 11577 18245 11611
rect 18245 11577 18279 11611
rect 18279 11577 18288 11611
rect 18236 11568 18288 11577
rect 19340 11568 19392 11620
rect 21548 11568 21600 11620
rect 6644 11543 6696 11552
rect 6644 11509 6653 11543
rect 6653 11509 6687 11543
rect 6687 11509 6696 11543
rect 6644 11500 6696 11509
rect 7840 11500 7892 11552
rect 9036 11500 9088 11552
rect 17776 11543 17828 11552
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 19156 11543 19208 11552
rect 19156 11509 19165 11543
rect 19165 11509 19199 11543
rect 19199 11509 19208 11543
rect 19156 11500 19208 11509
rect 19984 11500 20036 11552
rect 20812 11500 20864 11552
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 24676 11500 24728 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4344 11296 4396 11348
rect 5540 11296 5592 11348
rect 9036 11296 9088 11348
rect 12348 11296 12400 11348
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 14556 11296 14608 11348
rect 14924 11296 14976 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 6368 11228 6420 11280
rect 6460 11228 6512 11280
rect 7840 11228 7892 11280
rect 9864 11271 9916 11280
rect 9864 11237 9873 11271
rect 9873 11237 9907 11271
rect 9907 11237 9916 11271
rect 9864 11228 9916 11237
rect 9956 11228 10008 11280
rect 10600 11228 10652 11280
rect 11428 11228 11480 11280
rect 15384 11271 15436 11280
rect 15384 11237 15393 11271
rect 15393 11237 15427 11271
rect 15427 11237 15436 11271
rect 15384 11228 15436 11237
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 18236 11296 18288 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 20628 11339 20680 11348
rect 20628 11305 20637 11339
rect 20637 11305 20671 11339
rect 20671 11305 20680 11339
rect 20628 11296 20680 11305
rect 15476 11228 15528 11237
rect 21088 11271 21140 11280
rect 21088 11237 21097 11271
rect 21097 11237 21131 11271
rect 21131 11237 21140 11271
rect 21088 11228 21140 11237
rect 1308 11160 1360 11212
rect 2872 11160 2924 11212
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 2320 11092 2372 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 1584 11024 1636 11076
rect 2412 11067 2464 11076
rect 2412 11033 2421 11067
rect 2421 11033 2455 11067
rect 2455 11033 2464 11067
rect 2412 11024 2464 11033
rect 3792 11024 3844 11076
rect 4160 11024 4212 11076
rect 4436 11024 4488 11076
rect 7380 11092 7432 11144
rect 8024 11092 8076 11144
rect 17868 11160 17920 11212
rect 18420 11203 18472 11212
rect 18420 11169 18429 11203
rect 18429 11169 18463 11203
rect 18463 11169 18472 11203
rect 18420 11160 18472 11169
rect 8944 11024 8996 11076
rect 10968 11024 11020 11076
rect 16764 11092 16816 11144
rect 17592 11092 17644 11144
rect 22284 11160 22336 11212
rect 23112 11160 23164 11212
rect 20076 11092 20128 11144
rect 20444 11092 20496 11144
rect 22008 11092 22060 11144
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 15936 11067 15988 11076
rect 15936 11033 15945 11067
rect 15945 11033 15979 11067
rect 15979 11033 15988 11067
rect 15936 11024 15988 11033
rect 17132 11024 17184 11076
rect 22192 11024 22244 11076
rect 3332 10956 3384 11008
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6644 10956 6696 11008
rect 7012 10956 7064 11008
rect 12992 10956 13044 11008
rect 14096 10956 14148 11008
rect 19064 10956 19116 11008
rect 20996 10956 21048 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1952 10752 2004 10804
rect 3424 10752 3476 10804
rect 4344 10752 4396 10804
rect 5080 10795 5132 10804
rect 5080 10761 5089 10795
rect 5089 10761 5123 10795
rect 5123 10761 5132 10795
rect 5080 10752 5132 10761
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 9956 10752 10008 10804
rect 14648 10752 14700 10804
rect 15384 10752 15436 10804
rect 18420 10752 18472 10804
rect 21088 10795 21140 10804
rect 21088 10761 21097 10795
rect 21097 10761 21131 10795
rect 21131 10761 21140 10795
rect 21088 10752 21140 10761
rect 10600 10684 10652 10736
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 14556 10684 14608 10736
rect 15476 10684 15528 10736
rect 15936 10727 15988 10736
rect 15936 10693 15945 10727
rect 15945 10693 15979 10727
rect 15979 10693 15988 10727
rect 15936 10684 15988 10693
rect 24768 10727 24820 10736
rect 3056 10616 3108 10668
rect 4620 10659 4672 10668
rect 4620 10625 4629 10659
rect 4629 10625 4663 10659
rect 4663 10625 4672 10659
rect 4620 10616 4672 10625
rect 5540 10616 5592 10668
rect 1676 10591 1728 10600
rect 1676 10557 1685 10591
rect 1685 10557 1719 10591
rect 1719 10557 1728 10591
rect 1676 10548 1728 10557
rect 1860 10548 1912 10600
rect 5080 10548 5132 10600
rect 8484 10616 8536 10668
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 8208 10548 8260 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 3056 10523 3108 10532
rect 3056 10489 3065 10523
rect 3065 10489 3099 10523
rect 3099 10489 3108 10523
rect 3056 10480 3108 10489
rect 3700 10523 3752 10532
rect 1308 10412 1360 10464
rect 2872 10455 2924 10464
rect 2872 10421 2881 10455
rect 2881 10421 2915 10455
rect 2915 10421 2924 10455
rect 2872 10412 2924 10421
rect 3700 10489 3709 10523
rect 3709 10489 3743 10523
rect 3743 10489 3752 10523
rect 3700 10480 3752 10489
rect 6092 10480 6144 10532
rect 6920 10523 6972 10532
rect 6920 10489 6929 10523
rect 6929 10489 6963 10523
rect 6963 10489 6972 10523
rect 6920 10480 6972 10489
rect 7564 10523 7616 10532
rect 5172 10412 5224 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 7564 10489 7573 10523
rect 7573 10489 7607 10523
rect 7607 10489 7616 10523
rect 7564 10480 7616 10489
rect 8116 10480 8168 10532
rect 9588 10480 9640 10532
rect 14096 10616 14148 10668
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 15568 10616 15620 10668
rect 17224 10616 17276 10668
rect 18512 10616 18564 10668
rect 19984 10616 20036 10668
rect 24768 10693 24777 10727
rect 24777 10693 24811 10727
rect 24811 10693 24820 10727
rect 24768 10684 24820 10693
rect 21916 10616 21968 10668
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 12716 10548 12768 10600
rect 10692 10523 10744 10532
rect 9864 10455 9916 10464
rect 6552 10412 6604 10421
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 10692 10489 10701 10523
rect 10701 10489 10735 10523
rect 10735 10489 10744 10523
rect 10692 10480 10744 10489
rect 11980 10480 12032 10532
rect 13084 10480 13136 10532
rect 13728 10523 13780 10532
rect 13728 10489 13737 10523
rect 13737 10489 13771 10523
rect 13771 10489 13780 10523
rect 13728 10480 13780 10489
rect 15384 10523 15436 10532
rect 15384 10489 15393 10523
rect 15393 10489 15427 10523
rect 15427 10489 15436 10523
rect 15384 10480 15436 10489
rect 15476 10523 15528 10532
rect 15476 10489 15485 10523
rect 15485 10489 15519 10523
rect 15519 10489 15528 10523
rect 15476 10480 15528 10489
rect 16856 10548 16908 10600
rect 19064 10548 19116 10600
rect 17776 10455 17828 10464
rect 9864 10412 9916 10421
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 19156 10412 19208 10464
rect 24124 10548 24176 10600
rect 22284 10412 22336 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1676 10208 1728 10260
rect 3056 10208 3108 10260
rect 6460 10208 6512 10260
rect 6552 10208 6604 10260
rect 3148 10140 3200 10192
rect 3424 10183 3476 10192
rect 3424 10149 3433 10183
rect 3433 10149 3467 10183
rect 3467 10149 3476 10183
rect 3424 10140 3476 10149
rect 5540 10140 5592 10192
rect 7380 10208 7432 10260
rect 7840 10251 7892 10260
rect 7840 10217 7849 10251
rect 7849 10217 7883 10251
rect 7883 10217 7892 10251
rect 7840 10208 7892 10217
rect 12992 10251 13044 10260
rect 6828 10140 6880 10192
rect 9220 10140 9272 10192
rect 9956 10183 10008 10192
rect 9956 10149 9965 10183
rect 9965 10149 9999 10183
rect 9999 10149 10008 10183
rect 9956 10140 10008 10149
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 13728 10208 13780 10260
rect 14648 10208 14700 10260
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20444 10208 20496 10260
rect 21916 10251 21968 10260
rect 21916 10217 21925 10251
rect 21925 10217 21959 10251
rect 21959 10217 21968 10251
rect 21916 10208 21968 10217
rect 11704 10140 11756 10192
rect 2044 10072 2096 10124
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 4252 10072 4304 10124
rect 7196 10072 7248 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 12624 10072 12676 10124
rect 18420 10140 18472 10192
rect 19064 10183 19116 10192
rect 19064 10149 19073 10183
rect 19073 10149 19107 10183
rect 19107 10149 19116 10183
rect 19064 10140 19116 10149
rect 21088 10183 21140 10192
rect 21088 10149 21097 10183
rect 21097 10149 21131 10183
rect 21131 10149 21140 10183
rect 21088 10140 21140 10149
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 14740 10072 14792 10124
rect 15660 10072 15712 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 17592 10072 17644 10124
rect 22468 10115 22520 10124
rect 22468 10081 22512 10115
rect 22512 10081 22520 10115
rect 22468 10072 22520 10081
rect 24216 10072 24268 10124
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 8760 10047 8812 10056
rect 7012 9936 7064 9988
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 9680 10004 9732 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 11520 10004 11572 10056
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18972 10047 19024 10056
rect 18972 10013 18981 10047
rect 18981 10013 19015 10047
rect 19015 10013 19024 10047
rect 18972 10004 19024 10013
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 6828 9868 6880 9920
rect 11060 9936 11112 9988
rect 10692 9868 10744 9920
rect 10968 9868 11020 9920
rect 14740 9868 14792 9920
rect 15384 9868 15436 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 22100 9868 22152 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 4712 9664 4764 9716
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 8024 9707 8076 9716
rect 8024 9673 8033 9707
rect 8033 9673 8067 9707
rect 8067 9673 8076 9707
rect 8024 9664 8076 9673
rect 9864 9707 9916 9716
rect 9864 9673 9873 9707
rect 9873 9673 9907 9707
rect 9907 9673 9916 9707
rect 9864 9664 9916 9673
rect 9956 9664 10008 9716
rect 10140 9707 10192 9716
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 13360 9664 13412 9716
rect 15660 9664 15712 9716
rect 15844 9664 15896 9716
rect 5172 9639 5224 9648
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 5172 9605 5181 9639
rect 5181 9605 5215 9639
rect 5215 9605 5224 9639
rect 5172 9596 5224 9605
rect 10876 9596 10928 9648
rect 11060 9596 11112 9648
rect 13544 9596 13596 9648
rect 6828 9528 6880 9580
rect 7472 9528 7524 9580
rect 8760 9528 8812 9580
rect 15200 9596 15252 9648
rect 17316 9664 17368 9716
rect 19064 9664 19116 9716
rect 21088 9664 21140 9716
rect 22468 9707 22520 9716
rect 22468 9673 22477 9707
rect 22477 9673 22511 9707
rect 22511 9673 22520 9707
rect 22468 9664 22520 9673
rect 19616 9596 19668 9648
rect 21272 9596 21324 9648
rect 21456 9596 21508 9648
rect 22928 9596 22980 9648
rect 17224 9528 17276 9580
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 20260 9528 20312 9580
rect 22100 9528 22152 9580
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 1492 9460 1544 9512
rect 2044 9460 2096 9512
rect 2228 9460 2280 9512
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 2504 9460 2556 9469
rect 2596 9460 2648 9512
rect 4804 9392 4856 9444
rect 5540 9392 5592 9444
rect 2596 9324 2648 9376
rect 2964 9324 3016 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 7104 9435 7156 9444
rect 7104 9401 7113 9435
rect 7113 9401 7147 9435
rect 7147 9401 7156 9435
rect 7104 9392 7156 9401
rect 7288 9392 7340 9444
rect 7840 9324 7892 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9956 9392 10008 9444
rect 10784 9435 10836 9444
rect 10784 9401 10793 9435
rect 10793 9401 10827 9435
rect 10827 9401 10836 9435
rect 10784 9392 10836 9401
rect 10876 9435 10928 9444
rect 10876 9401 10885 9435
rect 10885 9401 10919 9435
rect 10919 9401 10928 9435
rect 10876 9392 10928 9401
rect 12808 9392 12860 9444
rect 14832 9435 14884 9444
rect 14832 9401 14841 9435
rect 14841 9401 14875 9435
rect 14875 9401 14884 9435
rect 14832 9392 14884 9401
rect 14924 9435 14976 9444
rect 14924 9401 14933 9435
rect 14933 9401 14967 9435
rect 14967 9401 14976 9435
rect 15476 9435 15528 9444
rect 14924 9392 14976 9401
rect 15476 9401 15485 9435
rect 15485 9401 15519 9435
rect 15519 9401 15528 9435
rect 15476 9392 15528 9401
rect 16488 9435 16540 9444
rect 16488 9401 16497 9435
rect 16497 9401 16531 9435
rect 16531 9401 16540 9435
rect 16488 9392 16540 9401
rect 16580 9435 16632 9444
rect 16580 9401 16589 9435
rect 16589 9401 16623 9435
rect 16623 9401 16632 9435
rect 16580 9392 16632 9401
rect 18236 9392 18288 9444
rect 11612 9324 11664 9376
rect 12624 9324 12676 9376
rect 13728 9324 13780 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 17316 9324 17368 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 21456 9435 21508 9444
rect 17776 9324 17828 9333
rect 21456 9401 21465 9435
rect 21465 9401 21499 9435
rect 21499 9401 21508 9435
rect 21456 9392 21508 9401
rect 21548 9435 21600 9444
rect 21548 9401 21557 9435
rect 21557 9401 21591 9435
rect 21591 9401 21600 9435
rect 22100 9435 22152 9444
rect 21548 9392 21600 9401
rect 22100 9401 22109 9435
rect 22109 9401 22143 9435
rect 22143 9401 22152 9435
rect 22100 9392 22152 9401
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 7104 9120 7156 9172
rect 8760 9120 8812 9172
rect 9956 9120 10008 9172
rect 10140 9120 10192 9172
rect 11428 9120 11480 9172
rect 13728 9120 13780 9172
rect 18052 9120 18104 9172
rect 18972 9120 19024 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20996 9120 21048 9172
rect 21548 9120 21600 9172
rect 4712 9095 4764 9104
rect 4712 9061 4721 9095
rect 4721 9061 4755 9095
rect 4755 9061 4764 9095
rect 4712 9052 4764 9061
rect 5540 9052 5592 9104
rect 6644 9052 6696 9104
rect 6828 9052 6880 9104
rect 9680 9052 9732 9104
rect 12992 9052 13044 9104
rect 13268 9052 13320 9104
rect 14556 9052 14608 9104
rect 14924 9052 14976 9104
rect 19892 9052 19944 9104
rect 21732 9052 21784 9104
rect 112 8984 164 9036
rect 1768 8984 1820 9036
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 2504 8916 2556 8968
rect 3148 8984 3200 9036
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8576 9027 8628 9036
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 8576 8984 8628 8993
rect 11520 8984 11572 9036
rect 17592 8984 17644 9036
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 18880 9027 18932 9036
rect 18880 8993 18889 9027
rect 18889 8993 18923 9027
rect 18923 8993 18932 9027
rect 18880 8984 18932 8993
rect 21824 8984 21876 9036
rect 23112 8984 23164 9036
rect 3884 8916 3936 8968
rect 2964 8848 3016 8900
rect 3700 8848 3752 8900
rect 7288 8916 7340 8968
rect 9404 8916 9456 8968
rect 11060 8916 11112 8968
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 11980 8848 12032 8900
rect 15200 8848 15252 8900
rect 15292 8848 15344 8900
rect 15936 8891 15988 8900
rect 15936 8857 15945 8891
rect 15945 8857 15979 8891
rect 15979 8857 15988 8891
rect 15936 8848 15988 8857
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 17224 8959 17276 8968
rect 16948 8916 17000 8925
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 17684 8916 17736 8968
rect 18972 8916 19024 8968
rect 20260 8916 20312 8968
rect 2044 8780 2096 8832
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 4896 8780 4948 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 9956 8780 10008 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 16580 8780 16632 8832
rect 17684 8780 17736 8832
rect 18236 8848 18288 8900
rect 21180 8848 21232 8900
rect 21272 8848 21324 8900
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 3332 8576 3384 8628
rect 4712 8576 4764 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9864 8576 9916 8628
rect 11060 8619 11112 8628
rect 1584 8508 1636 8560
rect 7564 8551 7616 8560
rect 7564 8517 7573 8551
rect 7573 8517 7607 8551
rect 7607 8517 7616 8551
rect 10692 8551 10744 8560
rect 7564 8508 7616 8517
rect 10692 8517 10701 8551
rect 10701 8517 10735 8551
rect 10735 8517 10744 8551
rect 10692 8508 10744 8517
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 14556 8576 14608 8628
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 19892 8619 19944 8628
rect 19892 8585 19901 8619
rect 19901 8585 19935 8619
rect 19935 8585 19944 8619
rect 19892 8576 19944 8585
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 21732 8619 21784 8628
rect 21732 8585 21741 8619
rect 21741 8585 21775 8619
rect 21775 8585 21784 8619
rect 21732 8576 21784 8585
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 12992 8508 13044 8560
rect 14648 8551 14700 8560
rect 2044 8440 2096 8492
rect 2964 8440 3016 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 7748 8440 7800 8492
rect 2320 8372 2372 8424
rect 12624 8440 12676 8492
rect 14648 8517 14657 8551
rect 14657 8517 14691 8551
rect 14691 8517 14700 8551
rect 14648 8508 14700 8517
rect 21456 8508 21508 8560
rect 18052 8440 18104 8492
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 21640 8440 21692 8492
rect 1492 8304 1544 8356
rect 2688 8304 2740 8356
rect 3424 8304 3476 8356
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 5448 8304 5500 8356
rect 4804 8236 4856 8245
rect 5356 8236 5408 8288
rect 6736 8304 6788 8356
rect 8576 8372 8628 8424
rect 9220 8347 9272 8356
rect 9220 8313 9229 8347
rect 9229 8313 9263 8347
rect 9263 8313 9272 8347
rect 9220 8304 9272 8313
rect 9956 8304 10008 8356
rect 10232 8347 10284 8356
rect 10232 8313 10241 8347
rect 10241 8313 10275 8347
rect 10275 8313 10284 8347
rect 10232 8304 10284 8313
rect 12992 8304 13044 8356
rect 14188 8304 14240 8356
rect 15384 8304 15436 8356
rect 15936 8304 15988 8356
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 13084 8236 13136 8288
rect 15660 8236 15712 8288
rect 22008 8372 22060 8424
rect 17316 8304 17368 8356
rect 19156 8304 19208 8356
rect 20904 8347 20956 8356
rect 20904 8313 20913 8347
rect 20913 8313 20947 8347
rect 20947 8313 20956 8347
rect 20904 8304 20956 8313
rect 21180 8304 21232 8356
rect 21640 8236 21692 8288
rect 22100 8279 22152 8288
rect 22100 8245 22109 8279
rect 22109 8245 22143 8279
rect 22143 8245 22152 8279
rect 22100 8236 22152 8245
rect 22192 8236 22244 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1676 8032 1728 8084
rect 3424 8032 3476 8084
rect 4620 8032 4672 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 7748 8032 7800 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 112 7964 164 8016
rect 3976 7964 4028 8016
rect 5356 7964 5408 8016
rect 6736 8007 6788 8016
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 6736 7973 6745 8007
rect 6745 7973 6779 8007
rect 6779 7973 6788 8007
rect 6736 7964 6788 7973
rect 9864 7964 9916 8016
rect 11060 8032 11112 8084
rect 12900 8032 12952 8084
rect 15292 8032 15344 8084
rect 15384 8032 15436 8084
rect 16488 8032 16540 8084
rect 16948 8032 17000 8084
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 21456 8032 21508 8084
rect 22836 8032 22888 8084
rect 10416 7964 10468 8016
rect 2504 7828 2556 7880
rect 7840 7896 7892 7948
rect 9036 7896 9088 7948
rect 9404 7896 9456 7948
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12072 7896 12124 7948
rect 12624 7896 12676 7948
rect 13636 7896 13688 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 6184 7828 6236 7880
rect 3884 7760 3936 7812
rect 7012 7828 7064 7880
rect 8484 7828 8536 7880
rect 12992 7828 13044 7880
rect 17316 7964 17368 8016
rect 17776 7964 17828 8016
rect 21088 8007 21140 8016
rect 21088 7973 21097 8007
rect 21097 7973 21131 8007
rect 21131 7973 21140 8007
rect 21088 7964 21140 7973
rect 21180 7964 21232 8016
rect 16304 7896 16356 7948
rect 18420 7896 18472 7948
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 21272 7828 21324 7880
rect 1768 7692 1820 7744
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 11612 7692 11664 7744
rect 14464 7692 14516 7744
rect 22008 7692 22060 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2964 7488 3016 7540
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 4804 7488 4856 7540
rect 6736 7488 6788 7540
rect 1676 7420 1728 7472
rect 2688 7420 2740 7472
rect 4160 7420 4212 7472
rect 7656 7488 7708 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 9588 7488 9640 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 9956 7420 10008 7472
rect 2136 7352 2188 7404
rect 3056 7352 3108 7404
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 1584 7284 1636 7336
rect 1860 7284 1912 7336
rect 4620 7284 4672 7336
rect 11520 7488 11572 7540
rect 11704 7488 11756 7540
rect 10416 7463 10468 7472
rect 10416 7429 10425 7463
rect 10425 7429 10459 7463
rect 10459 7429 10468 7463
rect 10416 7420 10468 7429
rect 11428 7420 11480 7472
rect 13636 7463 13688 7472
rect 13636 7429 13645 7463
rect 13645 7429 13679 7463
rect 13679 7429 13688 7463
rect 13636 7420 13688 7429
rect 11152 7352 11204 7404
rect 12072 7352 12124 7404
rect 12808 7352 12860 7404
rect 14096 7488 14148 7540
rect 14740 7488 14792 7540
rect 15384 7488 15436 7540
rect 15568 7488 15620 7540
rect 15752 7488 15804 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 18972 7531 19024 7540
rect 18972 7497 18981 7531
rect 18981 7497 19015 7531
rect 19015 7497 19024 7531
rect 18972 7488 19024 7497
rect 19156 7488 19208 7540
rect 21088 7488 21140 7540
rect 15476 7420 15528 7472
rect 16028 7420 16080 7472
rect 20904 7420 20956 7472
rect 18052 7395 18104 7404
rect 10048 7284 10100 7336
rect 14464 7284 14516 7336
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 19248 7352 19300 7404
rect 4988 7216 5040 7268
rect 6000 7216 6052 7268
rect 7932 7259 7984 7268
rect 7932 7225 7941 7259
rect 7941 7225 7975 7259
rect 7975 7225 7984 7259
rect 7932 7216 7984 7225
rect 5356 7191 5408 7200
rect 5356 7157 5365 7191
rect 5365 7157 5399 7191
rect 5399 7157 5408 7191
rect 5356 7148 5408 7157
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 8668 7216 8720 7268
rect 10784 7259 10836 7268
rect 10784 7225 10793 7259
rect 10793 7225 10827 7259
rect 10827 7225 10836 7259
rect 12624 7259 12676 7268
rect 10784 7216 10836 7225
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 15384 7259 15436 7268
rect 15384 7225 15393 7259
rect 15393 7225 15427 7259
rect 15427 7225 15436 7259
rect 15384 7216 15436 7225
rect 15568 7216 15620 7268
rect 19156 7216 19208 7268
rect 8208 7148 8260 7200
rect 9036 7148 9088 7200
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 12440 7148 12492 7200
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 18420 7148 18472 7200
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1492 6944 1544 6996
rect 2504 6987 2556 6996
rect 2504 6953 2513 6987
rect 2513 6953 2547 6987
rect 2547 6953 2556 6987
rect 2504 6944 2556 6953
rect 6920 6944 6972 6996
rect 8208 6987 8260 6996
rect 8208 6953 8217 6987
rect 8217 6953 8251 6987
rect 8251 6953 8260 6987
rect 8208 6944 8260 6953
rect 9864 6944 9916 6996
rect 1952 6876 2004 6928
rect 2780 6876 2832 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 3792 6808 3844 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 5540 6808 5592 6860
rect 5908 6808 5960 6860
rect 7840 6876 7892 6928
rect 10784 6944 10836 6996
rect 16764 6944 16816 6996
rect 19248 6944 19300 6996
rect 21272 6944 21324 6996
rect 11612 6919 11664 6928
rect 11612 6885 11621 6919
rect 11621 6885 11655 6919
rect 11655 6885 11664 6919
rect 11612 6876 11664 6885
rect 12624 6876 12676 6928
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 13820 6919 13872 6928
rect 13820 6885 13829 6919
rect 13829 6885 13863 6919
rect 13863 6885 13872 6919
rect 13820 6876 13872 6885
rect 15568 6876 15620 6928
rect 16028 6919 16080 6928
rect 16028 6885 16037 6919
rect 16037 6885 16071 6919
rect 16071 6885 16080 6919
rect 16028 6876 16080 6885
rect 20996 6876 21048 6928
rect 21732 6876 21784 6928
rect 7196 6808 7248 6860
rect 8576 6808 8628 6860
rect 9220 6808 9272 6860
rect 9864 6808 9916 6860
rect 4344 6740 4396 6792
rect 7380 6740 7432 6792
rect 11980 6740 12032 6792
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 17224 6808 17276 6860
rect 17776 6808 17828 6860
rect 18604 6851 18656 6860
rect 18604 6817 18613 6851
rect 18613 6817 18647 6851
rect 18647 6817 18656 6851
rect 18604 6808 18656 6817
rect 18972 6851 19024 6860
rect 18972 6817 18981 6851
rect 18981 6817 19015 6851
rect 19015 6817 19024 6851
rect 18972 6808 19024 6817
rect 20628 6808 20680 6860
rect 21640 6851 21692 6860
rect 21640 6817 21649 6851
rect 21649 6817 21683 6851
rect 21683 6817 21692 6851
rect 21640 6808 21692 6817
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 16396 6740 16448 6792
rect 21364 6740 21416 6792
rect 22192 6740 22244 6792
rect 8852 6672 8904 6724
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 15660 6672 15712 6724
rect 11152 6604 11204 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 15384 6604 15436 6656
rect 15844 6604 15896 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3148 6400 3200 6452
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 5540 6332 5592 6384
rect 7472 6332 7524 6384
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 8208 6400 8260 6452
rect 8944 6400 8996 6452
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 10784 6400 10836 6452
rect 11612 6443 11664 6452
rect 11612 6409 11621 6443
rect 11621 6409 11655 6443
rect 11655 6409 11664 6443
rect 11612 6400 11664 6409
rect 13820 6400 13872 6452
rect 17132 6400 17184 6452
rect 19064 6400 19116 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 8116 6332 8168 6384
rect 8668 6332 8720 6384
rect 12072 6332 12124 6384
rect 17224 6332 17276 6384
rect 17316 6332 17368 6384
rect 19984 6332 20036 6384
rect 8300 6264 8352 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 11428 6264 11480 6316
rect 19524 6264 19576 6316
rect 21180 6264 21232 6316
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2780 6060 2832 6112
rect 3516 6171 3568 6180
rect 3516 6137 3525 6171
rect 3525 6137 3559 6171
rect 3559 6137 3568 6171
rect 3516 6128 3568 6137
rect 5356 6128 5408 6180
rect 7196 6196 7248 6248
rect 7748 6196 7800 6248
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 18604 6196 18656 6248
rect 8024 6128 8076 6180
rect 8944 6171 8996 6180
rect 8944 6137 8953 6171
rect 8953 6137 8987 6171
rect 8987 6137 8996 6171
rect 8944 6128 8996 6137
rect 10048 6128 10100 6180
rect 10784 6128 10836 6180
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 7840 6103 7892 6112
rect 7840 6069 7849 6103
rect 7849 6069 7883 6103
rect 7883 6069 7892 6103
rect 7840 6060 7892 6069
rect 9772 6060 9824 6112
rect 13360 6128 13412 6180
rect 19984 6171 20036 6180
rect 19984 6137 19993 6171
rect 19993 6137 20027 6171
rect 20027 6137 20036 6171
rect 19984 6128 20036 6137
rect 11980 6103 12032 6112
rect 11980 6069 11989 6103
rect 11989 6069 12023 6103
rect 12023 6069 12032 6103
rect 11980 6060 12032 6069
rect 15568 6060 15620 6112
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 10876 5856 10928 5908
rect 12624 5856 12676 5908
rect 14096 5856 14148 5908
rect 18052 5856 18104 5908
rect 19524 5856 19576 5908
rect 4160 5788 4212 5840
rect 5264 5788 5316 5840
rect 6368 5788 6420 5840
rect 8208 5831 8260 5840
rect 8208 5797 8217 5831
rect 8217 5797 8251 5831
rect 8251 5797 8260 5831
rect 8208 5788 8260 5797
rect 10692 5831 10744 5840
rect 10692 5797 10701 5831
rect 10701 5797 10735 5831
rect 10735 5797 10744 5831
rect 10692 5788 10744 5797
rect 13360 5788 13412 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 17040 5831 17092 5840
rect 17040 5797 17049 5831
rect 17049 5797 17083 5831
rect 17083 5797 17092 5831
rect 17040 5788 17092 5797
rect 3516 5720 3568 5772
rect 12164 5720 12216 5772
rect 18328 5720 18380 5772
rect 18972 5763 19024 5772
rect 18972 5729 18981 5763
rect 18981 5729 19015 5763
rect 19015 5729 19024 5763
rect 18972 5720 19024 5729
rect 21180 5720 21232 5772
rect 23848 5720 23900 5772
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 6460 5652 6512 5704
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 11428 5652 11480 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 11244 5584 11296 5636
rect 15936 5584 15988 5636
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 10048 5516 10100 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 24216 5516 24268 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4528 5312 4580 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 6644 5244 6696 5296
rect 5448 5040 5500 5092
rect 9772 5312 9824 5364
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 11428 5355 11480 5364
rect 11428 5321 11437 5355
rect 11437 5321 11471 5355
rect 11471 5321 11480 5355
rect 11428 5312 11480 5321
rect 12164 5355 12216 5364
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 13360 5312 13412 5364
rect 12992 5219 13044 5228
rect 9956 5108 10008 5160
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 12624 5108 12676 5160
rect 13544 5108 13596 5160
rect 14372 5312 14424 5364
rect 15476 5312 15528 5364
rect 15568 5312 15620 5364
rect 17040 5312 17092 5364
rect 18328 5312 18380 5364
rect 19156 5312 19208 5364
rect 22376 5312 22428 5364
rect 23848 5355 23900 5364
rect 23848 5321 23857 5355
rect 23857 5321 23891 5355
rect 23891 5321 23900 5355
rect 23848 5312 23900 5321
rect 14280 5244 14332 5296
rect 15660 5244 15712 5296
rect 16028 5176 16080 5228
rect 16948 5176 17000 5228
rect 14004 5151 14056 5160
rect 14004 5117 14013 5151
rect 14013 5117 14047 5151
rect 14047 5117 14056 5151
rect 14004 5108 14056 5117
rect 2320 4972 2372 5024
rect 4160 4972 4212 5024
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 19156 5108 19208 5160
rect 24216 5108 24268 5160
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 27344 4972 27396 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5448 4768 5500 4820
rect 8208 4768 8260 4820
rect 8668 4768 8720 4820
rect 12808 4768 12860 4820
rect 13176 4768 13228 4820
rect 13452 4768 13504 4820
rect 7840 4700 7892 4752
rect 8024 4700 8076 4752
rect 8852 4700 8904 4752
rect 9496 4700 9548 4752
rect 11428 4700 11480 4752
rect 12440 4700 12492 4752
rect 14004 4768 14056 4820
rect 15384 4768 15436 4820
rect 16028 4768 16080 4820
rect 16396 4768 16448 4820
rect 18972 4768 19024 4820
rect 15568 4700 15620 4752
rect 2872 4632 2924 4684
rect 4712 4675 4764 4684
rect 4712 4641 4730 4675
rect 4730 4641 4764 4675
rect 4712 4632 4764 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 12164 4675 12216 4684
rect 12164 4641 12182 4675
rect 12182 4641 12216 4675
rect 12164 4632 12216 4641
rect 13084 4632 13136 4684
rect 13544 4675 13596 4684
rect 6000 4564 6052 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 10692 4564 10744 4616
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 15384 4607 15436 4616
rect 6460 4496 6512 4548
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 13728 4496 13780 4548
rect 6000 4428 6052 4480
rect 13268 4428 13320 4480
rect 13452 4428 13504 4480
rect 18604 4428 18656 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 6092 4267 6144 4276
rect 6092 4233 6101 4267
rect 6101 4233 6135 4267
rect 6135 4233 6144 4267
rect 6092 4224 6144 4233
rect 6552 4224 6604 4276
rect 7840 4224 7892 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 11244 4267 11296 4276
rect 4712 4199 4764 4208
rect 4712 4165 4721 4199
rect 4721 4165 4755 4199
rect 4755 4165 4764 4199
rect 4712 4156 4764 4165
rect 5540 4156 5592 4208
rect 6000 4156 6052 4208
rect 8024 4156 8076 4208
rect 8668 4156 8720 4208
rect 7380 4063 7432 4072
rect 7380 4029 7389 4063
rect 7389 4029 7423 4063
rect 7423 4029 7432 4063
rect 7380 4020 7432 4029
rect 8208 3995 8260 4004
rect 8208 3961 8217 3995
rect 8217 3961 8251 3995
rect 8251 3961 8260 3995
rect 8208 3952 8260 3961
rect 8300 3995 8352 4004
rect 8300 3961 8309 3995
rect 8309 3961 8343 3995
rect 8343 3961 8352 3995
rect 9496 4020 9548 4072
rect 8300 3952 8352 3961
rect 11244 4233 11253 4267
rect 11253 4233 11287 4267
rect 11287 4233 11296 4267
rect 11244 4224 11296 4233
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 13452 4224 13504 4276
rect 13544 4224 13596 4276
rect 14832 4224 14884 4276
rect 15476 4224 15528 4276
rect 15844 4224 15896 4276
rect 14556 4156 14608 4208
rect 14740 4088 14792 4140
rect 11520 4020 11572 4072
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 14464 4020 14516 4072
rect 15568 4156 15620 4208
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 19156 4088 19208 4140
rect 20720 4088 20772 4140
rect 19064 4020 19116 4072
rect 22008 4020 22060 4072
rect 17316 3952 17368 4004
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 12624 3884 12676 3936
rect 16856 3884 16908 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 7472 3723 7524 3732
rect 7472 3689 7481 3723
rect 7481 3689 7515 3723
rect 7515 3689 7524 3723
rect 7472 3680 7524 3689
rect 8208 3680 8260 3732
rect 10692 3680 10744 3732
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 13360 3680 13412 3732
rect 8300 3612 8352 3664
rect 9496 3612 9548 3664
rect 13452 3612 13504 3664
rect 15384 3680 15436 3732
rect 19984 3680 20036 3732
rect 7656 3587 7708 3596
rect 7656 3553 7665 3587
rect 7665 3553 7699 3587
rect 7699 3553 7708 3587
rect 7656 3544 7708 3553
rect 7748 3544 7800 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 18420 3612 18472 3664
rect 13912 3544 13964 3596
rect 16856 3544 16908 3596
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 10140 3383 10192 3392
rect 10140 3349 10149 3383
rect 10149 3349 10183 3383
rect 10183 3349 10192 3383
rect 10140 3340 10192 3349
rect 11428 3383 11480 3392
rect 11428 3349 11437 3383
rect 11437 3349 11471 3383
rect 11471 3349 11480 3383
rect 11428 3340 11480 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 6552 3179 6604 3188
rect 6552 3145 6561 3179
rect 6561 3145 6595 3179
rect 6595 3145 6604 3179
rect 6552 3136 6604 3145
rect 7932 3136 7984 3188
rect 11152 3136 11204 3188
rect 11980 3136 12032 3188
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 14280 3179 14332 3188
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 19708 3179 19760 3188
rect 19708 3145 19717 3179
rect 19717 3145 19751 3179
rect 19751 3145 19760 3179
rect 19708 3136 19760 3145
rect 11244 3068 11296 3120
rect 22008 3068 22060 3120
rect 27620 3068 27672 3120
rect 7656 3000 7708 3052
rect 10140 3000 10192 3052
rect 3976 2932 4028 2984
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 11704 2932 11756 2984
rect 12532 2932 12584 2984
rect 13728 3000 13780 3052
rect 14280 2932 14332 2984
rect 19340 2932 19392 2984
rect 12624 2864 12676 2916
rect 24032 2932 24084 2984
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 18144 2796 18196 2848
rect 19156 2796 19208 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 6184 2592 6236 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 10048 2592 10100 2644
rect 12900 2592 12952 2644
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 4712 2456 4764 2508
rect 11336 2524 11388 2576
rect 7840 2456 7892 2508
rect 9312 2456 9364 2508
rect 19156 2499 19208 2508
rect 6276 2388 6328 2440
rect 19156 2465 19165 2499
rect 19165 2465 19199 2499
rect 19199 2465 19208 2499
rect 19156 2456 19208 2465
rect 21456 2456 21508 2508
rect 10048 2320 10100 2372
rect 16856 2320 16908 2372
rect 27620 2320 27672 2372
rect 4712 2295 4764 2304
rect 4712 2261 4721 2295
rect 4721 2261 4755 2295
rect 4755 2261 4764 2295
rect 4712 2252 4764 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 17776 2252 17828 2304
rect 23020 2252 23072 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 664 76 716 128
rect 1308 76 1360 128
<< metal2 >>
rect 478 27520 534 28000
rect 1398 27520 1454 28000
rect 1964 27526 2360 27554
rect 110 25800 166 25809
rect 110 25735 166 25744
rect 124 24138 152 25735
rect 112 24132 164 24138
rect 112 24074 164 24080
rect 110 22808 166 22817
rect 110 22743 166 22752
rect 124 22710 152 22743
rect 112 22704 164 22710
rect 112 22646 164 22652
rect 492 20602 520 27520
rect 1122 26752 1178 26761
rect 1122 26687 1178 26696
rect 1136 23662 1164 26687
rect 1124 23656 1176 23662
rect 1124 23598 1176 23604
rect 480 20596 532 20602
rect 480 20538 532 20544
rect 1412 20330 1440 27520
rect 1582 24032 1638 24041
rect 1582 23967 1638 23976
rect 1596 22778 1624 23967
rect 1964 23474 1992 27526
rect 2332 27520 2360 27526
rect 2410 27520 2466 28000
rect 3422 27554 3478 28000
rect 3068 27526 3478 27554
rect 2332 27492 2452 27520
rect 3068 23474 3096 27526
rect 3422 27520 3478 27526
rect 4434 27554 4490 28000
rect 4434 27526 4752 27554
rect 4434 27520 4490 27526
rect 4436 27124 4488 27130
rect 4436 27066 4488 27072
rect 3792 23588 3844 23594
rect 3792 23530 3844 23536
rect 1872 23446 1992 23474
rect 2976 23446 3096 23474
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1492 22432 1544 22438
rect 1492 22374 1544 22380
rect 1400 20324 1452 20330
rect 1400 20266 1452 20272
rect 1504 19922 1532 22374
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 110 19816 166 19825
rect 110 19751 166 19760
rect 124 18970 152 19751
rect 112 18964 164 18970
rect 112 18906 164 18912
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 17270 1440 18702
rect 1504 18630 1532 19858
rect 1780 19514 1808 20334
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1400 17264 1452 17270
rect 1400 17206 1452 17212
rect 1688 17202 1716 17682
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 112 15904 164 15910
rect 112 15846 164 15852
rect 124 12481 152 15846
rect 1688 13530 1716 16050
rect 1872 15162 1900 23446
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2700 22642 2728 22918
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2700 22234 2728 22578
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 1950 21176 2006 21185
rect 2240 21146 2268 21286
rect 1950 21111 2006 21120
rect 2228 21140 2280 21146
rect 1964 21078 1992 21111
rect 2228 21082 2280 21088
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1964 20058 1992 20266
rect 2148 20058 2176 20742
rect 2240 20398 2268 21082
rect 2516 21010 2544 21830
rect 2700 21350 2728 22034
rect 2884 21690 2912 22034
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2872 21480 2924 21486
rect 2872 21422 2924 21428
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2700 21049 2728 21286
rect 2686 21040 2742 21049
rect 2412 21004 2464 21010
rect 2412 20946 2464 20952
rect 2504 21004 2556 21010
rect 2686 20975 2742 20984
rect 2504 20946 2556 20952
rect 2424 20602 2452 20946
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2240 19854 2268 20334
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 19922 2452 20198
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2044 19780 2096 19786
rect 2044 19722 2096 19728
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1964 17610 1992 19654
rect 2056 18358 2084 19722
rect 2240 18698 2268 19790
rect 2424 19446 2452 19858
rect 2516 19700 2544 20946
rect 2700 20874 2728 20975
rect 2688 20868 2740 20874
rect 2688 20810 2740 20816
rect 2596 19712 2648 19718
rect 2516 19672 2596 19700
rect 2596 19654 2648 19660
rect 2412 19440 2464 19446
rect 2412 19382 2464 19388
rect 2424 18834 2452 19382
rect 2700 19334 2728 20810
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2792 19446 2820 19722
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 2700 19306 2820 19334
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2044 18352 2096 18358
rect 2044 18294 2096 18300
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 2056 17542 2084 17614
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 17134 2084 17478
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1964 16590 1992 17070
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1964 16250 1992 16526
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2056 15162 2084 17070
rect 2148 16153 2176 18566
rect 2424 17796 2452 18770
rect 2608 18426 2636 18838
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2700 18698 2728 18770
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2504 17808 2556 17814
rect 2424 17768 2504 17796
rect 2504 17750 2556 17756
rect 2688 17740 2740 17746
rect 2792 17728 2820 19306
rect 2884 18766 2912 21422
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2740 17700 2820 17728
rect 2688 17682 2740 17688
rect 2700 16998 2728 17682
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2884 16658 2912 18702
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2504 16584 2556 16590
rect 2976 16538 3004 23446
rect 3804 23118 3832 23530
rect 4344 23520 4396 23526
rect 4344 23462 4396 23468
rect 4252 23248 4304 23254
rect 4252 23190 4304 23196
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 4264 22778 4292 23190
rect 4356 22778 4384 23462
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4356 22506 4384 22714
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4172 22166 4200 22442
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 21554 3648 21830
rect 4172 21690 4200 22102
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3790 20496 3846 20505
rect 3790 20431 3846 20440
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 3712 19786 3740 20334
rect 3804 19922 3832 20431
rect 3896 20398 3924 20878
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3896 19990 3924 20334
rect 4080 20262 4108 20946
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4172 20602 4200 20810
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4172 20330 4200 20538
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 4080 19922 4108 20198
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3700 19780 3752 19786
rect 3700 19722 3752 19728
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3712 18834 3740 19246
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18086 3280 18566
rect 3344 18426 3372 18702
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3146 17640 3202 17649
rect 3146 17575 3202 17584
rect 2504 16526 2556 16532
rect 2134 16144 2190 16153
rect 2134 16079 2190 16088
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1872 14618 1900 15098
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 110 12472 166 12481
rect 110 12407 166 12416
rect 1308 11212 1360 11218
rect 1308 11154 1360 11160
rect 110 10976 166 10985
rect 110 10911 166 10920
rect 124 9042 152 10911
rect 1320 10470 1348 11154
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1308 10464 1360 10470
rect 1308 10406 1360 10412
rect 112 9036 164 9042
rect 112 8978 164 8984
rect 110 8120 166 8129
rect 110 8055 166 8064
rect 124 8022 152 8055
rect 112 8016 164 8022
rect 112 7958 164 7964
rect 662 128 718 480
rect 1320 134 1348 10406
rect 1490 9752 1546 9761
rect 1490 9687 1546 9696
rect 1504 9625 1532 9687
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1504 9518 1532 9551
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1596 8566 1624 11018
rect 1688 10606 1716 12582
rect 1872 12102 1900 12718
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 10690 1900 12038
rect 1964 11898 1992 13466
rect 2056 12306 2084 14826
rect 2134 14648 2190 14657
rect 2240 14618 2268 15506
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 14958 2360 15302
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2134 14583 2190 14592
rect 2228 14612 2280 14618
rect 2148 14482 2176 14583
rect 2228 14554 2280 14560
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2148 13530 2176 14418
rect 2332 14346 2360 14894
rect 2228 14340 2280 14346
rect 2228 14282 2280 14288
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2136 13388 2188 13394
rect 2240 13376 2268 14282
rect 2424 13802 2452 14894
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2188 13348 2268 13376
rect 2136 13330 2188 13336
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2056 11898 2084 12242
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1964 11694 1992 11834
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2056 11370 2084 11834
rect 1964 11342 2084 11370
rect 1964 10810 1992 11342
rect 2042 11248 2098 11257
rect 2042 11183 2098 11192
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1872 10662 1992 10690
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1688 10266 1716 10542
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 7002 1532 8298
rect 1688 8090 1716 10202
rect 1872 9926 1900 10542
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1688 7478 1716 8026
rect 1780 7750 1808 8978
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1596 6866 1624 7278
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6118 1624 6802
rect 1780 6225 1808 7686
rect 1872 7342 1900 9862
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1964 6934 1992 10662
rect 2056 10130 2084 11183
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2056 9722 2084 10066
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 8838 2084 9454
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8498 2084 8774
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2148 7410 2176 13330
rect 2424 13258 2452 13738
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12918 2360 13126
rect 2320 12912 2372 12918
rect 2320 12854 2372 12860
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 12102 2268 12582
rect 2332 12102 2360 12854
rect 2424 12170 2452 13194
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2240 11830 2268 12038
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2240 9518 2268 11766
rect 2332 11762 2360 12038
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11150 2360 11698
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2226 9344 2282 9353
rect 2226 9279 2282 9288
rect 2240 8634 2268 9279
rect 2332 8838 2360 11086
rect 2424 11082 2452 12106
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2516 10130 2544 16526
rect 2884 16510 3004 16538
rect 2884 16250 2912 16510
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2884 16046 2912 16186
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15502 2912 15982
rect 2976 15502 3004 16390
rect 2872 15496 2924 15502
rect 2792 15456 2872 15484
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 15094 2728 15302
rect 2792 15162 2820 15456
rect 2872 15438 2924 15444
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2424 9625 2452 9658
rect 2410 9616 2466 9625
rect 2410 9551 2466 9560
rect 2608 9518 2636 14554
rect 2700 14278 2728 15030
rect 2976 15008 3004 15438
rect 2792 14980 3004 15008
rect 2792 14890 2820 14980
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2872 14884 2924 14890
rect 3068 14872 3096 16390
rect 3160 15638 3188 17575
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 2924 14844 3096 14872
rect 2872 14826 2924 14832
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 14074 2728 14214
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2700 12986 2728 14010
rect 3068 13802 3096 14844
rect 3160 14346 3188 15030
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2792 11744 2820 13670
rect 3068 13394 3096 13738
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3068 12764 3096 13330
rect 3148 12776 3200 12782
rect 3068 12736 3148 12764
rect 3148 12718 3200 12724
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2700 11716 2820 11744
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2516 9178 2544 9454
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2504 8968 2556 8974
rect 2608 8956 2636 9318
rect 2700 9042 2728 11716
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2556 8928 2636 8956
rect 2504 8910 2556 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2332 8430 2360 8774
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2516 7886 2544 8910
rect 2700 8362 2728 8978
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2516 7002 2544 7822
rect 2700 7478 2728 7890
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2792 6934 2820 11562
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10470 2912 11154
rect 2976 10656 3004 12038
rect 3056 10668 3108 10674
rect 2976 10628 3056 10656
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 1964 6118 1992 6870
rect 2792 6118 2820 6870
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 1596 1329 1624 6054
rect 1964 2689 1992 6054
rect 2792 5914 2820 6054
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1950 2680 2006 2689
rect 1950 2615 2006 2624
rect 1582 1320 1638 1329
rect 1582 1255 1638 1264
rect 662 76 664 128
rect 716 76 718 128
rect 662 0 718 76
rect 1308 128 1360 134
rect 1308 70 1360 76
rect 1950 82 2006 480
rect 2332 82 2360 4966
rect 2884 4690 2912 10406
rect 2976 10130 3004 10628
rect 3056 10610 3108 10616
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10266 3096 10474
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 9382 3004 10066
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2976 8498 3004 8842
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 7546 3004 8434
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3068 7410 3096 10202
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3160 9042 3188 10134
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3160 6458 3188 8978
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3160 6361 3188 6394
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 3252 4154 3280 18022
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3436 14958 3464 15302
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3528 14482 3556 15914
rect 3516 14476 3568 14482
rect 3436 14436 3516 14464
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3344 12714 3372 13330
rect 3436 13326 3464 14436
rect 3516 14418 3568 14424
rect 3620 14362 3648 16934
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15570 3740 15846
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3528 14334 3648 14362
rect 3528 13734 3556 14334
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3620 13530 3648 13874
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3712 13394 3740 15506
rect 3804 15094 3832 19858
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3988 19145 4016 19450
rect 4172 19242 4200 19654
rect 4264 19514 4292 20266
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4356 19310 4384 19858
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 3974 19136 4030 19145
rect 3974 19071 4030 19080
rect 4172 18884 4200 19178
rect 4252 18896 4304 18902
rect 4172 18856 4252 18884
rect 4448 18873 4476 27066
rect 4724 24342 4752 27526
rect 5446 27520 5502 28000
rect 6458 27520 6514 28000
rect 7470 27520 7526 28000
rect 8390 27520 8446 28000
rect 9402 27520 9458 28000
rect 10414 27554 10470 28000
rect 10152 27526 10470 27554
rect 5460 27130 5488 27520
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4540 22778 4568 23054
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4252 18838 4304 18844
rect 4434 18864 4490 18873
rect 4908 18834 4936 23462
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 5184 22506 5212 23122
rect 5172 22500 5224 22506
rect 5172 22442 5224 22448
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 5000 22234 5028 22374
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5184 22098 5212 22442
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 5000 21350 5028 21422
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 5000 20505 5028 21286
rect 4986 20496 5042 20505
rect 4986 20431 5042 20440
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 5184 19718 5212 20334
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4434 18799 4490 18808
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 5000 18630 5028 19178
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3884 18352 3936 18358
rect 3884 18294 3936 18300
rect 3896 18154 3924 18294
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3896 17882 3924 18090
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3988 17202 4016 18362
rect 4160 18148 4212 18154
rect 4160 18090 4212 18096
rect 4172 17882 4200 18090
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4264 17814 4292 18022
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3882 16688 3938 16697
rect 3882 16623 3938 16632
rect 3896 16590 3924 16623
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3896 15162 3924 16526
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 14278 3924 14758
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14074 3924 14214
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3804 13433 3832 13738
rect 3790 13424 3846 13433
rect 3700 13388 3752 13394
rect 3790 13359 3846 13368
rect 3700 13330 3752 13336
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3436 12850 3464 13262
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3792 13184 3844 13190
rect 3896 13172 3924 14010
rect 3988 13814 4016 17138
rect 4080 16658 4108 17478
rect 4264 16658 4292 17546
rect 4448 16998 4476 17750
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16794 4476 16934
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 15570 4108 16458
rect 4250 16416 4306 16425
rect 4250 16351 4306 16360
rect 4264 15706 4292 16351
rect 4448 16250 4476 16730
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 4632 15978 4660 16730
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4724 15978 4752 16458
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 4080 15065 4108 15506
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 15366 4660 15438
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4172 14414 4200 14962
rect 4264 14822 4292 15302
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4172 13938 4200 14350
rect 4264 14278 4292 14758
rect 4632 14482 4660 15302
rect 5000 14618 5028 18566
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17134 5120 17478
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5080 15564 5132 15570
rect 5184 15552 5212 19654
rect 5368 18426 5396 23530
rect 5552 23322 5580 23598
rect 6196 23526 6224 24210
rect 6472 23866 6500 27520
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 5540 23316 5592 23322
rect 5540 23258 5592 23264
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6656 22642 6684 23122
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5552 21418 5580 21830
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21554 6040 21966
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5724 21412 5776 21418
rect 5724 21354 5776 21360
rect 5552 20806 5580 21354
rect 5736 21010 5764 21354
rect 5724 21004 5776 21010
rect 5724 20946 5776 20952
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 20398 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5460 19145 5488 19246
rect 5552 19242 5580 20334
rect 6012 20262 6040 20946
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6104 19514 6132 19790
rect 6092 19508 6144 19514
rect 6012 19468 6092 19496
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5446 19136 5502 19145
rect 5446 19071 5502 19080
rect 5460 18766 5488 19071
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5276 17184 5304 18090
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17882 5396 18022
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5460 17338 5488 18566
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18136 6040 19468
rect 6092 19450 6144 19456
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5920 18108 6040 18136
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 17196 5408 17202
rect 5276 17156 5356 17184
rect 5276 16726 5304 17156
rect 5356 17138 5408 17144
rect 5460 17066 5488 17274
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5552 16794 5580 18022
rect 5920 17524 5948 18108
rect 6104 18086 6132 18770
rect 6092 18080 6144 18086
rect 5998 18048 6054 18057
rect 6092 18022 6144 18028
rect 5998 17983 6054 17992
rect 6012 17882 6040 17983
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5920 17496 6040 17524
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 6012 16658 6040 17496
rect 6104 17105 6132 18022
rect 6090 17096 6146 17105
rect 6090 17031 6146 17040
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16182 6040 16594
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5132 15524 5212 15552
rect 5080 15506 5132 15512
rect 5092 15366 5120 15506
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 3988 13786 4108 13814
rect 3844 13144 3924 13172
rect 3792 13126 3844 13132
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3344 12102 3372 12650
rect 3436 12238 3464 12786
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11014 3372 12038
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 8634 3372 10950
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 10198 3464 10746
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8362 3464 9318
rect 3528 8945 3556 13126
rect 3804 12918 3832 13126
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 4080 12306 4108 13786
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3976 11892 4028 11898
rect 4080 11880 4108 12242
rect 4028 11852 4108 11880
rect 3976 11834 4028 11840
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 11354 3832 11630
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3804 11082 3832 11290
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3700 10532 3752 10538
rect 3700 10474 3752 10480
rect 3514 8936 3570 8945
rect 3712 8906 3740 10474
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3514 8871 3570 8880
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 3712 8498 3740 8842
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3436 8090 3464 8298
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3896 7818 3924 8910
rect 3988 8022 4016 11834
rect 4172 11082 4200 13330
rect 4448 13326 4476 13874
rect 4540 13734 4568 14282
rect 5092 13841 5120 15302
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5184 14618 5212 14894
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5078 13832 5134 13841
rect 5078 13767 5134 13776
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4448 12986 4476 13262
rect 4540 13258 4568 13670
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4540 12986 4568 13194
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4632 12918 4660 13194
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4632 12442 4660 12854
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4356 11762 4384 12174
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 11218 4384 11290
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 7546 3924 7754
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3528 5778 3556 6122
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 1950 54 2360 82
rect 3160 4126 3280 4154
rect 3160 82 3188 4126
rect 3988 2990 4016 7958
rect 4172 7478 4200 11018
rect 4356 10810 4384 11154
rect 4448 11082 4476 12378
rect 4724 11665 4752 13126
rect 5000 12782 5028 13126
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4710 11656 4766 11665
rect 4710 11591 4766 11600
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4632 10674 4660 11154
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4264 9586 4292 10066
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4264 6866 4292 8230
rect 4632 8090 4660 10610
rect 4724 10062 4752 11086
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9722 4752 9998
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4724 8634 4752 9046
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4816 8294 4844 9386
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4632 7342 4660 8026
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7546 4844 7822
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4908 7410 4936 8434
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 5000 7274 5028 12718
rect 5092 10810 5120 13767
rect 5184 13190 5212 14554
rect 5276 13462 5304 15914
rect 6000 15904 6052 15910
rect 6104 15892 6132 16594
rect 6052 15864 6132 15892
rect 6000 15846 6052 15852
rect 6012 15570 6040 15846
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 14958 6040 15506
rect 5448 14952 5500 14958
rect 6000 14952 6052 14958
rect 5448 14894 5500 14900
rect 5814 14920 5870 14929
rect 5460 14482 5488 14894
rect 6000 14894 6052 14900
rect 5814 14855 5870 14864
rect 5828 14618 5856 14855
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5368 13938 5396 14350
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 14006 6040 14418
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 6196 13814 6224 22578
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6472 21350 6500 22102
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6288 20466 6316 20742
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6472 20330 6500 21286
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6288 19417 6316 20198
rect 6472 19990 6500 20266
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6274 19408 6330 19417
rect 6274 19343 6330 19352
rect 6380 19310 6408 19790
rect 6472 19446 6500 19926
rect 6460 19440 6512 19446
rect 6460 19382 6512 19388
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6288 18068 6316 19110
rect 6380 18970 6408 19246
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6368 18080 6420 18086
rect 6288 18040 6368 18068
rect 6368 18022 6420 18028
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 16998 6316 17682
rect 6380 17678 6408 18022
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6380 17549 6408 17614
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6288 16017 6316 16934
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6274 16008 6330 16017
rect 6274 15943 6330 15952
rect 6656 14482 6684 16526
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 14074 6592 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5276 12850 5304 13398
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5368 12374 5396 13194
rect 5460 12782 5488 13806
rect 6000 13796 6052 13802
rect 6196 13786 6316 13814
rect 6000 13738 6052 13744
rect 6012 13326 6040 13738
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13462 6224 13670
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6090 13288 6146 13297
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 6012 12306 6040 13262
rect 6090 13223 6146 13232
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6104 12186 6132 13223
rect 6196 12986 6224 13398
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6012 12158 6132 12186
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 11354 5580 11630
rect 5540 11348 5592 11354
rect 5460 11308 5540 11336
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 5092 10606 5120 10746
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9654 5212 10406
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5460 8362 5488 11308
rect 5540 11290 5592 11296
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10674 5580 10950
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5552 9450 5580 10134
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 9110 5580 9386
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 8022 5396 8230
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5368 7206 5396 7958
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7392 6040 12158
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11626 6132 12038
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6104 9042 6132 10474
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8090 6132 8978
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 5920 7364 6040 7392
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5846 4200 6054
rect 4264 5914 4292 6802
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 6322 4384 6734
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 5368 6186 5396 7142
rect 5920 6866 5948 7364
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5552 6390 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 5276 5846 5304 6054
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 4172 5030 4200 5782
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 5370 4568 5646
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 5460 5098 5488 5510
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 5460 4826 5488 5034
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4724 4214 4752 4626
rect 6012 4622 6040 7210
rect 6196 7206 6224 7822
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4486 6040 4558
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4214 6040 4422
rect 6104 4282 6132 4626
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4724 2310 4752 2450
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 3238 82 3294 480
rect 3160 54 3294 82
rect 1950 0 2006 54
rect 3238 0 3294 54
rect 4618 82 4674 480
rect 4724 82 4752 2246
rect 4618 54 4752 82
rect 5552 82 5580 4150
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6196 2650 6224 7142
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6288 2446 6316 13786
rect 6564 12918 6592 14010
rect 6748 14006 6776 24278
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6840 22234 6868 22374
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6932 19334 6960 24006
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7392 22642 7420 22918
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7024 20602 7052 21014
rect 7392 20806 7420 22578
rect 7484 21185 7512 27520
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7564 24268 7616 24274
rect 7564 24210 7616 24216
rect 7576 23798 7604 24210
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7576 22098 7604 22442
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7470 21176 7526 21185
rect 7470 21111 7526 21120
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7116 19378 7144 19994
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7104 19372 7156 19378
rect 6932 19306 7052 19334
rect 7104 19314 7156 19320
rect 7024 18766 7052 19306
rect 7208 19242 7236 19654
rect 7392 19378 7420 20742
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7208 18902 7236 19178
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7484 18766 7512 21111
rect 7576 21078 7604 22034
rect 7760 21894 7788 22918
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7668 20942 7696 21558
rect 7760 21486 7788 21830
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7668 19718 7696 20878
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 18970 7696 19654
rect 7852 18986 7880 24006
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8036 22438 8064 23122
rect 8220 22982 8248 23122
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7944 21554 7972 21966
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7944 21146 7972 21490
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7852 18970 7972 18986
rect 7656 18964 7708 18970
rect 7852 18964 7984 18970
rect 7852 18958 7932 18964
rect 7656 18906 7708 18912
rect 7932 18906 7984 18912
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7024 18630 7052 18702
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6920 18216 6972 18222
rect 6840 18176 6920 18204
rect 6840 17542 6868 18176
rect 6920 18158 6972 18164
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17746 7144 18022
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6840 16658 6868 17478
rect 7484 17066 7512 17818
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7024 16454 7052 16934
rect 7668 16658 7696 18634
rect 7852 18426 7880 18838
rect 7932 18692 7984 18698
rect 7932 18634 7984 18640
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7944 18306 7972 18634
rect 7852 18278 7972 18306
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7760 16794 7788 17070
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7668 16454 7696 16594
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7024 15910 7052 16390
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15706 7052 15846
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7024 14822 7052 15642
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14550 7052 14758
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 12102 6408 12718
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11898 6408 12038
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6380 11286 6408 11562
rect 6472 11286 6500 12174
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6380 9926 6408 11222
rect 6656 11014 6684 11494
rect 6748 11257 6776 13942
rect 7024 13734 7052 14486
rect 7668 14414 7696 16390
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7116 13870 7144 13942
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7116 13394 7144 13806
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12238 6960 12582
rect 7116 12374 7144 12922
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11898 6960 12174
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7116 11626 7144 12310
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 6734 11248 6790 11257
rect 6734 11183 6790 11192
rect 6644 11008 6696 11014
rect 7012 11008 7064 11014
rect 6644 10950 6696 10956
rect 6932 10968 7012 10996
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10266 6592 10406
rect 6460 10260 6512 10266
rect 6552 10260 6604 10266
rect 6512 10220 6552 10248
rect 6460 10202 6512 10208
rect 6552 10202 6604 10208
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6472 9722 6500 10202
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6656 9110 6684 10950
rect 6932 10538 6960 10968
rect 7012 10950 7064 10956
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6840 9926 6868 10134
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9110 6868 9522
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6748 8022 6776 8298
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6748 7546 6776 7958
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6932 7002 6960 10474
rect 7208 10130 7236 14350
rect 7760 13546 7788 16458
rect 7852 13734 7880 18278
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7944 17338 7972 18090
rect 8036 17678 8064 22374
rect 8312 20913 8340 24686
rect 8404 23866 8432 27520
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8588 22642 8616 23054
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8760 22500 8812 22506
rect 8760 22442 8812 22448
rect 8668 22160 8720 22166
rect 8772 22148 8800 22442
rect 9048 22234 9076 24550
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 9140 23322 9168 23462
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 8720 22120 8800 22148
rect 8668 22102 8720 22108
rect 8772 21486 8800 22120
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 8864 21690 8892 22034
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8298 20904 8354 20913
rect 8298 20839 8354 20848
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8220 17338 8248 19790
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8312 16522 8340 20839
rect 8588 20602 8616 20946
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8496 18290 8524 18906
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8588 17202 8616 19382
rect 8680 19174 8708 20334
rect 8772 20312 8800 21422
rect 8864 21418 8892 21626
rect 9048 21554 9076 22170
rect 9232 22166 9260 24006
rect 9220 22160 9272 22166
rect 9220 22102 9272 22108
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8852 21412 8904 21418
rect 8852 21354 8904 21360
rect 8864 21146 8892 21354
rect 9232 21146 9260 22102
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 8852 20324 8904 20330
rect 8772 20284 8852 20312
rect 8852 20266 8904 20272
rect 8864 20058 8892 20266
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 9232 18970 9260 20810
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8864 18290 8892 18566
rect 9048 18358 9076 18566
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7944 15638 7972 15982
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7944 13938 7972 15574
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 15162 8156 15438
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7760 13518 7972 13546
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 12986 7788 13398
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12646 7512 12718
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7380 11144 7432 11150
rect 7484 11121 7512 12582
rect 7576 12374 7604 12582
rect 7668 12374 7696 12650
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7852 11558 7880 12106
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11286 7880 11494
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7380 11086 7432 11092
rect 7470 11112 7526 11121
rect 7392 10266 7420 11086
rect 7470 11047 7526 11056
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7024 7886 7052 9930
rect 7472 9580 7524 9586
rect 7576 9568 7604 10474
rect 7852 10266 7880 11222
rect 7944 10577 7972 13518
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12714 8064 13194
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 11150 8064 12650
rect 8128 12102 8156 13126
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7930 10568 7986 10577
rect 8128 10538 8156 12038
rect 8220 10810 8248 16186
rect 8404 15910 8432 16594
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8496 16046 8524 16458
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 15570 8432 15846
rect 8482 15600 8538 15609
rect 8392 15564 8444 15570
rect 8482 15535 8484 15544
rect 8392 15506 8444 15512
rect 8536 15535 8538 15544
rect 8484 15506 8536 15512
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15026 8340 15302
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8404 13870 8432 15506
rect 8496 14822 8524 15506
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14657 8524 14758
rect 8482 14648 8538 14657
rect 8482 14583 8538 14592
rect 8484 14544 8536 14550
rect 8588 14532 8616 17138
rect 8956 17066 8984 17478
rect 9140 17202 9168 18090
rect 9324 17678 9352 24550
rect 9416 24274 9444 27520
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 9404 24268 9456 24274
rect 9404 24210 9456 24216
rect 9416 23866 9444 24210
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9416 23225 9444 23802
rect 9402 23216 9458 23225
rect 9402 23151 9458 23160
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9416 20058 9444 20878
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9784 19990 9812 22374
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 20602 9904 21014
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9784 19514 9812 19926
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9678 19408 9734 19417
rect 9678 19343 9734 19352
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9416 18426 9444 18702
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 18193 9536 18702
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9494 18184 9550 18193
rect 9494 18119 9550 18128
rect 9508 17746 9536 18119
rect 9600 17814 9628 18566
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8772 16182 8800 16390
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8772 15978 8800 16118
rect 8956 16114 8984 16390
rect 9034 16144 9090 16153
rect 8944 16108 8996 16114
rect 9140 16114 9168 17138
rect 9324 16794 9352 17614
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9034 16079 9090 16088
rect 9128 16108 9180 16114
rect 8944 16050 8996 16056
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8536 14504 8616 14532
rect 8484 14486 8536 14492
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8680 14074 8708 14418
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8864 13938 8892 15302
rect 9048 14482 9076 16079
rect 9128 16050 9180 16056
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15366 9352 15846
rect 9508 15638 9536 16662
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9140 14618 9168 14826
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9232 14346 9260 14826
rect 9324 14521 9352 15302
rect 9416 14550 9444 15302
rect 9404 14544 9456 14550
rect 9310 14512 9366 14521
rect 9404 14486 9456 14492
rect 9310 14447 9366 14456
rect 9508 14414 9536 15370
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8220 10606 8248 10746
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7930 10503 7986 10512
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8036 9722 8064 10066
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7524 9540 7604 9568
rect 7472 9522 7524 9528
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7116 9178 7144 9386
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7300 8974 7328 9386
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7576 8566 7604 9540
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7760 8498 7788 8774
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 8090 7788 8434
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7954 7880 9318
rect 8036 9042 8064 9658
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8634 8064 8978
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7208 6254 7236 6802
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6322 7420 6734
rect 7472 6384 7524 6390
rect 7524 6344 7604 6372
rect 7472 6326 7524 6332
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7392 5914 7420 6258
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6380 5370 6408 5782
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6472 4554 6500 5646
rect 6656 5302 6684 5646
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6564 3194 6592 4218
rect 7208 3738 7236 4558
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7392 3913 7420 4014
rect 7378 3904 7434 3913
rect 7378 3839 7434 3848
rect 7484 3738 7512 4966
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 7576 2650 7604 6344
rect 7668 4049 7696 7482
rect 7944 7274 7972 7686
rect 8220 7562 8248 10542
rect 8036 7534 8248 7562
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 4264 7788 6190
rect 7852 6118 7880 6870
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5370 7880 6054
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7852 4758 7880 5306
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 7840 4276 7892 4282
rect 7760 4236 7840 4264
rect 7654 4040 7710 4049
rect 7654 3975 7710 3984
rect 7668 3602 7696 3975
rect 7760 3602 7788 4236
rect 7840 4218 7892 4224
rect 7838 4176 7894 4185
rect 7838 4111 7894 4120
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7668 3058 7696 3538
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7852 2514 7880 4111
rect 7944 3194 7972 7210
rect 8036 6186 8064 7534
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 7002 8248 7142
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8220 6458 8248 6938
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8128 5710 8156 6326
rect 8312 6322 8340 13670
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12714 8432 13126
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8404 12442 8432 12650
rect 8496 12442 8524 13262
rect 8864 12442 8892 13874
rect 8956 12986 8984 14214
rect 9508 13814 9536 14350
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9416 13786 9536 13814
rect 9692 13814 9720 19343
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9784 18698 9812 18770
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9784 18086 9812 18634
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9772 18080 9824 18086
rect 9876 18057 9904 18090
rect 9772 18022 9824 18028
rect 9862 18048 9918 18057
rect 9784 17649 9812 18022
rect 9862 17983 9918 17992
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9770 17640 9826 17649
rect 9770 17575 9826 17584
rect 9876 16998 9904 17750
rect 9968 17202 9996 22986
rect 10060 19854 10088 25094
rect 10152 23866 10180 27526
rect 10414 27520 10470 27526
rect 11426 27554 11482 28000
rect 12438 27554 12494 28000
rect 11426 27526 11744 27554
rect 11426 27520 11482 27526
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 10612 24886 10640 25298
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10600 24880 10652 24886
rect 10230 24848 10286 24857
rect 10600 24822 10652 24828
rect 10230 24783 10286 24792
rect 10244 24750 10272 24783
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10428 23866 10456 24210
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10152 23662 10180 23802
rect 10140 23656 10192 23662
rect 10140 23598 10192 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10152 22642 10180 23258
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10244 22574 10272 23122
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22030 10732 22578
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10152 20942 10180 21966
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10704 21418 10732 21830
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10796 20534 10824 25094
rect 11164 24682 11192 25298
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11152 24676 11204 24682
rect 11152 24618 11204 24624
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10888 23662 10916 24006
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10980 23168 11008 23598
rect 11152 23588 11204 23594
rect 11152 23530 11204 23536
rect 11060 23180 11112 23186
rect 10980 23140 11060 23168
rect 11060 23122 11112 23128
rect 11072 22982 11100 23122
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10876 22500 10928 22506
rect 10876 22442 10928 22448
rect 10888 22234 10916 22442
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10876 21956 10928 21962
rect 10876 21898 10928 21904
rect 10888 21486 10916 21898
rect 11072 21894 11100 22918
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 11164 21128 11192 23530
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11256 21554 11284 21966
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11072 21100 11192 21128
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10796 20058 10824 20470
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10980 19990 11008 20402
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 19514 10088 19790
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10060 18290 10088 18906
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10140 18148 10192 18154
rect 10060 18108 10140 18136
rect 10060 18057 10088 18108
rect 10140 18090 10192 18096
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10046 18048 10102 18057
rect 10046 17983 10102 17992
rect 10060 17882 10088 17983
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9968 16794 9996 17138
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 16726 10088 17818
rect 10704 17202 10732 18090
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9876 16250 9904 16662
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 14550 9812 15846
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9876 15162 9904 15574
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9968 14890 9996 16050
rect 10232 15972 10284 15978
rect 10152 15932 10232 15960
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15026 10088 15438
rect 10152 15366 10180 15932
rect 10232 15914 10284 15920
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14550 10732 17138
rect 10796 16697 10824 17478
rect 10782 16688 10838 16697
rect 10782 16623 10838 16632
rect 10888 16590 10916 17614
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10888 15978 10916 16526
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 15434 10916 15914
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10796 14890 10824 15030
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10888 14618 10916 15370
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 9784 14074 9812 14486
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10980 13841 11008 19110
rect 11072 16658 11100 21100
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11256 20992 11284 21354
rect 11348 21146 11376 24754
rect 11716 24750 11744 27526
rect 12360 27526 12494 27554
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11716 24410 11744 24550
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11532 23186 11560 23530
rect 11704 23248 11756 23254
rect 11704 23190 11756 23196
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11716 22438 11744 23190
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 22166 11744 22374
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 11716 21350 11744 22102
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11336 21004 11388 21010
rect 11256 20964 11336 20992
rect 11164 20534 11192 20946
rect 11152 20528 11204 20534
rect 11150 20496 11152 20505
rect 11204 20496 11206 20505
rect 11150 20431 11206 20440
rect 11164 20405 11192 20431
rect 11256 19718 11284 20964
rect 11336 20946 11388 20952
rect 11808 20505 11836 24822
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23322 12112 23462
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11992 22778 12020 23054
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11794 20496 11850 20505
rect 11794 20431 11850 20440
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19310 11284 19654
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11886 19272 11942 19281
rect 11256 18630 11284 19246
rect 11886 19207 11942 19216
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11624 18426 11652 18702
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11532 17338 11560 17614
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 15065 11100 15302
rect 11058 15056 11114 15065
rect 11164 15026 11192 15506
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11058 14991 11114 15000
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 14618 11100 14758
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10966 13832 11022 13841
rect 9692 13786 10088 13814
rect 9232 13190 9260 13738
rect 9416 13530 9444 13786
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9048 12753 9076 12786
rect 9034 12744 9090 12753
rect 9034 12679 9090 12688
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11354 9076 11494
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8496 10130 8524 10610
rect 8956 10606 8984 11018
rect 9140 10674 9168 11630
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 9232 10198 9260 13126
rect 9692 12628 9720 13330
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9862 13288 9918 13297
rect 9784 12850 9812 13262
rect 9862 13223 9918 13232
rect 9876 12889 9904 13223
rect 9862 12880 9918 12889
rect 9772 12844 9824 12850
rect 9862 12815 9918 12824
rect 9772 12786 9824 12792
rect 9772 12640 9824 12646
rect 9692 12600 9772 12628
rect 9772 12582 9824 12588
rect 9496 11620 9548 11626
rect 9784 11608 9812 12582
rect 9876 12306 9904 12815
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 11898 9904 12242
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9864 11620 9916 11626
rect 9784 11580 9864 11608
rect 9496 11562 9548 11568
rect 9864 11562 9916 11568
rect 9310 11112 9366 11121
rect 9310 11047 9366 11056
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8496 9382 8524 10066
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8772 9586 8800 9998
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 7886 8524 9318
rect 8772 9178 8800 9522
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8588 8430 8616 8978
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 8090 8616 8366
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8588 6866 8616 8026
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8680 6390 8708 7210
rect 9048 7206 9076 7890
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8220 4826 8248 5782
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8036 4214 8064 4694
rect 8024 4208 8076 4214
rect 8312 4185 8340 6258
rect 8680 4826 8708 6326
rect 8864 6322 8892 6666
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8956 6186 8984 6394
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 9048 5545 9076 7142
rect 9232 6866 9260 8298
rect 9324 6905 9352 11047
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 7954 9444 8910
rect 9508 8537 9536 11562
rect 9876 11286 9904 11562
rect 9968 11286 9996 12038
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 10810 9996 11222
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9494 8528 9550 8537
rect 9494 8463 9550 8472
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9416 7546 9444 7890
rect 9600 7546 9628 10474
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9110 9720 9998
rect 9876 9722 9904 10406
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9722 9996 10134
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9968 9178 9996 9386
rect 9956 9172 10008 9178
rect 9876 9132 9956 9160
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9876 8634 9904 9132
rect 9956 9114 10008 9120
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9876 8022 9904 8570
rect 9968 8362 9996 8774
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9876 7002 9904 7958
rect 9968 7478 9996 8298
rect 10060 7546 10088 13786
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10784 13796 10836 13802
rect 11256 13814 11284 15302
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11256 13786 11376 13814
rect 10966 13767 11022 13776
rect 10784 13738 10836 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13394 10732 13738
rect 10796 13530 10824 13738
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12918 10732 13330
rect 11256 12918 11284 13398
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10600 12708 10652 12714
rect 10652 12668 10732 12696
rect 10600 12650 10652 12656
rect 10152 12374 10180 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10704 12170 10732 12668
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11694 10548 12038
rect 10704 11762 10732 12106
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10600 11280 10652 11286
rect 10796 11268 10824 12854
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10888 11898 10916 12310
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10652 11240 10824 11268
rect 10600 11222 10652 11228
rect 10612 10742 10640 11222
rect 10980 11082 11008 12582
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 9926 10732 10474
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10152 9178 10180 9658
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10152 8344 10180 9114
rect 10704 8566 10732 9862
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10888 9450 10916 9590
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10796 9330 10824 9386
rect 10980 9330 11008 9862
rect 11072 9654 11100 9930
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10796 9302 11008 9330
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10232 8356 10284 8362
rect 10152 8316 10232 8344
rect 10152 8090 10180 8316
rect 10232 8298 10284 8304
rect 10796 8242 10824 9302
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10796 8214 10916 8242
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10060 7342 10088 7482
rect 10428 7478 10456 7958
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10796 7002 10824 7210
rect 9864 6996 9916 7002
rect 9784 6956 9864 6984
rect 9310 6896 9366 6905
rect 9220 6860 9272 6866
rect 9310 6831 9366 6840
rect 9220 6802 9272 6808
rect 9034 5536 9090 5545
rect 9034 5471 9090 5480
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8680 4214 8708 4762
rect 8864 4758 8892 4966
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8668 4208 8720 4214
rect 8024 4150 8076 4156
rect 8298 4176 8354 4185
rect 8668 4150 8720 4156
rect 8298 4111 8354 4120
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8220 3738 8248 3946
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3670 8340 3946
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8850 3088 8906 3097
rect 8850 3023 8906 3032
rect 8864 2990 8892 3023
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5906 82 5962 480
rect 5552 54 5962 82
rect 7116 82 7144 2246
rect 7286 82 7342 480
rect 7116 54 7342 82
rect 8404 82 8432 2790
rect 9324 2514 9352 6831
rect 9784 6458 9812 6956
rect 9864 6938 9916 6944
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9784 6118 9812 6394
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5370 9812 6054
rect 9876 5914 9904 6802
rect 10796 6458 10824 6938
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10796 6186 10824 6394
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10060 5574 10088 6122
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10888 5914 10916 8214
rect 11072 8090 11100 8570
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11164 6662 11192 7346
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9508 4078 9536 4694
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3670 9536 4014
rect 9968 3942 9996 5102
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 10060 2650 10088 5510
rect 10704 5370 10732 5782
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4282 10732 4558
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 4218
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3058 10180 3334
rect 11164 3194 11192 6598
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11256 4282 11284 5578
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11256 3126 11284 3538
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 11348 2582 11376 13786
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11440 13705 11468 13738
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11440 12782 11468 13631
rect 11808 13433 11836 14486
rect 11794 13424 11850 13433
rect 11794 13359 11850 13368
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12986 11652 13262
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11440 12374 11468 12718
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11440 11898 11468 12106
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11440 11286 11468 11834
rect 11808 11762 11836 12310
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11440 10146 11468 11222
rect 11704 10192 11756 10198
rect 11440 10118 11560 10146
rect 11704 10134 11756 10140
rect 11532 10062 11560 10118
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11440 9178 11468 9998
rect 11716 9722 11744 10134
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11612 9376 11664 9382
rect 11664 9336 11744 9364
rect 11612 9318 11664 9324
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8294 11560 8978
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11532 7857 11560 8230
rect 11518 7848 11574 7857
rect 11518 7783 11574 7792
rect 11532 7546 11560 7783
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11440 6322 11468 7414
rect 11624 6934 11652 7686
rect 11716 7546 11744 9336
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11624 6458 11652 6870
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11440 5710 11468 6258
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11440 5370 11468 5646
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11440 4758 11468 5306
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11900 4154 11928 19207
rect 11992 14618 12020 21898
rect 12176 19938 12204 24618
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23730 12296 24006
rect 12360 23866 12388 27526
rect 12438 27520 12494 27526
rect 13450 27520 13506 28000
rect 14462 27520 14518 28000
rect 15382 27520 15438 28000
rect 16394 27520 16450 28000
rect 17406 27520 17462 28000
rect 18418 27554 18474 28000
rect 18248 27526 18474 27554
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24818 12848 25094
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12636 24342 12664 24550
rect 12624 24336 12676 24342
rect 12624 24278 12676 24284
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12268 22234 12296 23462
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 20262 12296 21286
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19990 12296 20198
rect 12084 19910 12204 19938
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12084 19281 12112 19910
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12176 19310 12204 19790
rect 12164 19304 12216 19310
rect 12070 19272 12126 19281
rect 12164 19246 12216 19252
rect 12070 19207 12126 19216
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12084 18902 12112 19110
rect 12176 18970 12204 19246
rect 12268 19174 12296 19926
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12084 18086 12112 18838
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 18154 12204 18566
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12176 16998 12204 17818
rect 12268 17814 12296 18226
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12084 16250 12112 16594
rect 12360 16561 12388 23802
rect 12636 23322 12664 24278
rect 12820 23474 12848 24754
rect 13464 24342 13492 27520
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 14016 24750 14044 25298
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13096 23798 13124 24074
rect 13084 23792 13136 23798
rect 13084 23734 13136 23740
rect 12728 23446 12848 23474
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12728 21690 12756 23446
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13004 22642 13032 23122
rect 13096 22982 13124 23734
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13176 23520 13228 23526
rect 13176 23462 13228 23468
rect 13188 23322 13216 23462
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13556 23254 13584 23530
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13556 22778 13584 23190
rect 13740 23118 13768 24550
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13740 22234 13768 23054
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13096 21894 13124 22102
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12452 20466 12480 20878
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 13096 20058 13124 21830
rect 13544 21616 13596 21622
rect 13544 21558 13596 21564
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13188 19718 13216 20878
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19378 13216 19654
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18902 12572 19110
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 13176 18896 13228 18902
rect 13176 18838 13228 18844
rect 12346 16552 12402 16561
rect 12346 16487 12402 16496
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12084 16017 12112 16186
rect 12070 16008 12126 16017
rect 12070 15943 12126 15952
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 15162 12296 15506
rect 12544 15366 12572 18838
rect 13188 18426 13216 18838
rect 13176 18420 13228 18426
rect 13096 18380 13176 18408
rect 13096 17882 13124 18380
rect 13176 18362 13228 18368
rect 13174 18320 13230 18329
rect 13174 18255 13230 18264
rect 13188 18222 13216 18255
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12636 17066 12664 17818
rect 13188 17270 13216 18158
rect 13280 17270 13308 20470
rect 13464 20262 13492 21014
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19990 13492 20198
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13464 17814 13492 18022
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13556 17542 13584 21558
rect 13832 21418 13860 22374
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13648 21146 13676 21354
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13648 20058 13676 21082
rect 13832 21010 13860 21354
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13924 20754 13952 24278
rect 14016 24274 14044 24686
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14016 23798 14044 24210
rect 14004 23792 14056 23798
rect 14004 23734 14056 23740
rect 14108 23730 14136 25094
rect 14476 24857 14504 27520
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14462 24848 14518 24857
rect 14462 24783 14518 24792
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14476 23730 14504 24618
rect 14096 23724 14148 23730
rect 14096 23666 14148 23672
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14108 23322 14136 23666
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14016 21554 14044 22918
rect 14292 21894 14320 23530
rect 14476 23118 14504 23666
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14568 23050 14596 24686
rect 14752 24614 14780 25298
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14280 21888 14332 21894
rect 14280 21830 14332 21836
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13832 20726 13952 20754
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13832 18737 13860 20726
rect 14016 20534 14044 21490
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14476 20466 14504 21898
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14384 20058 14412 20402
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14292 19174 14320 19858
rect 14476 19446 14504 20402
rect 14464 19440 14516 19446
rect 14568 19417 14596 22986
rect 14464 19382 14516 19388
rect 14554 19408 14610 19417
rect 14554 19343 14610 19352
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13924 18766 13952 19110
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 13912 18760 13964 18766
rect 13818 18728 13874 18737
rect 13912 18702 13964 18708
rect 13818 18663 13874 18672
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13280 17116 13308 17206
rect 13096 17088 13308 17116
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16250 12664 16594
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12636 15026 12664 16186
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 14482 12020 14554
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11992 14074 12020 14418
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12162 13832 12218 13841
rect 12162 13767 12218 13776
rect 12176 12986 12204 13767
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12176 12782 12204 12922
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11354 12388 12174
rect 12452 11898 12480 14350
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 10538 12020 11154
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 7954 12020 8842
rect 12162 8528 12218 8537
rect 12162 8463 12218 8472
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11992 7206 12020 7890
rect 12084 7410 12112 7890
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6118 12020 6734
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12084 6390 12112 6666
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11716 4126 11928 4154
rect 11520 4072 11572 4078
rect 11440 4049 11520 4060
rect 11426 4040 11520 4049
rect 11482 4032 11520 4040
rect 11520 4014 11572 4020
rect 11426 3975 11482 3984
rect 11716 3505 11744 4126
rect 11702 3496 11758 3505
rect 11702 3431 11758 3440
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 8574 82 8630 480
rect 8404 54 8630 82
rect 4618 0 4674 54
rect 5906 0 5962 54
rect 7286 0 7342 54
rect 8574 0 8630 54
rect 9954 82 10010 480
rect 10060 82 10088 2314
rect 9954 54 10088 82
rect 11242 82 11298 480
rect 11440 82 11468 3334
rect 11716 2990 11744 3431
rect 11992 3194 12020 6054
rect 12176 5778 12204 8463
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 5370 12204 5714
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12452 5166 12480 7142
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4758 12480 5102
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4282 12204 4626
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12544 2990 12572 14826
rect 12636 14482 12664 14962
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12728 13938 12756 16526
rect 12820 16182 12848 16934
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12820 15706 12848 16118
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 14822 12848 15642
rect 13096 15162 13124 17088
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13096 14958 13124 15098
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14006 12848 14758
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12820 13802 12848 13942
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 13530 12848 13738
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 11898 12848 13466
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 12646 12940 12718
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 11626 12848 11834
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12636 9382 12664 10066
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 8498 12664 9318
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12636 7954 12664 8434
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 6934 12664 7210
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12636 5574 12664 5850
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5166 12664 5510
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12636 2922 12664 3878
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 11242 54 11468 82
rect 12622 82 12678 480
rect 12728 82 12756 10542
rect 13004 10266 13032 10950
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 8838 12848 9386
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 7528 12848 8774
rect 12912 8090 12940 8910
rect 13004 8566 13032 9046
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13004 8362 13032 8502
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13004 7886 13032 8298
rect 13096 8294 13124 10474
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12820 7500 12940 7528
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 6662 12848 7346
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 4826 12848 6598
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12912 2650 12940 7500
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5574 13032 6190
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5234 13032 5510
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13188 4978 13216 16186
rect 13280 13326 13308 16458
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15978 13400 16390
rect 13464 16114 13492 16662
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15978 13492 16050
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13372 14385 13400 15914
rect 13464 15706 13492 15914
rect 13740 15706 13768 16526
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13740 15473 13768 15642
rect 13832 15609 13860 18663
rect 13924 18426 13952 18702
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13924 17814 13952 18090
rect 14108 17814 14136 18838
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 14096 17808 14148 17814
rect 14096 17750 14148 17756
rect 13924 17338 13952 17750
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14016 16998 14044 17138
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 15706 14044 16934
rect 14094 16688 14150 16697
rect 14094 16623 14150 16632
rect 14108 16250 14136 16623
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13818 15600 13874 15609
rect 13818 15535 13874 15544
rect 13726 15464 13782 15473
rect 13726 15399 13782 15408
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 14482 13492 14758
rect 13912 14544 13964 14550
rect 13740 14504 13912 14532
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13358 14376 13414 14385
rect 13358 14311 13414 14320
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13462 13400 13670
rect 13464 13530 13492 14418
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 13870 13584 14350
rect 13740 14006 13768 14504
rect 13912 14486 13964 14492
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13544 13864 13596 13870
rect 14292 13814 14320 19110
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14384 15162 14412 15506
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14384 14890 14412 15098
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 13544 13806 13596 13812
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 12238 13400 13398
rect 13452 12640 13504 12646
rect 13556 12628 13584 13806
rect 14200 13786 14320 13814
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13504 12600 13584 12628
rect 13452 12582 13504 12588
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13372 11354 13400 11562
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13372 10742 13400 11290
rect 13360 10736 13412 10742
rect 13280 10696 13360 10724
rect 13280 9110 13308 10696
rect 13360 10678 13412 10684
rect 13360 10124 13412 10130
rect 13464 10112 13492 12582
rect 13648 12442 13676 13262
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 10538 13768 11766
rect 14200 11121 14228 13786
rect 14384 13462 14412 14214
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 11762 14320 13262
rect 14476 12714 14504 18022
rect 14660 16697 14688 23734
rect 14844 23254 14872 25094
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15396 24410 15424 27520
rect 16408 24954 16436 27520
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 15844 24676 15896 24682
rect 15844 24618 15896 24624
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 14832 23248 14884 23254
rect 14832 23190 14884 23196
rect 14844 22234 14872 23190
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22642 15332 22918
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15212 21049 15240 21422
rect 15304 21146 15332 22578
rect 15396 22098 15424 23734
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15488 22506 15516 23054
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15396 21622 15424 22034
rect 15488 22030 15516 22442
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15198 21040 15254 21049
rect 15198 20975 15254 20984
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15396 20602 15424 20946
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18873 14872 19246
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 14830 18864 14886 18873
rect 14830 18799 14886 18808
rect 15120 18766 15148 19178
rect 15488 18970 15516 19858
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 14844 18426 14872 18702
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14844 18154 14872 18362
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 15120 17610 15148 18158
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14738 17232 14794 17241
rect 14738 17167 14794 17176
rect 14752 17134 14780 17167
rect 14844 17134 14872 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14844 16794 14872 16934
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14936 16726 14964 17002
rect 14924 16720 14976 16726
rect 14646 16688 14702 16697
rect 14924 16662 14976 16668
rect 14646 16623 14702 16632
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14924 16040 14976 16046
rect 14646 16008 14702 16017
rect 14924 15982 14976 15988
rect 14646 15943 14702 15952
rect 14740 15972 14792 15978
rect 14660 13818 14688 15943
rect 14740 15914 14792 15920
rect 14752 15026 14780 15914
rect 14936 15706 14964 15982
rect 15304 15978 15332 16186
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15396 14414 15424 16050
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15200 13864 15252 13870
rect 14738 13832 14794 13841
rect 14660 13790 14738 13818
rect 15396 13814 15424 14350
rect 15200 13806 15252 13812
rect 14738 13767 14794 13776
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11801 14412 12242
rect 14370 11792 14426 11801
rect 14280 11756 14332 11762
rect 14370 11727 14426 11736
rect 14280 11698 14332 11704
rect 14186 11112 14242 11121
rect 14186 11047 14242 11056
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10674 14136 10950
rect 14292 10674 14320 11698
rect 14384 11626 14412 11727
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14384 10577 14412 11562
rect 14370 10568 14426 10577
rect 13728 10532 13780 10538
rect 14370 10503 14426 10512
rect 13728 10474 13780 10480
rect 13740 10266 13768 10474
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13412 10084 13492 10112
rect 13360 10066 13412 10072
rect 13372 9722 13400 10066
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13556 6934 13584 9590
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 13740 9178 13768 9318
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 14108 7954 14136 8871
rect 14200 8362 14228 9318
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14476 8242 14504 12650
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 10742 14596 11290
rect 14660 10810 14688 11766
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 9110 14596 9318
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14568 8634 14596 9046
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8566 14688 10202
rect 14752 10130 14780 13767
rect 15212 13734 15240 13806
rect 15304 13786 15424 13814
rect 15488 13802 15516 14486
rect 15580 13814 15608 24210
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15672 20058 15700 23462
rect 15752 23248 15804 23254
rect 15856 23225 15884 24618
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 23322 15976 24550
rect 17420 24410 17448 27520
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 16592 23866 16620 24210
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 15752 23190 15804 23196
rect 15842 23216 15898 23225
rect 15764 22778 15792 23190
rect 15842 23151 15898 23160
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15750 22536 15806 22545
rect 15750 22471 15806 22480
rect 15764 21010 15792 22471
rect 15856 22234 15884 23151
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 15844 22228 15896 22234
rect 15844 22170 15896 22176
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15856 21554 15884 21966
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15856 21146 15884 21490
rect 15948 21486 15976 22102
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16132 20534 16160 20742
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15672 19378 15700 19994
rect 16224 19922 16252 22374
rect 16684 22098 16712 22510
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 21078 16528 21490
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16684 21078 16712 21286
rect 16488 21072 16540 21078
rect 16488 21014 16540 21020
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16776 20942 16804 22918
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16592 20466 16620 20810
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 20058 16436 20198
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15856 18902 15884 19382
rect 16316 19174 16344 19926
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15856 18426 15884 18838
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 16028 18352 16080 18358
rect 16028 18294 16080 18300
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15638 15792 15846
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 15094 15700 15438
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15764 14890 15792 15574
rect 15660 14884 15712 14890
rect 15660 14826 15712 14832
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15672 14770 15700 14826
rect 15856 14770 15884 18090
rect 16040 17814 16068 18294
rect 16028 17808 16080 17814
rect 15934 17776 15990 17785
rect 16028 17750 16080 17756
rect 15934 17711 15990 17720
rect 15948 17678 15976 17711
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 17542 15976 17614
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16040 17338 16068 17750
rect 16224 17610 16252 18702
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16224 17066 16252 17546
rect 16592 17202 16620 20402
rect 16776 20058 16804 20878
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16868 18698 16896 22442
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17052 20874 17080 21422
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 17144 20602 17172 21014
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17236 19378 17264 23258
rect 17512 23186 17540 23530
rect 17696 23526 17724 24210
rect 18248 23866 18276 27526
rect 18418 27520 18474 27526
rect 19430 27520 19486 28000
rect 20442 27554 20498 28000
rect 20364 27526 20498 27554
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17420 22420 17448 23122
rect 17512 22778 17540 23122
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17500 22432 17552 22438
rect 17420 22392 17500 22420
rect 17500 22374 17552 22380
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17328 19514 17356 19790
rect 17420 19514 17448 19926
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17408 18896 17460 18902
rect 17222 18864 17278 18873
rect 17408 18838 17460 18844
rect 17222 18799 17278 18808
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16868 18426 16896 18634
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16486 17096 16542 17105
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16304 17060 16356 17066
rect 16486 17031 16542 17040
rect 16304 17002 16356 17008
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16132 16250 16160 16662
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16224 15434 16252 17002
rect 16316 16794 16344 17002
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16500 16182 16528 17031
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 15672 14742 15884 14770
rect 15476 13796 15528 13802
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15304 13530 15332 13786
rect 15580 13786 15792 13814
rect 15476 13738 15528 13744
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13398
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15672 12442 15700 12718
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14844 10169 14872 11562
rect 14936 11354 14964 11562
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15396 11286 15424 12038
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15488 11286 15516 11834
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15476 11280 15528 11286
rect 15528 11240 15608 11268
rect 15476 11222 15528 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11222
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15488 10538 15516 10678
rect 15580 10674 15608 11240
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 14830 10160 14886 10169
rect 14740 10124 14792 10130
rect 14830 10095 14886 10104
rect 14740 10066 14792 10072
rect 15396 9926 15424 10474
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14200 8214 14504 8242
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 13648 7478 13676 7890
rect 14108 7546 14136 7890
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 13372 5846 13400 6122
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13372 5370 13400 5782
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13096 4950 13216 4978
rect 13096 4690 13124 4950
rect 13464 4826 13492 5646
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13188 3738 13216 4762
rect 13556 4690 13584 5102
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13280 4154 13308 4422
rect 13464 4282 13492 4422
rect 13556 4282 13584 4626
rect 13740 4554 13768 6734
rect 13832 6458 13860 6870
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14108 5914 14136 7482
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14004 5160 14056 5166
rect 14200 5137 14228 8214
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7342 14504 7686
rect 14752 7546 14780 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15672 9722 15700 10066
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14844 8838 14872 9386
rect 14936 9110 14964 9386
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 15212 8906 15240 9590
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14384 5370 14412 5510
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14004 5102 14056 5108
rect 14186 5128 14242 5137
rect 14016 4826 14044 5102
rect 14186 5063 14242 5072
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13280 4126 13400 4154
rect 13372 3738 13400 4126
rect 13452 4072 13504 4078
rect 13556 4060 13584 4218
rect 13504 4032 13584 4060
rect 13452 4014 13504 4020
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13372 3602 13400 3674
rect 13464 3670 13492 4014
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13372 3194 13400 3538
rect 13924 3194 13952 3538
rect 14292 3194 14320 5238
rect 14476 4078 14504 7278
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 5574 14780 6190
rect 14740 5568 14792 5574
rect 14554 5536 14610 5545
rect 14740 5510 14792 5516
rect 14554 5471 14610 5480
rect 14568 4214 14596 5471
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14752 4146 14780 5510
rect 14844 4282 14872 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8090 15332 8842
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15396 8090 15424 8298
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7546 15424 8026
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15488 7478 15516 9386
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15580 7274 15608 7482
rect 15672 7426 15700 8230
rect 15764 7546 15792 13786
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 16040 12986 16068 13738
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15948 11082 15976 12786
rect 16040 12646 16068 12922
rect 16592 12753 16620 17138
rect 17236 16658 17264 18799
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17328 17610 17356 18702
rect 17420 18426 17448 18838
rect 17512 18630 17540 22374
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17604 19854 17632 20470
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17604 18766 17632 19790
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17406 18184 17462 18193
rect 17406 18119 17462 18128
rect 17420 17746 17448 18119
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17420 17338 17448 17682
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 16250 17264 16594
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17144 15162 17172 15302
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 13326 16804 14350
rect 16960 14074 16988 14554
rect 17144 14482 17172 15098
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17144 14006 17172 14418
rect 17132 14000 17184 14006
rect 17184 13960 17264 13988
rect 17132 13942 17184 13948
rect 17236 13814 17264 13960
rect 17328 13938 17356 14418
rect 17420 14074 17448 17274
rect 17512 16697 17540 18022
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17604 15026 17632 18702
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17236 13786 17356 13814
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16960 12986 16988 13398
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17052 12850 17080 13262
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16578 12744 16634 12753
rect 16396 12708 16448 12714
rect 16578 12679 16634 12688
rect 16396 12650 16448 12656
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 11762 16068 12038
rect 16408 11762 16436 12650
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12374 16620 12582
rect 17144 12374 17172 13194
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 16592 11898 16620 12310
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16684 11762 16712 12174
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16408 11354 16436 11698
rect 16684 11354 16712 11698
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15948 10742 15976 11018
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 16776 10266 16804 11086
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9722 15884 10066
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15856 8945 15884 9658
rect 16500 9450 16528 9862
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 15842 8936 15898 8945
rect 15842 8871 15898 8880
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15948 8362 15976 8842
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15672 7398 15792 7426
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15396 6662 15424 7210
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15580 6118 15608 6870
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 4826 15424 5646
rect 15488 5370 15516 5782
rect 15580 5370 15608 6054
rect 15672 5710 15700 6666
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15580 4758 15608 5306
rect 15672 5302 15700 5646
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 15396 4264 15424 4558
rect 15476 4276 15528 4282
rect 15396 4236 15476 4264
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12622 54 12756 82
rect 13740 82 13768 2994
rect 14292 2990 14320 3130
rect 14476 3097 14504 4014
rect 15396 3738 15424 4236
rect 15476 4218 15528 4224
rect 15580 4214 15608 4694
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14462 3088 14518 3097
rect 14462 3023 14518 3032
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 13910 82 13966 480
rect 13740 54 13966 82
rect 9954 0 10010 54
rect 11242 0 11298 54
rect 12622 0 12678 54
rect 13910 0 13966 54
rect 15290 82 15346 480
rect 15764 82 15792 7398
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15856 4282 15884 6598
rect 15948 5642 15976 8298
rect 16500 8090 16528 9386
rect 16592 8838 16620 9386
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 16040 6934 16068 7414
rect 16316 7206 16344 7890
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7206 16804 7822
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16040 5234 16068 6870
rect 16316 6225 16344 7142
rect 16776 7002 16804 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16302 6216 16358 6225
rect 16302 6151 16358 6160
rect 16408 6118 16436 6734
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16040 4826 16068 5170
rect 16408 4826 16436 6054
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16868 4690 16896 10542
rect 16946 9072 17002 9081
rect 16946 9007 17002 9016
rect 16960 8974 16988 9007
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8090 16988 8910
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17144 6866 17172 11018
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17236 10266 17264 10610
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 10130 17356 13786
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 8974 17264 9522
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17328 8362 17356 9318
rect 17512 9024 17540 14486
rect 17696 14346 17724 23462
rect 18984 23186 19012 26862
rect 19444 24410 19472 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17788 22098 17816 23054
rect 18984 22778 19012 23122
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18694 22672 18750 22681
rect 18694 22607 18750 22616
rect 18328 22432 18380 22438
rect 18248 22392 18328 22420
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17788 21690 17816 22034
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17972 21418 18000 22102
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17880 20602 17908 20878
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17880 19514 17908 20538
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17270 17908 17682
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17880 16794 17908 17206
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17880 16114 17908 16730
rect 17972 16182 18000 17206
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17880 15570 17908 16050
rect 18064 16017 18092 18158
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18050 16008 18106 16017
rect 18050 15943 18106 15952
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15162 17908 15506
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17880 13870 17908 14010
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17590 11656 17646 11665
rect 17590 11591 17646 11600
rect 17604 11150 17632 11591
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 10130 17632 11086
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17604 9194 17632 10066
rect 17696 9489 17724 13126
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11558 17816 12242
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11257 17816 11494
rect 17774 11248 17830 11257
rect 17880 11218 17908 13806
rect 17774 11183 17830 11192
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17682 9480 17738 9489
rect 17682 9415 17738 9424
rect 17788 9382 17816 10406
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17604 9166 17724 9194
rect 17592 9036 17644 9042
rect 17512 8996 17592 9024
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17328 8022 17356 8298
rect 17316 8016 17368 8022
rect 17316 7958 17368 7964
rect 17328 7546 17356 7958
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17144 6458 17172 6802
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17236 6390 17264 6802
rect 17328 6390 17356 7482
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17316 6384 17368 6390
rect 17316 6326 17368 6332
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5234 16988 5646
rect 17052 5370 17080 5782
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 4049 16160 4082
rect 16118 4040 16174 4049
rect 16118 3975 16174 3984
rect 16868 3942 16896 4626
rect 17512 4154 17540 8996
rect 17592 8978 17644 8984
rect 17696 8974 17724 9166
rect 17684 8968 17736 8974
rect 17736 8928 17816 8956
rect 17684 8910 17736 8916
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17696 8090 17724 8774
rect 17788 8634 17816 8928
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17788 8022 17816 8570
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17788 6866 17816 7958
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17328 4126 17540 4154
rect 17972 4154 18000 15370
rect 18064 12918 18092 15943
rect 18156 15502 18184 17614
rect 18248 16153 18276 22392
rect 18328 22374 18380 22380
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18432 20466 18460 21286
rect 18616 21078 18644 21830
rect 18708 21554 18736 22607
rect 19076 21622 19104 23462
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18616 20602 18644 21014
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 17338 18368 18566
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18234 16144 18290 16153
rect 18234 16079 18290 16088
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18340 13734 18368 16526
rect 18432 16046 18460 19654
rect 18524 18970 18552 20470
rect 18616 20312 18644 20538
rect 18696 20324 18748 20330
rect 18616 20284 18696 20312
rect 18616 20058 18644 20284
rect 18696 20266 18748 20272
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18800 19446 18828 20878
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18616 19281 18644 19314
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18800 18329 18828 19382
rect 18984 18970 19012 19722
rect 19076 19281 19104 21558
rect 19260 21554 19288 21830
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20040 19380 21286
rect 19444 20942 19472 22578
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19432 20052 19484 20058
rect 19352 20012 19432 20040
rect 19432 19994 19484 20000
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19260 19378 19288 19858
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19062 19272 19118 19281
rect 19062 19207 19118 19216
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18786 18320 18842 18329
rect 18786 18255 18842 18264
rect 18892 17814 18920 18634
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18984 17746 19012 18294
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18984 17338 19012 17682
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18602 16144 18658 16153
rect 18602 16079 18658 16088
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15162 18460 15982
rect 18512 15360 18564 15366
rect 18616 15337 18644 16079
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18512 15302 18564 15308
rect 18602 15328 18658 15337
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 14958 18460 15098
rect 18524 14958 18552 15302
rect 18602 15263 18658 15272
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18708 14890 18736 15438
rect 19076 15434 19104 19207
rect 19444 19174 19472 19994
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19260 18902 19288 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19260 18086 19288 18838
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 18086 19380 18158
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19260 16998 19288 18022
rect 19444 17882 19472 18090
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 19260 15910 19288 16934
rect 19536 16590 19564 23734
rect 20364 23497 20392 27526
rect 20442 27520 20498 27526
rect 21454 27520 21510 28000
rect 22374 27520 22430 28000
rect 23386 27520 23442 28000
rect 24398 27554 24454 28000
rect 25410 27554 25466 28000
rect 24136 27526 24454 27554
rect 20350 23488 20406 23497
rect 19622 23420 19918 23440
rect 20350 23423 20406 23432
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20364 23050 20392 23423
rect 21468 23322 21496 27520
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19904 22642 19932 22918
rect 19892 22636 19944 22642
rect 20260 22636 20312 22642
rect 19944 22596 20024 22624
rect 19892 22578 19944 22584
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19996 22234 20024 22596
rect 20260 22578 20312 22584
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 20088 21690 20116 22442
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 20088 18290 20116 21082
rect 20272 20466 20300 22578
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22166 21036 22374
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20364 21622 20392 22034
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20272 19922 20300 20402
rect 20364 20330 20392 20742
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20364 20058 20392 20266
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 21088 19984 21140 19990
rect 21088 19926 21140 19932
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20640 18970 20668 19450
rect 21008 19174 21036 19790
rect 21100 19514 21128 19926
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21192 19378 21220 21966
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 21010 21312 21286
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21284 20466 21312 20946
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21284 19854 21312 20266
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21284 19378 21312 19790
rect 21376 19718 21404 21422
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21272 19372 21324 19378
rect 21324 19332 21404 19360
rect 21272 19314 21324 19320
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18970 21036 19110
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18902 21220 19314
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20088 17814 20116 18226
rect 20640 17882 20668 18702
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20088 16833 20116 17614
rect 20916 17241 20944 18226
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 21008 17762 21036 18022
rect 21100 17882 21128 18838
rect 21284 18426 21312 19178
rect 21376 18766 21404 19332
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21284 17762 21312 18090
rect 21008 17734 21312 17762
rect 20902 17232 20958 17241
rect 20902 17167 20958 17176
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20074 16824 20130 16833
rect 20074 16759 20130 16768
rect 20088 16726 20116 16759
rect 20456 16726 20484 16934
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15638 19564 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19064 15428 19116 15434
rect 19064 15370 19116 15376
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18708 14618 18736 14826
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18892 14482 18920 14894
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18432 14074 18460 14418
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18892 13870 18920 14418
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18880 13864 18932 13870
rect 19352 13841 19380 15098
rect 19536 14822 19564 15574
rect 19892 15360 19944 15366
rect 19996 15348 20024 16050
rect 19944 15320 20024 15348
rect 19892 15302 19944 15308
rect 19904 15026 19932 15302
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 18880 13806 18932 13812
rect 19338 13832 19394 13841
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18524 13190 18552 13806
rect 19338 13767 19394 13776
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19168 13462 19196 13670
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18524 12345 18552 12718
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 11626 18276 12174
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18248 11354 18276 11562
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18432 10810 18460 11154
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18432 10198 18460 10746
rect 18524 10674 18552 11290
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 9586 18092 9998
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 9178 18092 9522
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18248 8906 18276 9386
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18432 8634 18460 8978
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 7410 18092 8434
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18432 7206 18460 7890
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18326 6352 18382 6361
rect 18326 6287 18382 6296
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18064 5914 18092 6190
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18340 5778 18368 6287
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18340 5370 18368 5714
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 17972 4126 18184 4154
rect 17328 4010 17356 4126
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3602 16896 3878
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 18156 2854 18184 4126
rect 18432 3670 18460 7142
rect 18616 6866 18644 12786
rect 19168 12646 19196 13398
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18984 10062 19012 12038
rect 19076 11014 19104 12038
rect 19168 11558 19196 12378
rect 19352 11898 19380 13767
rect 19444 13705 19472 13942
rect 19536 13802 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19720 13938 19748 14214
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19430 13696 19486 13705
rect 19430 13631 19486 13640
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20272 12374 20300 12582
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 10198 19104 10542
rect 19168 10470 19196 11494
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18984 9178 19012 9998
rect 19076 9722 19104 10134
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18892 7936 18920 8978
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18984 8498 19012 8910
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 18972 7948 19024 7954
rect 18892 7908 18972 7936
rect 18972 7890 19024 7896
rect 18984 7546 19012 7890
rect 19168 7546 19196 8298
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 18984 6866 19012 7482
rect 19168 7274 19196 7482
rect 19260 7410 19288 7822
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19260 7002 19288 7346
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 18616 6254 18644 6802
rect 18984 6440 19012 6802
rect 19064 6452 19116 6458
rect 18984 6412 19064 6440
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 4486 18644 6190
rect 18984 5778 19012 6412
rect 19064 6394 19116 6400
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18984 4826 19012 5714
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19168 5166 19196 5306
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 19168 5030 19196 5102
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 19168 4146 19196 4966
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18156 2417 18184 2790
rect 18142 2408 18198 2417
rect 16856 2372 16908 2378
rect 18142 2343 18198 2352
rect 16856 2314 16908 2320
rect 15290 54 15792 82
rect 16578 82 16634 480
rect 16868 82 16896 2314
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 16578 54 16896 82
rect 17788 82 17816 2246
rect 17958 82 18014 480
rect 17788 54 18014 82
rect 19076 82 19104 4014
rect 19352 3194 19380 11562
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 10674 20024 11494
rect 20088 11150 20116 11630
rect 20456 11150 20484 16526
rect 20548 16250 20576 16934
rect 20732 16454 20760 17002
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 16250 20760 16390
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20824 16182 20852 16662
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20916 15450 20944 17167
rect 21008 17066 21036 17734
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20996 16788 21048 16794
rect 21048 16748 21128 16776
rect 20996 16730 21048 16736
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 15638 21036 16390
rect 21100 16182 21128 16748
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 21100 15638 21128 16118
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15706 21312 15846
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 20720 15428 20772 15434
rect 20916 15422 21036 15450
rect 20720 15370 20772 15376
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14074 20576 14962
rect 20732 14414 20760 15370
rect 20904 15360 20956 15366
rect 20904 15302 20956 15308
rect 20916 14890 20944 15302
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20916 14618 20944 14826
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20548 13190 20576 13670
rect 20732 13530 20760 14350
rect 21008 13814 21036 15422
rect 21100 15162 21128 15574
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 21100 14890 21128 14962
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21100 14074 21128 14486
rect 21192 14385 21220 14758
rect 21178 14376 21234 14385
rect 21178 14311 21234 14320
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20916 13786 21036 13814
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 11898 20576 13126
rect 20824 12782 20852 13466
rect 20916 13394 20944 13786
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 12986 20944 13330
rect 21100 13258 21128 14010
rect 21468 13870 21496 20878
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 19786 21864 20198
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21652 16590 21680 17002
rect 21836 16998 21864 17750
rect 21928 17678 21956 24006
rect 22388 23866 22416 27520
rect 23400 26926 23428 27520
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 23124 23730 23152 24210
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 22020 22234 22048 22510
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22296 21690 22324 22102
rect 22664 21690 22692 22374
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22020 19990 22048 20334
rect 22480 20330 22508 20946
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22468 20324 22520 20330
rect 22468 20266 22520 20272
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 22020 18290 22048 19926
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 18834 22416 19178
rect 22480 19174 22508 19858
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22282 18728 22338 18737
rect 22282 18663 22338 18672
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21836 16726 21864 16934
rect 21928 16794 21956 17614
rect 22112 17610 22140 18090
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21822 16552 21878 16561
rect 21822 16487 21878 16496
rect 21836 15586 21864 16487
rect 21916 16108 21968 16114
rect 22020 16096 22048 17478
rect 22204 17338 22232 18022
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22296 17270 22324 18663
rect 22388 18358 22416 18770
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22296 17134 22324 17206
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 21968 16068 22048 16096
rect 21916 16050 21968 16056
rect 22020 15706 22048 16068
rect 22112 15978 22140 16526
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 21836 15558 21956 15586
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15162 21864 15438
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 15088 21784 15094
rect 21928 15042 21956 15558
rect 22112 15434 22140 15914
rect 22388 15910 22416 18022
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22204 15706 22232 15846
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 21732 15030 21784 15036
rect 21640 14884 21692 14890
rect 21640 14826 21692 14832
rect 21652 14550 21680 14826
rect 21744 14550 21772 15030
rect 21836 15014 21956 15042
rect 22376 15088 22428 15094
rect 22376 15030 22428 15036
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21180 13864 21232 13870
rect 21456 13864 21508 13870
rect 21232 13824 21456 13852
rect 21180 13806 21232 13812
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21192 13394 21220 13670
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 13138 21220 13194
rect 21100 13110 21220 13138
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20732 12442 20760 12582
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20640 11354 20668 12310
rect 20824 12306 20852 12718
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 21100 11694 21128 13110
rect 21284 12714 21312 13126
rect 21376 12850 21404 13824
rect 21652 13814 21680 14486
rect 21456 13806 21508 13812
rect 21560 13786 21680 13814
rect 21560 12850 21588 13786
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21192 12442 21220 12650
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21560 12170 21588 12786
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20824 11558 20852 11630
rect 21284 11558 21312 12106
rect 21560 11626 21588 12106
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10266 20024 10610
rect 20456 10266 20484 11086
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19628 9654 19656 9998
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20272 9178 20300 9522
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19904 8634 19932 9046
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8634 20300 8910
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20640 6866 20668 7142
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6390 20024 6598
rect 19984 6384 20036 6390
rect 20824 6361 20852 11494
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10062 21036 10950
rect 21100 10810 21128 11222
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21100 10198 21128 10746
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21008 9178 21036 9998
rect 21100 9722 21128 10134
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21284 9654 21312 9998
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 21284 8906 21312 9590
rect 21468 9450 21496 9590
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21192 8362 21220 8842
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 20916 7478 20944 8298
rect 21192 8022 21220 8298
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21100 7546 21128 7958
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20996 6928 21048 6934
rect 20996 6870 21048 6876
rect 21008 6458 21036 6870
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 19984 6326 20036 6332
rect 20810 6352 20866 6361
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19536 5914 19564 6258
rect 19996 6186 20024 6326
rect 21192 6322 21220 7958
rect 21284 7886 21312 8842
rect 21468 8566 21496 9386
rect 21560 9178 21588 9386
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 8634 21772 9046
rect 21836 9042 21864 15014
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21928 13394 21956 13806
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22204 12646 22232 13330
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22020 10674 22048 11086
rect 22204 11082 22232 12582
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21928 10266 21956 10610
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22020 9432 22048 10610
rect 22296 10470 22324 11154
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9586 22140 9862
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22100 9444 22152 9450
rect 22020 9404 22100 9432
rect 22100 9386 22152 9392
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21652 8294 21680 8434
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21284 7002 21312 7822
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21376 6458 21404 6734
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 20810 6287 20866 6296
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 21192 5778 21220 6258
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3738 20024 3975
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19720 3194 19748 3538
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19352 2990 19380 3130
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19168 2514 19196 2790
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 19246 82 19302 480
rect 19076 54 19302 82
rect 15290 0 15346 54
rect 16578 0 16634 54
rect 17958 0 18014 54
rect 19246 0 19302 54
rect 20626 82 20682 480
rect 20732 82 20760 4082
rect 21468 2514 21496 8026
rect 21652 6866 21680 8230
rect 21744 6934 21772 8570
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22020 7857 22048 8366
rect 22112 8294 22140 9386
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22006 7848 22062 7857
rect 22006 7783 22062 7792
rect 22020 7750 22048 7783
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 22204 6798 22232 8230
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22296 4154 22324 10406
rect 22388 5370 22416 15030
rect 22480 13258 22508 19110
rect 22756 18816 22784 20810
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22848 19922 22876 20402
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22848 19242 22876 19858
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 22836 18828 22888 18834
rect 22756 18788 22836 18816
rect 22836 18770 22888 18776
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22572 16726 22600 18566
rect 22848 18086 22876 18770
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22572 16182 22600 16662
rect 22560 16176 22612 16182
rect 22560 16118 22612 16124
rect 22664 16114 22692 16662
rect 22756 16590 22784 17546
rect 22848 16998 22876 17682
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22744 16584 22796 16590
rect 22848 16561 22876 16934
rect 22744 16526 22796 16532
rect 22834 16552 22890 16561
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22572 15638 22600 15914
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22572 15026 22600 15574
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22664 13394 22692 15846
rect 22756 15502 22784 16526
rect 22834 16487 22890 16496
rect 22940 16114 22968 23462
rect 23570 19272 23626 19281
rect 23570 19207 23626 19216
rect 23584 18222 23612 19207
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23676 18970 23704 19110
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 17678 23244 18022
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23216 16454 23244 16934
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22756 13802 22784 14418
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22756 13462 22784 13738
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22468 12912 22520 12918
rect 22468 12854 22520 12860
rect 22480 12306 22508 12854
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22480 11898 22508 12242
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22848 11801 22876 15982
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23032 13870 23060 15642
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23032 13394 23060 13806
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23032 12986 23060 13330
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22834 11792 22890 11801
rect 22834 11727 22890 11736
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 9722 22508 10066
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22480 9625 22508 9658
rect 22466 9616 22522 9625
rect 22466 9551 22522 9560
rect 22848 8090 22876 11727
rect 23124 11218 23152 16050
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23216 15162 23244 15574
rect 23308 15473 23336 17478
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23294 15464 23350 15473
rect 23294 15399 23350 15408
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23584 12889 23612 14894
rect 23570 12880 23626 12889
rect 23570 12815 23626 12824
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12442 23704 12582
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23768 12345 23796 17070
rect 23860 14074 23888 23462
rect 24136 22545 24164 27526
rect 24398 27520 24454 27526
rect 25056 27526 25466 27554
rect 24950 26752 25006 26761
rect 24950 26687 25006 26696
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24964 23866 24992 26687
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25056 23730 25084 27526
rect 25410 27520 25466 27526
rect 26422 27520 26478 28000
rect 27434 27520 27490 28000
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25148 23866 25176 24210
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22808 24822 22817
rect 24766 22743 24822 22752
rect 24780 22710 24808 22743
rect 24768 22704 24820 22710
rect 25148 22681 25176 23802
rect 26436 22778 26464 27520
rect 27448 23798 27476 27520
rect 27618 25936 27674 25945
rect 27618 25871 27674 25880
rect 27632 24206 27660 25871
rect 27710 24576 27766 24585
rect 27710 24511 27766 24520
rect 27724 24410 27752 24511
rect 27712 24404 27764 24410
rect 27712 24346 27764 24352
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 24768 22646 24820 22652
rect 25134 22672 25190 22681
rect 25134 22607 25190 22616
rect 24122 22536 24178 22545
rect 24122 22471 24178 22480
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24766 21312 24822 21321
rect 24766 21247 24822 21256
rect 24780 21146 24808 21247
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 20946
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24674 20496 24730 20505
rect 24674 20431 24730 20440
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24688 18834 24716 20431
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24122 18592 24178 18601
rect 24122 18527 24178 18536
rect 24136 18222 24164 18527
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18770
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17785 24624 18022
rect 27618 17912 27674 17921
rect 27618 17847 27674 17856
rect 24582 17776 24638 17785
rect 24124 17740 24176 17746
rect 24582 17711 24638 17720
rect 24124 17682 24176 17688
rect 24136 17377 24164 17682
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24122 17368 24178 17377
rect 24289 17360 24585 17380
rect 24122 17303 24178 17312
rect 24136 17270 24164 17303
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24044 16794 24072 17138
rect 27632 16833 27660 17847
rect 24214 16824 24270 16833
rect 24032 16788 24084 16794
rect 24214 16759 24270 16768
rect 27618 16824 27674 16833
rect 27618 16759 27674 16768
rect 24032 16730 24084 16736
rect 24228 16658 24256 16759
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24136 15706 24164 16458
rect 24228 16182 24256 16594
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 16176 24268 16182
rect 24216 16118 24268 16124
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24780 15706 24808 15943
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 14822 24716 15506
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23754 12336 23810 12345
rect 23754 12271 23810 12280
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23492 10169 23520 11086
rect 23478 10160 23534 10169
rect 23478 10095 23534 10104
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 22940 9081 22968 9590
rect 22926 9072 22982 9081
rect 22926 9007 22982 9016
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23124 8634 23152 8978
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23860 5370 23888 5714
rect 22376 5364 22428 5370
rect 22376 5306 22428 5312
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23952 4185 23980 14758
rect 24950 14512 25006 14521
rect 24124 14476 24176 14482
rect 24950 14447 25006 14456
rect 24124 14418 24176 14424
rect 24136 13734 24164 14418
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24964 14074 24992 14447
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24136 13376 24164 13670
rect 24688 13394 24716 13806
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24780 13530 24808 13631
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24044 13348 24164 13376
rect 24216 13388 24268 13394
rect 24044 9625 24072 13348
rect 24216 13330 24268 13336
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24228 12646 24256 13330
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24122 12336 24178 12345
rect 24122 12271 24178 12280
rect 24136 10606 24164 12271
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24228 10130 24256 12582
rect 24766 12064 24822 12073
rect 24289 11996 24585 12016
rect 24766 11999 24822 12008
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 11999
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24596 11257 24624 11630
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24582 11248 24638 11257
rect 24582 11183 24638 11192
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24030 9616 24086 9625
rect 24030 9551 24086 9560
rect 24124 9580 24176 9586
rect 24044 8537 24072 9551
rect 24124 9522 24176 9528
rect 24136 9489 24164 9522
rect 24122 9480 24178 9489
rect 24122 9415 24178 9424
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24030 8528 24086 8537
rect 24030 8463 24086 8472
rect 22020 4126 22324 4154
rect 23938 4176 23994 4185
rect 22020 4078 22048 4126
rect 23938 4111 23994 4120
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 20626 54 20760 82
rect 21914 82 21970 480
rect 22020 82 22048 3062
rect 24044 2990 24072 8463
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24228 5166 24256 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 24214 2408 24270 2417
rect 24214 2343 24270 2352
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 21914 54 22048 82
rect 23032 82 23060 2246
rect 23294 82 23350 480
rect 23032 54 23350 82
rect 24228 82 24256 2343
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1057 24716 11494
rect 24766 10840 24822 10849
rect 24766 10775 24822 10784
rect 24780 10742 24808 10775
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 25226 5400 25282 5409
rect 25226 5335 25282 5344
rect 25240 3505 25268 5335
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 25594 4176 25650 4185
rect 25594 4111 25650 4120
rect 25226 3496 25282 3505
rect 25226 3431 25282 3440
rect 25240 2650 25268 3431
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 24674 1048 24730 1057
rect 24674 983 24730 992
rect 24582 82 24638 480
rect 24228 54 24638 82
rect 25608 82 25636 4111
rect 25962 82 26018 480
rect 25608 54 26018 82
rect 20626 0 20682 54
rect 21914 0 21970 54
rect 23294 0 23350 54
rect 24582 0 24638 54
rect 25962 0 26018 54
rect 27250 82 27306 480
rect 27356 82 27384 4966
rect 27618 3224 27674 3233
rect 27618 3159 27674 3168
rect 27632 3126 27660 3159
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 27632 1873 27660 2314
rect 27618 1864 27674 1873
rect 27618 1799 27674 1808
rect 27250 54 27384 82
rect 27250 0 27306 54
<< via2 >>
rect 110 25744 166 25800
rect 110 22752 166 22808
rect 1122 26696 1178 26752
rect 1582 23976 1638 24032
rect 110 19760 166 19816
rect 1950 21120 2006 21176
rect 2686 20984 2742 21040
rect 3790 20440 3846 20496
rect 3146 17584 3202 17640
rect 2134 16088 2190 16144
rect 110 12416 166 12472
rect 110 10920 166 10976
rect 110 8064 166 8120
rect 1490 9696 1546 9752
rect 1490 9560 1546 9616
rect 2134 14592 2190 14648
rect 2042 11192 2098 11248
rect 2226 9288 2282 9344
rect 2410 9560 2466 9616
rect 1766 6160 1822 6216
rect 1950 2624 2006 2680
rect 1582 1264 1638 1320
rect 3146 6296 3202 6352
rect 3974 19080 4030 19136
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 4434 18808 4490 18864
rect 4986 20440 5042 20496
rect 3882 16632 3938 16688
rect 3790 13368 3846 13424
rect 4250 16360 4306 16416
rect 4066 15000 4122 15056
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5446 19080 5502 19136
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5998 17992 6054 18048
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6090 17040 6146 17096
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 3514 8880 3570 8936
rect 5078 13776 5134 13832
rect 4710 11600 4766 11656
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5814 14864 5870 14920
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6274 19352 6330 19408
rect 6274 15952 6330 16008
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6090 13232 6146 13288
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 7470 21120 7526 21176
rect 6734 11192 6790 11248
rect 8298 20848 8354 20904
rect 7470 11056 7526 11112
rect 7930 10512 7986 10568
rect 8482 15564 8538 15600
rect 8482 15544 8484 15564
rect 8484 15544 8536 15564
rect 8536 15544 8538 15564
rect 8482 14592 8538 14648
rect 9402 23160 9458 23216
rect 9678 19352 9734 19408
rect 9494 18128 9550 18184
rect 9034 16088 9090 16144
rect 9310 14456 9366 14512
rect 7378 3848 7434 3904
rect 7654 3984 7710 4040
rect 7838 4120 7894 4176
rect 9862 17992 9918 18048
rect 9770 17584 9826 17640
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10230 24792 10286 24848
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10046 17992 10102 18048
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10782 16632 10838 16688
rect 11150 20476 11152 20496
rect 11152 20476 11204 20496
rect 11204 20476 11206 20496
rect 11150 20440 11206 20476
rect 11794 20440 11850 20496
rect 11886 19216 11942 19272
rect 11058 15000 11114 15056
rect 9034 12688 9090 12744
rect 9862 13232 9918 13288
rect 9862 12824 9918 12880
rect 9310 11056 9366 11112
rect 9494 8472 9550 8528
rect 10966 13776 11022 13832
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9310 6840 9366 6896
rect 9034 5480 9090 5536
rect 8298 4120 8354 4176
rect 8850 3032 8906 3088
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11426 13640 11482 13696
rect 11794 13368 11850 13424
rect 11518 7792 11574 7848
rect 12070 19216 12126 19272
rect 12346 16496 12402 16552
rect 12070 15952 12126 16008
rect 13174 18264 13230 18320
rect 14462 24792 14518 24848
rect 14554 19352 14610 19408
rect 13818 18672 13874 18728
rect 12162 13776 12218 13832
rect 12162 8472 12218 8528
rect 11426 3984 11482 4040
rect 11702 3440 11758 3496
rect 14094 16632 14150 16688
rect 13818 15544 13874 15600
rect 13726 15408 13782 15464
rect 13358 14320 13414 14376
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15198 20984 15254 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14830 18808 14886 18864
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14738 17176 14794 17232
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14646 16632 14702 16688
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14646 15952 14702 16008
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14738 13776 14794 13832
rect 14370 11736 14426 11792
rect 14186 11056 14242 11112
rect 14370 10512 14426 10568
rect 14094 8880 14150 8936
rect 15842 23160 15898 23216
rect 15750 22480 15806 22536
rect 15934 17720 15990 17776
rect 17222 18808 17278 18864
rect 16486 17040 16542 17096
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14830 10104 14886 10160
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14186 5072 14242 5128
rect 14554 5480 14610 5536
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 17406 18128 17462 18184
rect 17498 16632 17554 16688
rect 16578 12688 16634 12744
rect 15842 8880 15898 8936
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14462 3032 14518 3088
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16302 6160 16358 6216
rect 16946 9016 17002 9072
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 18694 22616 18750 22672
rect 18050 15952 18106 16008
rect 17590 11600 17646 11656
rect 17774 11192 17830 11248
rect 17682 9424 17738 9480
rect 16118 3984 16174 4040
rect 18234 16088 18290 16144
rect 18602 19216 18658 19272
rect 19062 19216 19118 19272
rect 18786 18264 18842 18320
rect 18602 16088 18658 16144
rect 18602 15272 18658 15328
rect 20350 23432 20406 23488
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20902 17176 20958 17232
rect 20074 16768 20130 16824
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19338 13776 19394 13832
rect 18510 12280 18566 12336
rect 18326 6296 18382 6352
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13640 19486 13696
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 18142 2352 18198 2408
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 21178 14320 21234 14376
rect 22282 18672 22338 18728
rect 21822 16496 21878 16552
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20810 6296 20866 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19982 3984 20038 4040
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22006 7792 22062 7848
rect 22834 16496 22890 16552
rect 23570 19216 23626 19272
rect 22834 11736 22890 11792
rect 22466 9560 22522 9616
rect 23294 15408 23350 15464
rect 23570 12824 23626 12880
rect 24950 26696 25006 26752
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22752 24822 22808
rect 27618 25880 27674 25936
rect 27710 24520 27766 24576
rect 25134 22616 25190 22672
rect 24122 22480 24178 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 21256 24822 21312
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24674 20440 24730 20496
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 18536 24178 18592
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 27618 17856 27674 17912
rect 24582 17720 24638 17776
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24122 17312 24178 17368
rect 24214 16768 24270 16824
rect 27618 16768 27674 16824
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24766 15952 24822 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23754 12280 23810 12336
rect 23478 10104 23534 10160
rect 22926 9016 22982 9072
rect 24950 14456 25006 14512
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 13640 24822 13696
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24122 12280 24178 12336
rect 24766 12008 24822 12064
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24582 11192 24638 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24030 9560 24086 9616
rect 24122 9424 24178 9480
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24030 8472 24086 8528
rect 23938 4120 23994 4176
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24214 2352 24270 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24766 10784 24822 10840
rect 25226 5344 25282 5400
rect 25594 4120 25650 4176
rect 25226 3440 25282 3496
rect 24674 992 24730 1048
rect 27618 3168 27674 3224
rect 27618 1808 27674 1864
<< metal3 >>
rect 0 27208 480 27328
rect 27520 27208 28000 27328
rect 62 26754 122 27208
rect 1117 26754 1183 26757
rect 62 26752 1183 26754
rect 62 26696 1122 26752
rect 1178 26696 1183 26752
rect 62 26694 1183 26696
rect 1117 26691 1183 26694
rect 24945 26754 25011 26757
rect 27662 26754 27722 27208
rect 24945 26752 27722 26754
rect 24945 26696 24950 26752
rect 25006 26696 27722 26752
rect 24945 26694 27722 26696
rect 24945 26691 25011 26694
rect 27520 25936 28000 25968
rect 27520 25880 27618 25936
rect 27674 25880 28000 25936
rect 27520 25848 28000 25880
rect 0 25800 480 25832
rect 0 25744 110 25800
rect 166 25744 480 25800
rect 0 25712 480 25744
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 10225 24850 10291 24853
rect 14457 24850 14523 24853
rect 14590 24850 14596 24852
rect 10225 24848 14596 24850
rect 10225 24792 10230 24848
rect 10286 24792 14462 24848
rect 14518 24792 14596 24848
rect 10225 24790 14596 24792
rect 10225 24787 10291 24790
rect 14457 24787 14523 24790
rect 14590 24788 14596 24790
rect 14660 24788 14666 24852
rect 27520 24576 28000 24608
rect 27520 24520 27710 24576
rect 27766 24520 28000 24576
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24520
rect 19610 24447 19930 24448
rect 0 24216 480 24336
rect 62 24034 122 24216
rect 1577 24034 1643 24037
rect 62 24032 1643 24034
rect 62 23976 1582 24032
rect 1638 23976 1643 24032
rect 62 23974 1643 23976
rect 1577 23971 1643 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 20345 23490 20411 23493
rect 20478 23490 20484 23492
rect 20345 23488 20484 23490
rect 20345 23432 20350 23488
rect 20406 23432 20484 23488
rect 20345 23430 20484 23432
rect 20345 23427 20411 23430
rect 20478 23428 20484 23430
rect 20548 23428 20554 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 9397 23218 9463 23221
rect 15837 23218 15903 23221
rect 9397 23216 15903 23218
rect 9397 23160 9402 23216
rect 9458 23160 15842 23216
rect 15898 23160 15903 23216
rect 9397 23158 15903 23160
rect 9397 23155 9463 23158
rect 15837 23155 15903 23158
rect 27520 23128 28000 23248
rect 5610 22880 5930 22881
rect 0 22808 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22752 110 22808
rect 166 22752 480 22808
rect 0 22720 480 22752
rect 24761 22810 24827 22813
rect 27662 22810 27722 23128
rect 24761 22808 27722 22810
rect 24761 22752 24766 22808
rect 24822 22752 27722 22808
rect 24761 22750 27722 22752
rect 24761 22747 24827 22750
rect 18689 22674 18755 22677
rect 25129 22674 25195 22677
rect 18689 22672 25195 22674
rect 18689 22616 18694 22672
rect 18750 22616 25134 22672
rect 25190 22616 25195 22672
rect 18689 22614 25195 22616
rect 18689 22611 18755 22614
rect 25129 22611 25195 22614
rect 15745 22538 15811 22541
rect 24117 22538 24183 22541
rect 15745 22536 24183 22538
rect 15745 22480 15750 22536
rect 15806 22480 24122 22536
rect 24178 22480 24183 22536
rect 15745 22478 24183 22480
rect 15745 22475 15811 22478
rect 24117 22475 24183 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21888
rect 24277 21727 24597 21728
rect 0 21224 480 21344
rect 24761 21314 24827 21317
rect 27662 21314 27722 21768
rect 24761 21312 27722 21314
rect 24761 21256 24766 21312
rect 24822 21256 27722 21312
rect 24761 21254 27722 21256
rect 24761 21251 24827 21254
rect 10277 21248 10597 21249
rect 62 20906 122 21224
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1945 21178 2011 21181
rect 7465 21178 7531 21181
rect 1945 21176 7531 21178
rect 1945 21120 1950 21176
rect 2006 21120 7470 21176
rect 7526 21120 7531 21176
rect 1945 21118 7531 21120
rect 1945 21115 2011 21118
rect 7465 21115 7531 21118
rect 2681 21042 2747 21045
rect 15193 21042 15259 21045
rect 2681 21040 15259 21042
rect 2681 20984 2686 21040
rect 2742 20984 15198 21040
rect 15254 20984 15259 21040
rect 2681 20982 15259 20984
rect 2681 20979 2747 20982
rect 15193 20979 15259 20982
rect 8293 20906 8359 20909
rect 62 20904 8359 20906
rect 62 20848 8298 20904
rect 8354 20848 8359 20904
rect 62 20846 8359 20848
rect 8293 20843 8359 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20636 28000 20664
rect 27520 20572 27660 20636
rect 27724 20572 28000 20636
rect 27520 20544 28000 20572
rect 3785 20498 3851 20501
rect 4981 20498 5047 20501
rect 11145 20498 11211 20501
rect 3785 20496 11211 20498
rect 3785 20440 3790 20496
rect 3846 20440 4986 20496
rect 5042 20440 11150 20496
rect 11206 20440 11211 20496
rect 3785 20438 11211 20440
rect 3785 20435 3851 20438
rect 4981 20435 5047 20438
rect 11145 20435 11211 20438
rect 11789 20498 11855 20501
rect 24669 20498 24735 20501
rect 11789 20496 27354 20498
rect 11789 20440 11794 20496
rect 11850 20440 24674 20496
rect 24730 20440 27354 20496
rect 11789 20438 27354 20440
rect 11789 20435 11855 20438
rect 24669 20435 24735 20438
rect 27294 20362 27354 20438
rect 27654 20362 27660 20364
rect 27294 20302 27660 20362
rect 27654 20300 27660 20302
rect 27724 20300 27730 20364
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19816 480 19848
rect 0 19760 110 19816
rect 166 19760 480 19816
rect 0 19728 480 19760
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 6269 19410 6335 19413
rect 9673 19410 9739 19413
rect 14549 19410 14615 19413
rect 6269 19408 14615 19410
rect 6269 19352 6274 19408
rect 6330 19352 9678 19408
rect 9734 19352 14554 19408
rect 14610 19352 14615 19408
rect 6269 19350 14615 19352
rect 6269 19347 6335 19350
rect 9673 19347 9739 19350
rect 14549 19347 14615 19350
rect 11881 19274 11947 19277
rect 12065 19274 12131 19277
rect 18597 19274 18663 19277
rect 11881 19272 18663 19274
rect 11881 19216 11886 19272
rect 11942 19216 12070 19272
rect 12126 19216 18602 19272
rect 18658 19216 18663 19272
rect 11881 19214 18663 19216
rect 11881 19211 11947 19214
rect 12065 19211 12131 19214
rect 18597 19211 18663 19214
rect 19057 19274 19123 19277
rect 23565 19274 23631 19277
rect 19057 19272 23631 19274
rect 19057 19216 19062 19272
rect 19118 19216 23570 19272
rect 23626 19216 23631 19272
rect 19057 19214 23631 19216
rect 19057 19211 19123 19214
rect 23565 19211 23631 19214
rect 27520 19184 28000 19304
rect 3969 19138 4035 19141
rect 5441 19138 5507 19141
rect 3969 19136 5507 19138
rect 3969 19080 3974 19136
rect 4030 19080 5446 19136
rect 5502 19080 5507 19136
rect 3969 19078 5507 19080
rect 3969 19075 4035 19078
rect 5441 19075 5507 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 4429 18866 4495 18869
rect 14825 18866 14891 18869
rect 17217 18866 17283 18869
rect 4429 18864 17283 18866
rect 4429 18808 4434 18864
rect 4490 18808 14830 18864
rect 14886 18808 17222 18864
rect 17278 18808 17283 18864
rect 4429 18806 17283 18808
rect 4429 18803 4495 18806
rect 14825 18803 14891 18806
rect 17217 18803 17283 18806
rect 13813 18730 13879 18733
rect 22277 18730 22343 18733
rect 27662 18730 27722 19184
rect 13813 18728 21466 18730
rect 13813 18672 13818 18728
rect 13874 18672 21466 18728
rect 13813 18670 21466 18672
rect 13813 18667 13879 18670
rect 21406 18594 21466 18670
rect 22277 18728 27722 18730
rect 22277 18672 22282 18728
rect 22338 18672 27722 18728
rect 22277 18670 27722 18672
rect 22277 18667 22343 18670
rect 24117 18594 24183 18597
rect 21406 18592 24183 18594
rect 21406 18536 24122 18592
rect 24178 18536 24183 18592
rect 21406 18534 24183 18536
rect 24117 18531 24183 18534
rect 5610 18528 5930 18529
rect 0 18368 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 62 18050 122 18368
rect 13169 18322 13235 18325
rect 18781 18322 18847 18325
rect 13169 18320 18847 18322
rect 13169 18264 13174 18320
rect 13230 18264 18786 18320
rect 18842 18264 18847 18320
rect 13169 18262 18847 18264
rect 13169 18259 13235 18262
rect 18781 18259 18847 18262
rect 9489 18186 9555 18189
rect 17401 18186 17467 18189
rect 9489 18184 17467 18186
rect 9489 18128 9494 18184
rect 9550 18128 17406 18184
rect 17462 18128 17467 18184
rect 9489 18126 17467 18128
rect 9489 18123 9555 18126
rect 17401 18123 17467 18126
rect 5993 18050 6059 18053
rect 62 18048 6059 18050
rect 62 17992 5998 18048
rect 6054 17992 6059 18048
rect 62 17990 6059 17992
rect 5993 17987 6059 17990
rect 9857 18050 9923 18053
rect 10041 18050 10107 18053
rect 9857 18048 10107 18050
rect 9857 17992 9862 18048
rect 9918 17992 10046 18048
rect 10102 17992 10107 18048
rect 9857 17990 10107 17992
rect 9857 17987 9923 17990
rect 10041 17987 10107 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 27520 17912 28000 17944
rect 27520 17856 27618 17912
rect 27674 17856 28000 17912
rect 27520 17824 28000 17856
rect 15929 17778 15995 17781
rect 24577 17778 24643 17781
rect 15929 17776 24643 17778
rect 15929 17720 15934 17776
rect 15990 17720 24582 17776
rect 24638 17720 24643 17776
rect 15929 17718 24643 17720
rect 15929 17715 15995 17718
rect 24577 17715 24643 17718
rect 3141 17642 3207 17645
rect 9765 17642 9831 17645
rect 3141 17640 9831 17642
rect 3141 17584 3146 17640
rect 3202 17584 9770 17640
rect 9826 17584 9831 17640
rect 3141 17582 9831 17584
rect 3141 17579 3207 17582
rect 9765 17579 9831 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 23422 17308 23428 17372
rect 23492 17370 23498 17372
rect 24117 17370 24183 17373
rect 23492 17368 24183 17370
rect 23492 17312 24122 17368
rect 24178 17312 24183 17368
rect 23492 17310 24183 17312
rect 23492 17308 23498 17310
rect 24117 17307 24183 17310
rect 14733 17234 14799 17237
rect 20897 17234 20963 17237
rect 14733 17232 20963 17234
rect 14733 17176 14738 17232
rect 14794 17176 20902 17232
rect 20958 17176 20963 17232
rect 14733 17174 20963 17176
rect 14733 17171 14799 17174
rect 20897 17171 20963 17174
rect 6085 17098 6151 17101
rect 16481 17098 16547 17101
rect 6085 17096 16547 17098
rect 6085 17040 6090 17096
rect 6146 17040 16486 17096
rect 16542 17040 16547 17096
rect 6085 17038 16547 17040
rect 6085 17035 6151 17038
rect 16481 17035 16547 17038
rect 0 16872 480 16992
rect 10277 16896 10597 16897
rect 62 16418 122 16872
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 20069 16826 20135 16829
rect 24209 16826 24275 16829
rect 27613 16826 27679 16829
rect 20069 16824 24275 16826
rect 20069 16768 20074 16824
rect 20130 16768 24214 16824
rect 24270 16768 24275 16824
rect 20069 16766 24275 16768
rect 20069 16763 20135 16766
rect 24209 16763 24275 16766
rect 27294 16824 27679 16826
rect 27294 16768 27618 16824
rect 27674 16768 27679 16824
rect 27294 16766 27679 16768
rect 3877 16690 3943 16693
rect 10777 16690 10843 16693
rect 3877 16688 10843 16690
rect 3877 16632 3882 16688
rect 3938 16632 10782 16688
rect 10838 16632 10843 16688
rect 3877 16630 10843 16632
rect 3877 16627 3943 16630
rect 10777 16627 10843 16630
rect 14089 16690 14155 16693
rect 14641 16690 14707 16693
rect 17493 16690 17559 16693
rect 27294 16690 27354 16766
rect 27613 16763 27679 16766
rect 14089 16688 27354 16690
rect 14089 16632 14094 16688
rect 14150 16632 14646 16688
rect 14702 16632 17498 16688
rect 17554 16632 27354 16688
rect 14089 16630 27354 16632
rect 14089 16627 14155 16630
rect 14641 16627 14707 16630
rect 17493 16627 17559 16630
rect 12341 16554 12407 16557
rect 21817 16554 21883 16557
rect 22829 16554 22895 16557
rect 12341 16552 22895 16554
rect 12341 16496 12346 16552
rect 12402 16496 21822 16552
rect 21878 16496 22834 16552
rect 22890 16496 22895 16552
rect 12341 16494 22895 16496
rect 12341 16491 12407 16494
rect 21817 16491 21883 16494
rect 22829 16491 22895 16494
rect 27520 16464 28000 16584
rect 4245 16418 4311 16421
rect 62 16416 4311 16418
rect 62 16360 4250 16416
rect 4306 16360 4311 16416
rect 62 16358 4311 16360
rect 4245 16355 4311 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2129 16146 2195 16149
rect 9029 16146 9095 16149
rect 18229 16146 18295 16149
rect 18597 16146 18663 16149
rect 2129 16144 18663 16146
rect 2129 16088 2134 16144
rect 2190 16088 9034 16144
rect 9090 16088 18234 16144
rect 18290 16088 18602 16144
rect 18658 16088 18663 16144
rect 2129 16086 18663 16088
rect 2129 16083 2195 16086
rect 9029 16083 9095 16086
rect 18229 16083 18295 16086
rect 18597 16083 18663 16086
rect 6269 16010 6335 16013
rect 6494 16010 6500 16012
rect 6269 16008 6500 16010
rect 6269 15952 6274 16008
rect 6330 15952 6500 16008
rect 6269 15950 6500 15952
rect 6269 15947 6335 15950
rect 6494 15948 6500 15950
rect 6564 15948 6570 16012
rect 12065 16010 12131 16013
rect 14641 16010 14707 16013
rect 12065 16008 14707 16010
rect 12065 15952 12070 16008
rect 12126 15952 14646 16008
rect 14702 15952 14707 16008
rect 12065 15950 14707 15952
rect 12065 15947 12131 15950
rect 14641 15947 14707 15950
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 18045 16010 18111 16013
rect 17972 16008 18111 16010
rect 17972 15952 18050 16008
rect 18106 15952 18111 16008
rect 17972 15950 18111 15952
rect 17972 15948 17978 15950
rect 18045 15947 18111 15950
rect 24761 16010 24827 16013
rect 27662 16010 27722 16464
rect 24761 16008 27722 16010
rect 24761 15952 24766 16008
rect 24822 15952 27722 16008
rect 24761 15950 27722 15952
rect 24761 15947 24827 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 8477 15602 8543 15605
rect 13813 15602 13879 15605
rect 8477 15600 13879 15602
rect 8477 15544 8482 15600
rect 8538 15544 13818 15600
rect 13874 15544 13879 15600
rect 8477 15542 13879 15544
rect 8477 15539 8543 15542
rect 13813 15539 13879 15542
rect 0 15376 480 15496
rect 13721 15466 13787 15469
rect 23289 15466 23355 15469
rect 13721 15464 23355 15466
rect 13721 15408 13726 15464
rect 13782 15408 23294 15464
rect 23350 15408 23355 15464
rect 13721 15406 23355 15408
rect 13721 15403 13787 15406
rect 23289 15403 23355 15406
rect 23430 15406 27722 15466
rect 62 14922 122 15376
rect 18597 15330 18663 15333
rect 23430 15330 23490 15406
rect 18597 15328 23490 15330
rect 18597 15272 18602 15328
rect 18658 15272 23490 15328
rect 18597 15270 23490 15272
rect 18597 15267 18663 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 27662 15224 27722 15406
rect 24277 15199 24597 15200
rect 27520 15104 28000 15224
rect 4061 15058 4127 15061
rect 11053 15058 11119 15061
rect 4061 15056 11119 15058
rect 4061 15000 4066 15056
rect 4122 15000 11058 15056
rect 11114 15000 11119 15056
rect 4061 14998 11119 15000
rect 4061 14995 4127 14998
rect 11053 14995 11119 14998
rect 5809 14922 5875 14925
rect 62 14920 5875 14922
rect 62 14864 5814 14920
rect 5870 14864 5875 14920
rect 62 14862 5875 14864
rect 5809 14859 5875 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 2129 14650 2195 14653
rect 8477 14650 8543 14653
rect 2129 14648 8543 14650
rect 2129 14592 2134 14648
rect 2190 14592 8482 14648
rect 8538 14592 8543 14648
rect 2129 14590 8543 14592
rect 2129 14587 2195 14590
rect 8477 14587 8543 14590
rect 9305 14514 9371 14517
rect 24945 14514 25011 14517
rect 9305 14512 25011 14514
rect 9305 14456 9310 14512
rect 9366 14456 24950 14512
rect 25006 14456 25011 14512
rect 9305 14454 25011 14456
rect 9305 14451 9371 14454
rect 24945 14451 25011 14454
rect 13353 14378 13419 14381
rect 21173 14378 21239 14381
rect 13353 14376 21239 14378
rect 13353 14320 13358 14376
rect 13414 14320 21178 14376
rect 21234 14320 21239 14376
rect 13353 14318 21239 14320
rect 13353 14315 13419 14318
rect 21173 14315 21239 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13880 480 14000
rect 27520 13880 28000 14000
rect 62 13290 122 13880
rect 5073 13834 5139 13837
rect 10961 13834 11027 13837
rect 12157 13834 12223 13837
rect 5073 13832 12223 13834
rect 5073 13776 5078 13832
rect 5134 13776 10966 13832
rect 11022 13776 12162 13832
rect 12218 13776 12223 13832
rect 5073 13774 12223 13776
rect 5073 13771 5139 13774
rect 10961 13771 11027 13774
rect 12157 13771 12223 13774
rect 14733 13834 14799 13837
rect 19333 13834 19399 13837
rect 14733 13832 19399 13834
rect 14733 13776 14738 13832
rect 14794 13776 19338 13832
rect 19394 13776 19399 13832
rect 14733 13774 19399 13776
rect 14733 13771 14799 13774
rect 19333 13771 19399 13774
rect 11421 13698 11487 13701
rect 19425 13698 19491 13701
rect 11421 13696 19491 13698
rect 11421 13640 11426 13696
rect 11482 13640 19430 13696
rect 19486 13640 19491 13696
rect 11421 13638 19491 13640
rect 11421 13635 11487 13638
rect 19425 13635 19491 13638
rect 24761 13698 24827 13701
rect 27662 13698 27722 13880
rect 24761 13696 27722 13698
rect 24761 13640 24766 13696
rect 24822 13640 27722 13696
rect 24761 13638 27722 13640
rect 24761 13635 24827 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3785 13426 3851 13429
rect 11789 13426 11855 13429
rect 3785 13424 11855 13426
rect 3785 13368 3790 13424
rect 3846 13368 11794 13424
rect 11850 13368 11855 13424
rect 3785 13366 11855 13368
rect 3785 13363 3851 13366
rect 11789 13363 11855 13366
rect 6085 13290 6151 13293
rect 9857 13290 9923 13293
rect 62 13288 9923 13290
rect 62 13232 6090 13288
rect 6146 13232 9862 13288
rect 9918 13232 9923 13288
rect 62 13230 9923 13232
rect 6085 13227 6151 13230
rect 9857 13227 9923 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 9857 12882 9923 12885
rect 23565 12882 23631 12885
rect 9857 12880 23631 12882
rect 9857 12824 9862 12880
rect 9918 12824 23570 12880
rect 23626 12824 23631 12880
rect 9857 12822 23631 12824
rect 9857 12819 9923 12822
rect 23565 12819 23631 12822
rect 9029 12746 9095 12749
rect 16573 12746 16639 12749
rect 9029 12744 16639 12746
rect 9029 12688 9034 12744
rect 9090 12688 16578 12744
rect 16634 12688 16639 12744
rect 9029 12686 16639 12688
rect 9029 12683 9095 12686
rect 16573 12683 16639 12686
rect 10277 12544 10597 12545
rect 0 12472 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12640
rect 19610 12479 19930 12480
rect 0 12416 110 12472
rect 166 12416 480 12472
rect 0 12384 480 12416
rect 18505 12338 18571 12341
rect 23749 12338 23815 12341
rect 24117 12338 24183 12341
rect 18505 12336 24183 12338
rect 18505 12280 18510 12336
rect 18566 12280 23754 12336
rect 23810 12280 24122 12336
rect 24178 12280 24183 12336
rect 18505 12278 24183 12280
rect 18505 12275 18571 12278
rect 23749 12275 23815 12278
rect 24117 12275 24183 12278
rect 24761 12066 24827 12069
rect 27662 12066 27722 12520
rect 24761 12064 27722 12066
rect 24761 12008 24766 12064
rect 24822 12008 27722 12064
rect 24761 12006 27722 12008
rect 24761 12003 24827 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 14365 11794 14431 11797
rect 22829 11794 22895 11797
rect 14365 11792 22895 11794
rect 14365 11736 14370 11792
rect 14426 11736 22834 11792
rect 22890 11736 22895 11792
rect 14365 11734 22895 11736
rect 14365 11731 14431 11734
rect 22829 11731 22895 11734
rect 4705 11658 4771 11661
rect 17585 11658 17651 11661
rect 4705 11656 17651 11658
rect 4705 11600 4710 11656
rect 4766 11600 17590 11656
rect 17646 11600 17651 11656
rect 4705 11598 17651 11600
rect 4705 11595 4771 11598
rect 17585 11595 17651 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2037 11250 2103 11253
rect 6729 11250 6795 11253
rect 17769 11250 17835 11253
rect 24577 11250 24643 11253
rect 2037 11248 17835 11250
rect 2037 11192 2042 11248
rect 2098 11192 6734 11248
rect 6790 11192 17774 11248
rect 17830 11192 17835 11248
rect 2037 11190 17835 11192
rect 2037 11187 2103 11190
rect 6729 11187 6795 11190
rect 17769 11187 17835 11190
rect 19198 11248 24643 11250
rect 19198 11192 24582 11248
rect 24638 11192 24643 11248
rect 19198 11190 24643 11192
rect 7465 11114 7531 11117
rect 9305 11114 9371 11117
rect 14181 11114 14247 11117
rect 19198 11114 19258 11190
rect 24577 11187 24643 11190
rect 27520 11160 28000 11280
rect 7465 11112 19258 11114
rect 7465 11056 7470 11112
rect 7526 11056 9310 11112
rect 9366 11056 14186 11112
rect 14242 11056 19258 11112
rect 7465 11054 19258 11056
rect 7465 11051 7531 11054
rect 9305 11051 9371 11054
rect 14181 11051 14247 11054
rect 0 10976 480 11008
rect 0 10920 110 10976
rect 166 10920 480 10976
rect 0 10888 480 10920
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 24761 10842 24827 10845
rect 27662 10842 27722 11160
rect 24761 10840 27722 10842
rect 24761 10784 24766 10840
rect 24822 10784 27722 10840
rect 24761 10782 27722 10784
rect 24761 10779 24827 10782
rect 7925 10570 7991 10573
rect 14365 10570 14431 10573
rect 7925 10568 14431 10570
rect 7925 10512 7930 10568
rect 7986 10512 14370 10568
rect 14426 10512 14431 10568
rect 7925 10510 14431 10512
rect 7925 10507 7991 10510
rect 14365 10507 14431 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 14825 10162 14891 10165
rect 23473 10162 23539 10165
rect 14825 10160 23539 10162
rect 14825 10104 14830 10160
rect 14886 10104 23478 10160
rect 23534 10104 23539 10160
rect 14825 10102 23539 10104
rect 14825 10099 14891 10102
rect 23473 10099 23539 10102
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27520 9800 28000 9920
rect 24277 9759 24597 9760
rect 1485 9754 1551 9757
rect 614 9752 1551 9754
rect 614 9696 1490 9752
rect 1546 9696 1551 9752
rect 614 9694 1551 9696
rect 614 9690 674 9694
rect 1485 9691 1551 9694
rect 62 9648 674 9690
rect 0 9630 674 9648
rect 0 9528 480 9630
rect 1485 9618 1551 9621
rect 2405 9618 2471 9621
rect 22461 9618 22527 9621
rect 1485 9616 22527 9618
rect 1485 9560 1490 9616
rect 1546 9560 2410 9616
rect 2466 9560 22466 9616
rect 22522 9560 22527 9616
rect 1485 9558 22527 9560
rect 1485 9555 1551 9558
rect 2405 9555 2471 9558
rect 22461 9555 22527 9558
rect 24025 9618 24091 9621
rect 27662 9618 27722 9800
rect 24025 9616 27722 9618
rect 24025 9560 24030 9616
rect 24086 9560 27722 9616
rect 24025 9558 27722 9560
rect 24025 9555 24091 9558
rect 17677 9482 17743 9485
rect 4110 9480 17743 9482
rect 4110 9424 17682 9480
rect 17738 9424 17743 9480
rect 4110 9422 17743 9424
rect 2221 9346 2287 9349
rect 4110 9346 4170 9422
rect 17677 9419 17743 9422
rect 20478 9420 20484 9484
rect 20548 9482 20554 9484
rect 24117 9482 24183 9485
rect 20548 9480 24183 9482
rect 20548 9424 24122 9480
rect 24178 9424 24183 9480
rect 20548 9422 24183 9424
rect 20548 9420 20554 9422
rect 24117 9419 24183 9422
rect 2221 9344 4170 9346
rect 2221 9288 2226 9344
rect 2282 9288 4170 9344
rect 2221 9286 4170 9288
rect 2221 9283 2287 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 16941 9074 17007 9077
rect 22921 9074 22987 9077
rect 16941 9072 22987 9074
rect 16941 9016 16946 9072
rect 17002 9016 22926 9072
rect 22982 9016 22987 9072
rect 16941 9014 22987 9016
rect 16941 9011 17007 9014
rect 22921 9011 22987 9014
rect 3509 8938 3575 8941
rect 14089 8938 14155 8941
rect 15837 8938 15903 8941
rect 3509 8936 15903 8938
rect 3509 8880 3514 8936
rect 3570 8880 14094 8936
rect 14150 8880 15842 8936
rect 15898 8880 15903 8936
rect 3509 8878 15903 8880
rect 3509 8875 3575 8878
rect 14089 8875 14155 8878
rect 15837 8875 15903 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 9489 8530 9555 8533
rect 12157 8530 12223 8533
rect 24025 8530 24091 8533
rect 9489 8528 24091 8530
rect 9489 8472 9494 8528
rect 9550 8472 12162 8528
rect 12218 8472 24030 8528
rect 24086 8472 24091 8528
rect 9489 8470 24091 8472
rect 9489 8467 9555 8470
rect 12157 8467 12223 8470
rect 24025 8467 24091 8470
rect 27520 8532 28000 8560
rect 27520 8468 27660 8532
rect 27724 8468 28000 8532
rect 27520 8440 28000 8468
rect 10277 8192 10597 8193
rect 0 8120 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 0 8064 110 8120
rect 166 8064 480 8120
rect 0 8032 480 8064
rect 11513 7850 11579 7853
rect 11646 7850 11652 7852
rect 11513 7848 11652 7850
rect 11513 7792 11518 7848
rect 11574 7792 11652 7848
rect 11513 7790 11652 7792
rect 11513 7787 11579 7790
rect 11646 7788 11652 7790
rect 11716 7788 11722 7852
rect 22001 7850 22067 7853
rect 22001 7848 27722 7850
rect 22001 7792 22006 7848
rect 22062 7792 27722 7848
rect 22001 7790 27722 7792
rect 22001 7787 22067 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27662 7336 27722 7790
rect 27520 7216 28000 7336
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 54 6836 60 6900
rect 124 6898 130 6900
rect 9305 6898 9371 6901
rect 124 6896 9371 6898
rect 124 6840 9310 6896
rect 9366 6840 9371 6896
rect 124 6838 9371 6840
rect 124 6836 130 6838
rect 9305 6835 9371 6838
rect 0 6628 480 6656
rect 0 6564 60 6628
rect 124 6564 480 6628
rect 0 6536 480 6564
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 3141 6354 3207 6357
rect 18321 6354 18387 6357
rect 20805 6354 20871 6357
rect 3141 6352 20871 6354
rect 3141 6296 3146 6352
rect 3202 6296 18326 6352
rect 18382 6296 20810 6352
rect 20866 6296 20871 6352
rect 3141 6294 20871 6296
rect 3141 6291 3207 6294
rect 18321 6291 18387 6294
rect 20805 6291 20871 6294
rect 1761 6218 1827 6221
rect 16297 6218 16363 6221
rect 1761 6216 16363 6218
rect 1761 6160 1766 6216
rect 1822 6160 16302 6216
rect 16358 6160 16363 6216
rect 1761 6158 16363 6160
rect 1761 6155 1827 6158
rect 16297 6155 16363 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 27520 5856 28000 5976
rect 9029 5538 9095 5541
rect 14549 5538 14615 5541
rect 9029 5536 14615 5538
rect 9029 5480 9034 5536
rect 9090 5480 14554 5536
rect 14610 5480 14615 5536
rect 9029 5478 14615 5480
rect 9029 5475 9095 5478
rect 14549 5475 14615 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 25221 5402 25287 5405
rect 27662 5402 27722 5856
rect 25221 5400 27722 5402
rect 25221 5344 25226 5400
rect 25282 5344 27722 5400
rect 25221 5342 27722 5344
rect 25221 5339 25287 5342
rect 0 5132 480 5160
rect 0 5068 60 5132
rect 124 5068 480 5132
rect 14181 5130 14247 5133
rect 0 5040 480 5068
rect 9630 5128 14247 5130
rect 9630 5072 14186 5128
rect 14242 5072 14247 5128
rect 9630 5070 14247 5072
rect 54 4796 60 4860
rect 124 4858 130 4860
rect 9630 4858 9690 5070
rect 14181 5067 14247 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 124 4798 9690 4858
rect 124 4796 130 4798
rect 27520 4496 28000 4616
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7833 4178 7899 4181
rect 8293 4178 8359 4181
rect 23933 4178 23999 4181
rect 25589 4178 25655 4181
rect 7833 4176 8359 4178
rect 7833 4120 7838 4176
rect 7894 4120 8298 4176
rect 8354 4120 8359 4176
rect 7833 4118 8359 4120
rect 7833 4115 7899 4118
rect 8293 4115 8359 4118
rect 19290 4176 25655 4178
rect 19290 4120 23938 4176
rect 23994 4120 25594 4176
rect 25650 4120 25655 4176
rect 19290 4118 25655 4120
rect 7649 4042 7715 4045
rect 11421 4042 11487 4045
rect 7649 4040 11487 4042
rect 7649 3984 7654 4040
rect 7710 3984 11426 4040
rect 11482 3984 11487 4040
rect 7649 3982 11487 3984
rect 7649 3979 7715 3982
rect 11421 3979 11487 3982
rect 16113 4042 16179 4045
rect 19290 4042 19350 4118
rect 23933 4115 23999 4118
rect 25589 4115 25655 4118
rect 16113 4040 19350 4042
rect 16113 3984 16118 4040
rect 16174 3984 19350 4040
rect 16113 3982 19350 3984
rect 19977 4042 20043 4045
rect 27662 4042 27722 4496
rect 19977 4040 27722 4042
rect 19977 3984 19982 4040
rect 20038 3984 27722 4040
rect 19977 3982 27722 3984
rect 16113 3979 16179 3982
rect 19977 3979 20043 3982
rect 7373 3906 7439 3909
rect 62 3904 7439 3906
rect 62 3848 7378 3904
rect 7434 3848 7439 3904
rect 62 3846 7439 3848
rect 62 3664 122 3846
rect 7373 3843 7439 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3544 480 3664
rect 11697 3498 11763 3501
rect 25221 3498 25287 3501
rect 11697 3496 25287 3498
rect 11697 3440 11702 3496
rect 11758 3440 25226 3496
rect 25282 3440 25287 3496
rect 11697 3438 25287 3440
rect 11697 3435 11763 3438
rect 25221 3435 25287 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27520 3224 28000 3256
rect 27520 3168 27618 3224
rect 27674 3168 28000 3224
rect 27520 3136 28000 3168
rect 8845 3090 8911 3093
rect 14457 3090 14523 3093
rect 8845 3088 14523 3090
rect 8845 3032 8850 3088
rect 8906 3032 14462 3088
rect 14518 3032 14523 3088
rect 8845 3030 14523 3032
rect 8845 3027 8911 3030
rect 14457 3027 14523 3030
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 1945 2682 2011 2685
rect 62 2680 2011 2682
rect 62 2624 1950 2680
rect 2006 2624 2011 2680
rect 62 2622 2011 2624
rect 62 2168 122 2622
rect 1945 2619 2011 2622
rect 18137 2410 18203 2413
rect 24209 2410 24275 2413
rect 18137 2408 24275 2410
rect 18137 2352 18142 2408
rect 18198 2352 24214 2408
rect 24270 2352 24275 2408
rect 18137 2350 24275 2352
rect 18137 2347 18203 2350
rect 24209 2347 24275 2350
rect 5610 2208 5930 2209
rect 0 2048 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 27520 1864 28000 1896
rect 27520 1808 27618 1864
rect 27674 1808 28000 1864
rect 27520 1776 28000 1808
rect 1577 1322 1643 1325
rect 62 1320 1643 1322
rect 62 1264 1582 1320
rect 1638 1264 1643 1320
rect 62 1262 1643 1264
rect 62 808 122 1262
rect 1577 1259 1643 1262
rect 24669 1050 24735 1053
rect 24669 1048 27722 1050
rect 24669 992 24674 1048
rect 24730 992 27722 1048
rect 24669 990 27722 992
rect 24669 987 24735 990
rect 0 688 480 808
rect 27662 672 27722 990
rect 27520 552 28000 672
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 14596 24788 14660 24852
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 20484 23428 20548 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 27660 20572 27724 20636
rect 27660 20300 27724 20364
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 23428 17308 23492 17372
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 6500 15948 6564 16012
rect 17908 15948 17972 16012
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 20484 9420 20548 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 27660 8468 27724 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 11652 7788 11716 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 60 6836 124 6900
rect 60 6564 124 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 60 5068 124 5132
rect 60 4796 124 4860
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14595 24852 14661 24853
rect 14595 24788 14596 24852
rect 14660 24788 14661 24852
rect 14595 24787 14661 24788
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 14598 17458 14658 24787
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 59 6900 125 6901
rect 59 6836 60 6900
rect 124 6836 125 6900
rect 59 6835 125 6836
rect 62 6629 122 6835
rect 59 6628 125 6629
rect 59 6564 60 6628
rect 124 6564 125 6628
rect 59 6563 125 6564
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 59 5132 125 5133
rect 59 5068 60 5132
rect 124 5068 125 5132
rect 59 5067 125 5068
rect 62 4861 122 5067
rect 59 4860 125 4861
rect 59 4796 60 4860
rect 124 4796 125 4860
rect 59 4795 125 4796
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 20483 23492 20549 23493
rect 20483 23428 20484 23492
rect 20548 23428 20549 23492
rect 20483 23427 20549 23428
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 20486 9485 20546 23427
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 27659 20636 27725 20637
rect 27659 20572 27660 20636
rect 27724 20572 27725 20636
rect 27659 20571 27725 20572
rect 27662 20365 27722 20571
rect 27659 20364 27725 20365
rect 27659 20300 27660 20364
rect 27724 20300 27725 20364
rect 27659 20299 27725 20300
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 20483 9484 20549 9485
rect 20483 9420 20484 9484
rect 20548 9420 20549 9484
rect 20483 9419 20549 9420
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 27659 8532 27725 8533
rect 27659 8468 27660 8532
rect 27724 8468 27725 8532
rect 27659 8467 27725 8468
rect 27662 7938 27722 8467
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 14510 17222 14746 17458
rect 6414 16012 6650 16098
rect 6414 15948 6500 16012
rect 6500 15948 6564 16012
rect 6564 15948 6650 16012
rect 6414 15862 6650 15948
rect 17822 16012 18058 16098
rect 17822 15948 17908 16012
rect 17908 15948 17972 16012
rect 17972 15948 18058 16012
rect 17822 15862 18058 15948
rect 11566 7852 11802 7938
rect 11566 7788 11652 7852
rect 11652 7788 11716 7852
rect 11716 7788 11802 7852
rect 11566 7702 11802 7788
rect 23342 17372 23578 17458
rect 23342 17308 23428 17372
rect 23428 17308 23492 17372
rect 23492 17308 23578 17372
rect 23342 17222 23578 17308
rect 27574 7702 27810 7938
<< metal5 >>
rect 14468 17458 23620 17500
rect 14468 17222 14510 17458
rect 14746 17222 23342 17458
rect 23578 17222 23620 17458
rect 14468 17180 23620 17222
rect 6372 16098 18100 16140
rect 6372 15862 6414 16098
rect 6650 15862 17822 16098
rect 18058 15862 18100 16098
rect 6372 15820 18100 15862
rect 11524 7938 27852 7980
rect 11524 7702 11566 7938
rect 11802 7702 27574 7938
rect 27810 7702 27852 7938
rect 11524 7660 27852 7702
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_buf_2  _179_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_53
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_61 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_68
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_72
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 774 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_79
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_118 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_120
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_0_152
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_145
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_169
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_169
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_192
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_200
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_212
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_224
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_224
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _178_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_85
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_139
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_170
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_35
timestamp 1586364061
transform 1 0 4324 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_89
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_62
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_4_77
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_52
timestamp 1586364061
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_65
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_85
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_151
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_155
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_190
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_194
timestamp 1586364061
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_222
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_28
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_111
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_122
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_140
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_144
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_197
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_241
timestamp 1586364061
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_246
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_or2_4  _050_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 682 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_53
timestamp 1586364061
transform 1 0 5980 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_85
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_180
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_188
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_248
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_or2_4  _113_
timestamp 1586364061
transform 1 0 1472 0 1 7072
box -38 -48 682 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _162_
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _164_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_195
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_11
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_37
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_162
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_236
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_248
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_260
timestamp 1586364061
transform 1 0 25024 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_or4_4  _076_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__D
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_72
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_76
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_165
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_222
timestamp 1586364061
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_273
timestamp 1586364061
transform 1 0 26220 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_65
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_69
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_184
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_235
timestamp 1586364061
transform 1 0 22724 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_45
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_238
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_248
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_252
timestamp 1586364061
transform 1 0 24288 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_264
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_nand2_4  _085_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_131
timestamp 1586364061
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _048_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 4140 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_42
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_50
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_16_140
timestamp 1586364061
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 774 592
use scs8hd_conb_1  _161_
timestamp 1586364061
transform 1 0 23460 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_246
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_258
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_113
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_157
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_210
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_227
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_231
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_234
timestamp 1586364061
transform 1 0 22632 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_242
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__C
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__067__D
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_55
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_78
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_82
timestamp 1586364061
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_96
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_100
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_160
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_224
timestamp 1586364061
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_258
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_270
timestamp 1586364061
transform 1 0 25944 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_274
timestamp 1586364061
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _132_
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 866 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _067_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_30
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__132__C
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_85
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_109
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_122
timestamp 1586364061
transform 1 0 12328 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_150
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_209
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_234
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_238
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_241
timestamp 1586364061
transform 1 0 23276 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _166_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_253
timestamp 1586364061
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_17
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 4876 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_50
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_54
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_58
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 11868 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_233
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_237
timestamp 1586364061
transform 1 0 22908 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_77
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_130
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_133
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use scs8hd_nor2_4  _083_
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_180
timestamp 1586364061
transform 1 0 17664 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_197
timestamp 1586364061
transform 1 0 19228 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_235
timestamp 1586364061
transform 1 0 22724 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_246
timestamp 1586364061
transform 1 0 23736 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_or4_4  _086_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_or4_4  _114_
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_37
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_41
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_205
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_234
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_238
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_242
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_or4_4  _051_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_53
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_72
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_113
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_134
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_138
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_224
timestamp 1586364061
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_228
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 774 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_13
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_26
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_30
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_46
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_50
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_54
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_58
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_164
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_212
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_216
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_238
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_248
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__D
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__D
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_17
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_78
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_87
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_141
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_155
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_176
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_182
timestamp 1586364061
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_189
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_228
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_241
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_248
timestamp 1586364061
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_252
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_256
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_268
timestamp 1586364061
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_270
timestamp 1586364061
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_276
timestamp 1586364061
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_10
timestamp 1586364061
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_55
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_89
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_158
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_173
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _060_
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_203
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_207
timestamp 1586364061
transform 1 0 20148 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_252
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_264
timestamp 1586364061
transform 1 0 25392 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_272
timestamp 1586364061
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_20
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_24
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_28
timestamp 1586364061
transform 1 0 3680 0 1 17952
box -38 -48 130 592
use scs8hd_conb_1  _163_
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_167
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_189
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_230
timestamp 1586364061
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_248
timestamp 1586364061
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_252
timestamp 1586364061
transform 1 0 24288 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _168_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use scs8hd_or3_4  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _062_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_184
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _054_
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_241
timestamp 1586364061
transform 1 0 23276 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_252
timestamp 1586364061
transform 1 0 24288 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_264
timestamp 1586364061
transform 1 0 25392 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_272
timestamp 1586364061
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_or3_4  _061_
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__C
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_77
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_166
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_177
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_213
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_226
timestamp 1586364061
transform 1 0 21896 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_238
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use scs8hd_conb_1  _169_
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_248
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_260
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_272
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_12
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_or3_4  _055_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use scs8hd_or3_4  _059_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_29
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_41
timestamp 1586364061
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_50
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_54
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _167_
timestamp 1586364061
transform 1 0 8188 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_85
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_89
timestamp 1586364061
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_131
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_135
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_167
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_184
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_191
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_228
timestamp 1586364061
transform 1 0 22080 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _052_
timestamp 1586364061
transform 1 0 22448 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_32_241
timestamp 1586364061
transform 1 0 23276 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_253
timestamp 1586364061
transform 1 0 24380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_265
timestamp 1586364061
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_273
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_10
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_or3_4  _057_
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 866 592
use scs8hd_or3_4  _053_
timestamp 1586364061
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__C
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__C
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 406 592
use scs8hd_or3_4  _063_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_or3_4  _065_
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_29
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_54
timestamp 1586364061
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_58
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_71
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_75
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_79
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_134
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_151
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_157
timestamp 1586364061
transform 1 0 15548 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_161
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_177
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _058_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_216
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _056_
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_233
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_235
timestamp 1586364061
transform 1 0 22724 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_259
timestamp 1586364061
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_28
timestamp 1586364061
transform 1 0 3680 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_34
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_81
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_99
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_116
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_126
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_151
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_155
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_178
timestamp 1586364061
transform 1 0 17480 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_188
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_192
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_207
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_224
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_228
timestamp 1586364061
transform 1 0 22080 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_11
timestamp 1586364061
transform 1 0 2116 0 -1 22304
box -38 -48 130 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_43
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_51
timestamp 1586364061
transform 1 0 5796 0 -1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_67
timestamp 1586364061
transform 1 0 7268 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_70
timestamp 1586364061
transform 1 0 7544 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_150
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_167
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_179
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17664 0 -1 22304
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_195
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_198
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_203
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_236
timestamp 1586364061
transform 1 0 22816 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_248
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_260
timestamp 1586364061
transform 1 0 25024 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_272
timestamp 1586364061
transform 1 0 26128 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2668 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_28
timestamp 1586364061
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_32
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_45
timestamp 1586364061
transform 1 0 5244 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_96
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_37_140
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_157
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_174
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_178
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_195
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_223
timestamp 1586364061
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_275
timestamp 1586364061
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_52
timestamp 1586364061
transform 1 0 5888 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_60
timestamp 1586364061
transform 1 0 6624 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_81
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_85
timestamp 1586364061
transform 1 0 8924 0 -1 23392
box -38 -48 590 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 10028 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_131
timestamp 1586364061
transform 1 0 13156 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 17112 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  FILLER_38_171
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_183
timestamp 1586364061
transform 1 0 17940 0 -1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_194
timestamp 1586364061
transform 1 0 18952 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _165_
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_33
timestamp 1586364061
transform 1 0 4140 0 1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_49
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_62
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_68
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_72
timestamp 1586364061
transform 1 0 7728 0 1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_73
timestamp 1586364061
transform 1 0 7820 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_80
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_90
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_109
timestamp 1586364061
transform 1 0 11132 0 -1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_132
timestamp 1586364061
transform 1 0 13248 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_153
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_162
timestamp 1586364061
transform 1 0 16008 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 16468 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_171
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_181
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_195
timestamp 1586364061
transform 1 0 19044 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_207
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23000 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_241
timestamp 1586364061
transform 1 0 23276 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_253
timestamp 1586364061
transform 1 0 24380 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_85
timestamp 1586364061
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_89
timestamp 1586364061
transform 1 0 9292 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_96
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_100
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_104
timestamp 1586364061
transform 1 0 10672 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_134
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_138
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 406 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_145
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_149
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_157
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_161
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_173
timestamp 1586364061
transform 1 0 17020 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_181
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_100
timestamp 1586364061
transform 1 0 10304 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_111
timestamp 1586364061
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_123
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_136
timestamp 1586364061
transform 1 0 13616 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_147
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 478 27520 534 28000 6 address[0]
port 0 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 address[1]
port 1 nsew default input
rlabel metal2 s 3238 0 3294 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 2410 27520 2466 28000 6 address[3]
port 3 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 688 480 808 6 address[5]
port 5 nsew default input
rlabel metal3 s 0 2048 480 2168 6 address[6]
port 6 nsew default input
rlabel metal2 s 4618 0 4674 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 0 3544 480 3664 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 4434 27520 4490 28000 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal2 s 5446 27520 5502 28000 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 27520 552 28000 672 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 7286 0 7342 480 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 27520 1776 28000 1896 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 8574 0 8630 480 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 6458 27520 6514 28000 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 27520 3136 28000 3256 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 27520 4496 28000 4616 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 11242 0 11298 480 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 5856 28000 5976 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 27520 9800 28000 9920 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal2 s 7470 27520 7526 28000 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal2 s 15290 0 15346 480 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 8390 27520 8446 28000 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 9402 27520 9458 28000 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 12438 27520 12494 28000 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal2 s 13450 27520 13506 28000 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 14462 27520 14518 28000 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 15382 27520 15438 28000 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal2 s 16394 27520 16450 28000 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 18418 27520 18474 28000 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal3 s 27520 16464 28000 16584 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 23294 0 23350 480 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 19430 27520 19486 28000 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chany_top_in[0]
port 63 nsew default input
rlabel metal2 s 20442 27520 20498 28000 6 chany_top_in[1]
port 64 nsew default input
rlabel metal3 s 27520 19184 28000 19304 6 chany_top_in[2]
port 65 nsew default input
rlabel metal2 s 21454 27520 21510 28000 6 chany_top_in[3]
port 66 nsew default input
rlabel metal2 s 24582 0 24638 480 6 chany_top_in[4]
port 67 nsew default input
rlabel metal2 s 25962 0 26018 480 6 chany_top_in[5]
port 68 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chany_top_in[6]
port 69 nsew default input
rlabel metal3 s 0 22720 480 22840 6 chany_top_in[7]
port 70 nsew default input
rlabel metal3 s 27520 20544 28000 20664 6 chany_top_in[8]
port 71 nsew default input
rlabel metal3 s 27520 21768 28000 21888 6 chany_top_out[0]
port 72 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 27250 0 27306 480 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal3 s 27520 24488 28000 24608 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal3 s 0 25712 480 25832 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal3 s 27520 27208 28000 27328 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 1950 0 2006 480 6 data_in
port 81 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 82 nsew default input
rlabel metal3 s 0 27208 480 27328 6 left_bottom_grid_pin_12_
port 83 nsew default input
rlabel metal2 s 23386 27520 23442 28000 6 left_top_grid_pin_10_
port 84 nsew default input
rlabel metal2 s 24398 27520 24454 28000 6 right_bottom_grid_pin_12_
port 85 nsew default input
rlabel metal2 s 25410 27520 25466 28000 6 right_top_grid_pin_10_
port 86 nsew default input
rlabel metal2 s 26422 27520 26478 28000 6 top_left_grid_pin_13_
port 87 nsew default input
rlabel metal2 s 27434 27520 27490 28000 6 top_right_grid_pin_11_
port 88 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 89 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 90 nsew default input
<< end >>
