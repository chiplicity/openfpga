* NGSPICE file created from sb_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

.subckt sb_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ chanx_left_in[0] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ right_bottom_grid_pin_12_ right_top_grid_pin_11_ right_top_grid_pin_13_ right_top_grid_pin_15_
+ right_top_grid_pin_1_ right_top_grid_pin_3_ right_top_grid_pin_5_ right_top_grid_pin_7_
+ right_top_grid_pin_9_ vpwr vgnd
XFILLER_22_144 vgnd vpwr scs8hd_decap_8
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_96 vgnd vpwr scs8hd_decap_4
XFILLER_26_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_41 vgnd vpwr scs8hd_fill_1
XFILLER_13_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_155 vpwr vgnd scs8hd_fill_2
XFILLER_13_199 vgnd vpwr scs8hd_decap_6
XFILLER_27_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_147 vgnd vpwr scs8hd_decap_6
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_95 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_269 vgnd vpwr scs8hd_decap_6
XFILLER_5_173 vgnd vpwr scs8hd_decap_8
XANTENNA__124__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_228 vpwr vgnd scs8hd_fill_2
XFILLER_24_206 vgnd vpwr scs8hd_decap_8
XFILLER_32_250 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_31 vpwr vgnd scs8hd_fill_2
X_131_ _157_/A _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_12_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _188_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_64 vpwr vgnd scs8hd_fill_2
XFILLER_34_96 vgnd vpwr scs8hd_decap_3
XFILLER_34_85 vgnd vpwr scs8hd_decap_6
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
XFILLER_11_264 vgnd vpwr scs8hd_decap_12
X_114_ _114_/A address[4] _114_/C _114_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
XANTENNA__105__C _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_128 vgnd vpwr scs8hd_decap_6
XFILLER_38_117 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_7 vgnd vpwr scs8hd_decap_3
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XANTENNA__222__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_28_183 vgnd vpwr scs8hd_fill_1
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _112_/X vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_45 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_4
XFILLER_19_172 vgnd vpwr scs8hd_decap_4
XFILLER_34_186 vgnd vpwr scs8hd_fill_1
XFILLER_34_120 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_252 vpwr vgnd scs8hd_fill_2
XFILLER_0_241 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A address[6] vgnd vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_75 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_55 vgnd vpwr scs8hd_decap_4
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XANTENNA__230__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_6
XFILLER_33_207 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_5_152 vpwr vgnd scs8hd_fill_2
XFILLER_5_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _184_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _119_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_54 vgnd vpwr scs8hd_fill_1
XFILLER_15_218 vpwr vgnd scs8hd_fill_2
XFILLER_15_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _119_/A _133_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__225__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_144 vgnd vpwr scs8hd_decap_8
XANTENNA__119__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA__135__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vgnd vpwr scs8hd_decap_3
XFILLER_20_210 vpwr vgnd scs8hd_fill_2
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_3
X_113_ address[3] _114_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
XFILLER_11_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_7 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_151 vpwr vgnd scs8hd_fill_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__116__C _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_76 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_132 vpwr vgnd scs8hd_fill_2
XFILLER_31_179 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_5_ mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_143 vgnd vpwr scs8hd_decap_8
XFILLER_16_154 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B address[5] vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_157 vpwr vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_3
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_3_58 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_fill_1
XFILLER_12_190 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_45 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_6 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _139_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_22 vpwr vgnd scs8hd_fill_2
XFILLER_23_99 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_77 vgnd vpwr scs8hd_decap_12
XFILLER_34_76 vpwr vgnd scs8hd_fill_2
XANTENNA__236__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_204 vgnd vpwr scs8hd_decap_12
XFILLER_7_248 vpwr vgnd scs8hd_fill_2
XFILLER_11_200 vpwr vgnd scs8hd_fill_2
X_112_ address[5] _112_/X vgnd vpwr scs8hd_buf_1
XANTENNA__146__A _145_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_91 vpwr vgnd scs8hd_fill_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_45 vgnd vpwr scs8hd_decap_8
XFILLER_29_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_69 vpwr vgnd scs8hd_fill_2
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XFILLER_34_133 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_188 vpwr vgnd scs8hd_fill_2
XFILLER_25_155 vpwr vgnd scs8hd_fill_2
XFILLER_25_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_23 vpwr vgnd scs8hd_fill_2
XFILLER_31_99 vpwr vgnd scs8hd_fill_2
XFILLER_31_11 vgnd vpwr scs8hd_decap_12
XFILLER_0_276 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _217_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_158 vpwr vgnd scs8hd_fill_2
XFILLER_31_136 vgnd vpwr scs8hd_decap_4
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _174_/C vgnd vpwr scs8hd_diode_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_225 vgnd vpwr scs8hd_decap_12
XFILLER_39_214 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vpwr vgnd scs8hd_fill_2
XFILLER_30_191 vgnd vpwr scs8hd_decap_6
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__244__A _244_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_128 vgnd vpwr scs8hd_decap_4
XFILLER_37_10 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_261 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _203_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_78 vpwr vgnd scs8hd_fill_2
XFILLER_2_157 vgnd vpwr scs8hd_decap_12
XFILLER_2_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_223 vgnd vpwr scs8hd_decap_3
XFILLER_20_256 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_18_89 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_216 vgnd vpwr scs8hd_decap_12
X_111_ address[6] _161_/A vgnd vpwr scs8hd_buf_1
XANTENNA__162__A _112_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_175 vpwr vgnd scs8hd_fill_2
XFILLER_37_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_99 vpwr vgnd scs8hd_fill_2
XFILLER_28_186 vgnd vpwr scs8hd_fill_1
XFILLER_28_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_59 vgnd vpwr scs8hd_decap_3
XFILLER_34_167 vgnd vpwr scs8hd_decap_4
XFILLER_34_145 vpwr vgnd scs8hd_fill_2
XFILLER_34_101 vgnd vpwr scs8hd_decap_8
XANTENNA__157__A _157_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_197 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_134 vgnd vpwr scs8hd_fill_1
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_89 vgnd vpwr scs8hd_decap_4
XFILLER_31_34 vgnd vpwr scs8hd_decap_4
XFILLER_31_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_233 vgnd vpwr scs8hd_fill_1
XFILLER_16_101 vgnd vpwr scs8hd_decap_3
XFILLER_16_189 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_248 vpwr vgnd scs8hd_fill_2
XFILLER_39_237 vgnd vpwr scs8hd_decap_6
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_23 vgnd vpwr scs8hd_decap_8
XFILLER_13_115 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_137 vgnd vpwr scs8hd_decap_3
XFILLER_3_49 vgnd vpwr scs8hd_fill_1
XFILLER_8_163 vgnd vpwr scs8hd_decap_8
XFILLER_8_174 vgnd vpwr scs8hd_decap_12
XANTENNA__170__A _161_/X vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_107 vpwr vgnd scs8hd_fill_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_111 vgnd vpwr scs8hd_decap_4
XANTENNA__149__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_273 vgnd vpwr scs8hd_decap_4
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_32_254 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vpwr vgnd scs8hd_fill_2
XFILLER_23_254 vpwr vgnd scs8hd_fill_2
XFILLER_23_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_46 vpwr vgnd scs8hd_fill_2
XFILLER_2_169 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_235 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_213 vgnd vpwr scs8hd_decap_12
X_110_ _097_/A _123_/A _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_228 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_239_ _239_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_187 vpwr vgnd scs8hd_fill_2
XFILLER_29_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_198 vpwr vgnd scs8hd_fill_2
XFILLER_28_165 vgnd vpwr scs8hd_decap_12
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_3_253 vpwr vgnd scs8hd_fill_2
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_34_124 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_176 vgnd vpwr scs8hd_fill_1
XANTENNA__173__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_116 vgnd vpwr scs8hd_decap_12
XFILLER_40_105 vgnd vpwr scs8hd_decap_8
XFILLER_33_190 vpwr vgnd scs8hd_fill_2
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_256 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_113 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_205 vpwr vgnd scs8hd_fill_2
XFILLER_21_90 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_171 vgnd vpwr scs8hd_decap_3
XFILLER_22_138 vgnd vpwr scs8hd_decap_4
XFILLER_7_92 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_26_79 vpwr vgnd scs8hd_fill_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_9_109 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_208 vgnd vpwr scs8hd_decap_6
XFILLER_8_186 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_9 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_9_ mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_241 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_156 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_222 vpwr vgnd scs8hd_fill_2
XFILLER_32_200 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_211 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_14_211 vgnd vpwr scs8hd_decap_3
X_186_ _145_/A _112_/X _177_/C _102_/C _186_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__176__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_203 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_8
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_225 vgnd vpwr scs8hd_decap_4
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
X_238_ _238_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_24_90 vpwr vgnd scs8hd_fill_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
X_169_ _145_/B _174_/B vgnd vpwr scs8hd_buf_1
Xmem_bottom_track_7.LATCH_0_.latch data_in _194_/A _175_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vgnd vpwr scs8hd_decap_4
XFILLER_28_177 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_90 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__173__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_40_128 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_268 vgnd vpwr scs8hd_decap_8
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_136 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_80 vgnd vpwr scs8hd_decap_3
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_183 vpwr vgnd scs8hd_fill_2
XANTENNA__184__A _181_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_180 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__094__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_172 vgnd vpwr scs8hd_decap_4
XFILLER_8_121 vpwr vgnd scs8hd_fill_2
XFILLER_12_194 vgnd vpwr scs8hd_decap_8
XFILLER_8_198 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_275 vpwr vgnd scs8hd_fill_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_12_49 vgnd vpwr scs8hd_fill_1
XFILLER_26_253 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__089__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_4
XFILLER_17_220 vpwr vgnd scs8hd_fill_2
XANTENNA__181__B _181_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_4_61 vgnd vpwr scs8hd_fill_1
XFILLER_23_234 vpwr vgnd scs8hd_fill_2
XFILLER_3_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_138 vgnd vpwr scs8hd_decap_4
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XANTENNA__091__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_185_ _145_/A _112_/X _177_/C _099_/C _185_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XANTENNA__086__B _083_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _201_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_11_248 vpwr vgnd scs8hd_fill_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
X_168_ _161_/X _181_/B _177_/C _175_/D _168_/Y vgnd vpwr scs8hd_nor4_4
X_237_ _237_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ _102_/A address[2] _099_/C _100_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_1_95 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_29_36 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_6
XFILLER_28_123 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _202_/A _184_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_fill_1
XFILLER_19_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_156 vgnd vpwr scs8hd_decap_3
XANTENNA__173__C _145_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_25_159 vpwr vgnd scs8hd_fill_2
XFILLER_25_148 vpwr vgnd scs8hd_fill_2
XFILLER_25_126 vpwr vgnd scs8hd_fill_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_225 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_159 vgnd vpwr scs8hd_decap_3
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA__184__B _112_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_37 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_151 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_19 vgnd vpwr scs8hd_decap_12
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_144 vgnd vpwr scs8hd_decap_6
XANTENNA__170__D _174_/D vgnd vpwr scs8hd_diode_2
XANTENNA__179__B _181_/B vgnd vpwr scs8hd_diode_2
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_14 vgnd vpwr scs8hd_decap_12
XANTENNA__089__B address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_58 vgnd vpwr scs8hd_decap_3
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_265 vgnd vpwr scs8hd_decap_8
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _244_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_213 vgnd vpwr scs8hd_fill_1
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XANTENNA__181__C _145_/C vgnd vpwr scs8hd_diode_2
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XANTENNA__091__C _137_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_224 vgnd vpwr scs8hd_decap_8
XFILLER_14_235 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_184_ _181_/A _112_/X _174_/C _102_/C _184_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__176__C _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XANTENNA__086__C _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_81 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
X_236_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_167_ _102_/C _175_/D vgnd vpwr scs8hd_buf_1
X_098_ address[1] _102_/A vgnd vpwr scs8hd_inv_8
XFILLER_37_179 vpwr vgnd scs8hd_fill_2
XFILLER_37_168 vpwr vgnd scs8hd_fill_2
XFILLER_37_135 vpwr vgnd scs8hd_fill_2
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_8
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B _119_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_149 vpwr vgnd scs8hd_fill_2
XFILLER_34_127 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_168 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__173__D _175_/D vgnd vpwr scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_27 vpwr vgnd scs8hd_fill_2
XFILLER_0_237 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_3.LATCH_0_.latch data_in _190_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_193 vpwr vgnd scs8hd_fill_2
XFILLER_24_171 vgnd vpwr scs8hd_decap_8
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _204_/A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA__184__C _174_/C vgnd vpwr scs8hd_diode_2
XANTENNA__168__D _175_/D vgnd vpwr scs8hd_diode_2
XFILLER_30_163 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XFILLER_38_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _215_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_263 vgnd vpwr scs8hd_decap_12
XFILLER_29_241 vgnd vpwr scs8hd_decap_3
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_32_70 vpwr vgnd scs8hd_fill_2
XFILLER_12_163 vgnd vpwr scs8hd_decap_12
XFILLER_12_185 vgnd vpwr scs8hd_decap_3
XANTENNA__179__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_37_26 vgnd vpwr scs8hd_decap_12
XANTENNA__089__C _114_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_115 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_233 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA__181__D _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_85 vgnd vpwr scs8hd_decap_4
XFILLER_4_30 vgnd vpwr scs8hd_fill_1
XFILLER_23_258 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_129 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_203 vgnd vpwr scs8hd_decap_6
XFILLER_14_247 vgnd vpwr scs8hd_decap_8
XFILLER_14_258 vgnd vpwr scs8hd_decap_12
X_183_ _181_/A _112_/X _174_/C _099_/C _183_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
XFILLER_13_94 vpwr vgnd scs8hd_fill_2
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_38_80 vgnd vpwr scs8hd_fill_1
XANTENNA__176__D _174_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_262 vgnd vpwr scs8hd_decap_12
XFILLER_20_206 vpwr vgnd scs8hd_fill_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_4
X_235_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ _161_/X _181_/B _177_/C _174_/D _166_/Y vgnd vpwr scs8hd_nor4_4
X_097_ _097_/A _119_/A _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_147 vpwr vgnd scs8hd_fill_2
XFILLER_34_6 vgnd vpwr scs8hd_decap_12
XFILLER_1_31 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_86 vgnd vpwr scs8hd_fill_1
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
X_149_ _157_/A _150_/B _149_/Y vgnd vpwr scs8hd_nor2_4
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_194 vpwr vgnd scs8hd_fill_2
XFILLER_33_161 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_205 vgnd vpwr scs8hd_fill_1
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _198_/A _180_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_131 vpwr vgnd scs8hd_fill_2
XFILLER_22_109 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XANTENNA__184__D _102_/C vgnd vpwr scs8hd_diode_2
XFILLER_15_172 vpwr vgnd scs8hd_fill_2
XFILLER_7_30 vpwr vgnd scs8hd_fill_2
XFILLER_38_242 vgnd vpwr scs8hd_decap_12
XFILLER_26_17 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_275 vpwr vgnd scs8hd_fill_2
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_16_61 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vgnd vpwr scs8hd_decap_4
XFILLER_12_175 vgnd vpwr scs8hd_fill_1
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA__179__D _174_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_38 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XFILLER_32_259 vgnd vpwr scs8hd_decap_12
XFILLER_32_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_20 vpwr vgnd scs8hd_fill_2
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XFILLER_4_53 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
X_182_ _181_/A _181_/B _145_/C _102_/C _182_/Y vgnd vpwr scs8hd_nor4_4
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _100_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_274 vgnd vpwr scs8hd_decap_3
XFILLER_20_218 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_229 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_7 vgnd vpwr scs8hd_decap_12
X_165_ _099_/C _174_/D vgnd vpwr scs8hd_buf_1
XFILLER_6_211 vgnd vpwr scs8hd_decap_3
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_234_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_40_71 vgnd vpwr scs8hd_decap_12
X_096_ _095_/X _119_/A vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_43 vgnd vpwr scs8hd_decap_12
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _199_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_148_ _119_/A _150_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XFILLER_18_170 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_3
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _156_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_73 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_187 vpwr vgnd scs8hd_fill_2
XFILLER_30_143 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vpwr vgnd scs8hd_fill_2
XFILLER_38_254 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_176 vgnd vpwr scs8hd_fill_1
XFILLER_29_221 vgnd vpwr scs8hd_decap_12
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_32_83 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _185_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_7_ mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_202 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _203_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_224 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_238 vgnd vpwr scs8hd_decap_12
XFILLER_32_205 vpwr vgnd scs8hd_fill_2
XFILLER_27_50 vgnd vpwr scs8hd_decap_4
XFILLER_17_202 vgnd vpwr scs8hd_decap_3
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_238 vgnd vpwr scs8hd_decap_4
XFILLER_23_19 vgnd vpwr scs8hd_fill_1
XFILLER_13_52 vgnd vpwr scs8hd_decap_3
X_181_ _181_/A _181_/B _145_/C _099_/C _181_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_153 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_34_18 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_233_ _233_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr
+ scs8hd_diode_2
X_164_ _163_/X _177_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_095_ address[1] _083_/Y _102_/C _095_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_83 vgnd vpwr scs8hd_decap_8
XFILLER_1_55 vgnd vpwr scs8hd_decap_6
XANTENNA__111__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
X_147_ _118_/A _150_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _105_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XFILLER_18_193 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_4
XFILLER_0_229 vgnd vpwr scs8hd_decap_4
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_266 vgnd vpwr scs8hd_decap_8
XFILLER_38_200 vgnd vpwr scs8hd_decap_12
XFILLER_21_188 vgnd vpwr scs8hd_decap_3
XFILLER_29_233 vgnd vpwr scs8hd_decap_8
XFILLER_32_51 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_104 vpwr vgnd scs8hd_fill_2
XFILLER_16_96 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_214 vgnd vpwr scs8hd_decap_12
XFILLER_7_170 vgnd vpwr scs8hd_fill_1
XFILLER_7_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _202_/A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_5_107 vpwr vgnd scs8hd_fill_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_77 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_6
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_228 vgnd vpwr scs8hd_decap_4
XFILLER_23_206 vgnd vpwr scs8hd_decap_3
XFILLER_22_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_180_ _181_/A _181_/B _137_/C _175_/D _180_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_232_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_163_ _114_/A _124_/Y _114_/C _163_/X vgnd vpwr scs8hd_or3_4
X_094_ address[0] _102_/C vgnd vpwr scs8hd_buf_1
XFILLER_37_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_10_21 vgnd vpwr scs8hd_decap_4
XFILLER_10_32 vgnd vpwr scs8hd_decap_4
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_34_109 vpwr vgnd scs8hd_fill_2
XFILLER_19_85 vgnd vpwr scs8hd_decap_3
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_146_ _145_/X _150_/B vgnd vpwr scs8hd_buf_1
XFILLER_33_175 vpwr vgnd scs8hd_fill_2
XFILLER_33_153 vpwr vgnd scs8hd_fill_2
XFILLER_33_142 vpwr vgnd scs8hd_fill_2
XFILLER_18_150 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_24_142 vgnd vpwr scs8hd_decap_8
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_86 vpwr vgnd scs8hd_fill_2
XFILLER_30_101 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_142 vgnd vpwr scs8hd_decap_4
XFILLER_15_153 vpwr vgnd scs8hd_fill_2
XFILLER_30_167 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _116_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_55 vpwr vgnd scs8hd_fill_2
XFILLER_7_11 vgnd vpwr scs8hd_decap_3
XFILLER_7_88 vgnd vpwr scs8hd_decap_4
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _118_/A _133_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _195_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_134 vpwr vgnd scs8hd_fill_2
XFILLER_21_156 vgnd vpwr scs8hd_decap_3
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_7.LATCH_1_.latch data_in _193_/A _174_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_53 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_138 vgnd vpwr scs8hd_decap_4
XFILLER_12_145 vgnd vpwr scs8hd_decap_8
XFILLER_35_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__220__A _220_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_237 vgnd vpwr scs8hd_decap_6
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_32_218 vpwr vgnd scs8hd_fill_2
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XFILLER_27_85 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_163 vgnd vpwr scs8hd_decap_12
XFILLER_4_89 vgnd vpwr scs8hd_fill_1
XFILLER_4_12 vgnd vpwr scs8hd_decap_6
XANTENNA__130__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_87 vpwr vgnd scs8hd_fill_2
XFILLER_13_98 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_166 vgnd vpwr scs8hd_decap_12
XFILLER_38_84 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_231_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_24_64 vpwr vgnd scs8hd_fill_2
X_162_ _112_/X _181_/B vgnd vpwr scs8hd_buf_1
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _118_/A _097_/A _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_4
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ _145_/A _145_/B _145_/C _145_/X vgnd vpwr scs8hd_or3_4
XANTENNA__122__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _205_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XFILLER_24_121 vgnd vpwr scs8hd_decap_8
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_10 vpwr vgnd scs8hd_fill_2
XANTENNA__223__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_135 vgnd vpwr scs8hd_decap_4
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _122_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _133_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _197_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_21_113 vgnd vpwr scs8hd_decap_6
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_29_213 vpwr vgnd scs8hd_fill_2
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XFILLER_35_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_15.LATCH_1_.latch data_in _201_/A _183_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_31 vgnd vpwr scs8hd_decap_4
XFILLER_27_20 vpwr vgnd scs8hd_fill_2
XFILLER_17_216 vpwr vgnd scs8hd_fill_2
XFILLER_17_249 vgnd vpwr scs8hd_decap_12
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_175 vgnd vpwr scs8hd_decap_12
XFILLER_4_24 vgnd vpwr scs8hd_decap_6
XANTENNA__114__C _114_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XFILLER_31_241 vgnd vpwr scs8hd_decap_3
XFILLER_22_252 vgnd vpwr scs8hd_decap_12
XFILLER_22_241 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _201_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_22 vgnd vpwr scs8hd_decap_3
XFILLER_38_30 vgnd vpwr scs8hd_fill_1
XANTENNA__231__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_156 vpwr vgnd scs8hd_fill_2
XFILLER_1_178 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_8
XANTENNA__141__A _157_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_193 vgnd vpwr scs8hd_decap_12
XFILLER_24_87 vgnd vpwr scs8hd_fill_1
XFILLER_24_43 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
X_161_ _161_/A _161_/X vgnd vpwr scs8hd_buf_1
X_230_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XANTENNA__226__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_40_64 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_092_ _091_/X _097_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_119 vgnd vpwr scs8hd_fill_1
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_54 vgnd vpwr scs8hd_decap_4
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_174 vgnd vpwr scs8hd_decap_3
XFILLER_27_163 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _123_/A _139_/B _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_174 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_111 vpwr vgnd scs8hd_fill_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_90 vpwr vgnd scs8hd_fill_2
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_188 vgnd vpwr scs8hd_decap_3
XFILLER_21_22 vpwr vgnd scs8hd_fill_2
XFILLER_21_77 vgnd vpwr scs8hd_fill_1
XFILLER_30_147 vgnd vpwr scs8hd_decap_4
XFILLER_30_114 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_188 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
X_127_ address[6] address[5] _174_/C _128_/A vgnd vpwr scs8hd_or3_4
XFILLER_16_3 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _246_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_6
XANTENNA__234__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vgnd vpwr scs8hd_decap_3
XFILLER_7_162 vgnd vpwr scs8hd_decap_8
XFILLER_7_173 vgnd vpwr scs8hd_decap_8
XFILLER_26_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_209 vgnd vpwr scs8hd_decap_4
XFILLER_27_65 vpwr vgnd scs8hd_fill_2
XFILLER_27_54 vgnd vpwr scs8hd_fill_1
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_187 vgnd vpwr scs8hd_decap_12
XFILLER_4_132 vgnd vpwr scs8hd_decap_4
Xmem_bottom_track_3.LATCH_1_.latch data_in _189_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_264 vgnd vpwr scs8hd_decap_8
XFILLER_1_113 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _200_/A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_220 vpwr vgnd scs8hd_fill_2
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XANTENNA__125__C _114_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_253 vpwr vgnd scs8hd_fill_2
XANTENNA__141__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_90 vpwr vgnd scs8hd_fill_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_160_ _123_/A _159_/B _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_091_ address[6] address[5] _137_/C _091_/X vgnd vpwr scs8hd_or3_4
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_175 vgnd vpwr scs8hd_decap_12
XFILLER_36_164 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_27_142 vgnd vpwr scs8hd_decap_4
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _122_/A _139_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _204_/Y mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_142 vgnd vpwr scs8hd_decap_8
XANTENNA__147__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_45 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_47 vpwr vgnd scs8hd_fill_2
X_126_ _125_/X _174_/C vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_29_259 vpwr vgnd scs8hd_fill_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_8_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _123_/A vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _123_/A vgnd vpwr scs8hd_buf_1
XFILLER_26_229 vgnd vpwr scs8hd_decap_3
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XFILLER_25_240 vgnd vpwr scs8hd_decap_4
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _193_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__245__A _245_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_199 vgnd vpwr scs8hd_decap_12
XFILLER_4_122 vgnd vpwr scs8hd_decap_3
XANTENNA__155__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_11.LATCH_1_.latch data_in _197_/A _179_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XFILLER_1_103 vpwr vgnd scs8hd_fill_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_6
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_203 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_39_184 vgnd vpwr scs8hd_fill_1
XFILLER_24_23 vgnd vpwr scs8hd_decap_6
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
X_090_ _089_/X _137_/C vgnd vpwr scs8hd_buf_1
XFILLER_10_202 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_8
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__152__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_12 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_132 vgnd vpwr scs8hd_decap_4
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
X_142_ _121_/A _139_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_179 vpwr vgnd scs8hd_fill_2
XFILLER_33_157 vpwr vgnd scs8hd_fill_2
XFILLER_33_146 vpwr vgnd scs8hd_fill_2
XFILLER_33_113 vpwr vgnd scs8hd_fill_2
XANTENNA__147__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_132 vgnd vpwr scs8hd_fill_1
XFILLER_18_154 vgnd vpwr scs8hd_decap_3
XANTENNA__163__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_70 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_113 vgnd vpwr scs8hd_decap_3
XFILLER_15_157 vpwr vgnd scs8hd_fill_2
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
X_125_ address[3] _124_/Y _114_/C _125_/X vgnd vpwr scs8hd_or3_4
XANTENNA__158__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_105 vpwr vgnd scs8hd_fill_2
XFILLER_21_138 vpwr vgnd scs8hd_fill_2
XFILLER_16_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_260 vgnd vpwr scs8hd_decap_12
XFILLER_11_193 vgnd vpwr scs8hd_decap_4
X_108_ address[1] address[2] address[0] _109_/A vgnd vpwr scs8hd_or3_4
XANTENNA__160__B _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _155_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_27_89 vpwr vgnd scs8hd_fill_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__155__B _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _206_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_215 vgnd vpwr scs8hd_decap_12
XFILLER_0_170 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _161_/X vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _207_/HI _199_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _196_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_10_59 vgnd vpwr scs8hd_decap_4
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_27_188 vgnd vpwr scs8hd_fill_1
XFILLER_27_100 vpwr vgnd scs8hd_fill_2
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
X_141_ _157_/A _139_/B _141_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_166 vpwr vgnd scs8hd_fill_2
XANTENNA__163__B _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_2_82 vgnd vpwr scs8hd_decap_8
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_14 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_139 vgnd vpwr scs8hd_fill_1
XFILLER_23_191 vpwr vgnd scs8hd_fill_2
X_124_ address[4] _124_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_16 vgnd vpwr scs8hd_decap_3
XFILLER_23_7 vgnd vpwr scs8hd_decap_12
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XANTENNA__158__B _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _161_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vgnd vpwr scs8hd_decap_6
XANTENNA__084__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_28_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _155_/Y vgnd vpwr scs8hd_diode_2
X_107_ _097_/A _122_/A _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_3
XANTENNA__169__A _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vgnd vpwr scs8hd_decap_4
XFILLER_27_35 vgnd vpwr scs8hd_fill_1
XFILLER_27_24 vpwr vgnd scs8hd_fill_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XFILLER_31_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__171__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_48 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_234 vgnd vpwr scs8hd_decap_8
XFILLER_13_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_182 vgnd vpwr scs8hd_decap_4
XANTENNA__166__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XANTENNA__182__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_164 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_47 vgnd vpwr scs8hd_decap_6
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_80 vpwr vgnd scs8hd_fill_2
XFILLER_36_145 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _198_/A mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__177__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_38 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_19_58 vgnd vpwr scs8hd_fill_1
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_140_ _119_/A _139_/B _140_/Y vgnd vpwr scs8hd_nor2_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_189 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__163__C _114_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_115 vgnd vpwr scs8hd_decap_3
XFILLER_21_26 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_181 vpwr vgnd scs8hd_fill_2
X_123_ _123_/A _121_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_70 vpwr vgnd scs8hd_fill_2
XFILLER_16_7 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__174__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _202_/Y mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_107 vgnd vpwr scs8hd_decap_6
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_58 vgnd vpwr scs8hd_decap_12
XFILLER_32_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
X_106_ _105_/X _122_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_188 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_82 vpwr vgnd scs8hd_fill_2
XFILLER_27_69 vgnd vpwr scs8hd_decap_3
XFILLER_25_232 vpwr vgnd scs8hd_fill_2
XFILLER_25_221 vpwr vgnd scs8hd_fill_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_91 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_180 vgnd vpwr scs8hd_decap_3
XANTENNA__171__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_224 vgnd vpwr scs8hd_decap_3
XFILLER_22_202 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_224 vgnd vpwr scs8hd_decap_8
XFILLER_9_239 vgnd vpwr scs8hd_decap_4
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_3_ mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _191_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__166__C _177_/C vgnd vpwr scs8hd_diode_2
XANTENNA__182__B _181_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_94 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XFILLER_1_19 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA__177__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_179 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_80 vgnd vpwr scs8hd_decap_6
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_138 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _195_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_182 vgnd vpwr scs8hd_fill_1
XFILLER_21_49 vgnd vpwr scs8hd_fill_1
XANTENNA__098__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
XFILLER_15_149 vpwr vgnd scs8hd_fill_2
X_122_ _122_/A _121_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__C _174_/C vgnd vpwr scs8hd_diode_2
XFILLER_21_119 vgnd vpwr scs8hd_fill_1
XFILLER_37_241 vgnd vpwr scs8hd_decap_3
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_16_49 vpwr vgnd scs8hd_fill_2
XFILLER_20_141 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_20_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_70 vgnd vpwr scs8hd_decap_8
XFILLER_7_112 vgnd vpwr scs8hd_decap_4
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_156 vgnd vpwr scs8hd_decap_3
XFILLER_11_152 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vpwr vgnd scs8hd_fill_2
X_105_ address[1] address[2] _105_/C _105_/X vgnd vpwr scs8hd_or3_4
XFILLER_22_81 vgnd vpwr scs8hd_decap_8
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XFILLER_19_263 vgnd vpwr scs8hd_decap_12
XFILLER_21_6 vpwr vgnd scs8hd_fill_2
XANTENNA__185__B _112_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XANTENNA__095__B _083_/Y vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_91 vpwr vgnd scs8hd_fill_2
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _175_/D vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_151 vgnd vpwr scs8hd_decap_4
XFILLER_0_162 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__D _174_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_73 vpwr vgnd scs8hd_fill_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_4
XANTENNA__182__C _145_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_3
XANTENNA__177__C _177_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_33_117 vgnd vpwr scs8hd_decap_4
XFILLER_18_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_125 vgnd vpwr scs8hd_decap_4
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _206_/HI _197_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_106 vgnd vpwr scs8hd_decap_3
XFILLER_32_194 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _194_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_121_ _121_/A _121_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_172 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_14_161 vgnd vpwr scs8hd_decap_3
XFILLER_21_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__D _174_/D vgnd vpwr scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_197 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_11_197 vgnd vpwr scs8hd_fill_1
X_104_ _097_/A _121_/A _104_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_242 vpwr vgnd scs8hd_fill_2
XFILLER_19_253 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XANTENNA__185__C _177_/C vgnd vpwr scs8hd_diode_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_27_38 vgnd vpwr scs8hd_fill_1
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XANTENNA__095__C _102_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_70 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _216_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_160 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_18 vpwr vgnd scs8hd_fill_2
XFILLER_21_270 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _207_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_270 vgnd vpwr scs8hd_decap_4
XANTENNA__182__D _102_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_189 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_82 vpwr vgnd scs8hd_fill_2
XANTENNA__177__D _175_/D vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_159 vpwr vgnd scs8hd_fill_2
XFILLER_27_104 vgnd vpwr scs8hd_fill_1
XFILLER_35_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_26_181 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_17_181 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _157_/A _121_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_62 vgnd vpwr scs8hd_fill_1
XFILLER_11_95 vgnd vpwr scs8hd_decap_3
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_121 vpwr vgnd scs8hd_fill_2
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vgnd vpwr scs8hd_decap_4
X_103_ _102_/X _121_/A vgnd vpwr scs8hd_buf_1
XANTENNA__185__D _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_8_74 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_128 vpwr vgnd scs8hd_fill_2
XFILLER_4_117 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _200_/Y mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_224 vgnd vpwr scs8hd_decap_8
XFILLER_16_235 vgnd vpwr scs8hd_decap_12
XFILLER_17_83 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vgnd vpwr scs8hd_decap_8
XFILLER_30_260 vgnd vpwr scs8hd_decap_12
XFILLER_1_109 vpwr vgnd scs8hd_fill_2
XFILLER_13_216 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vgnd vpwr scs8hd_decap_6
XFILLER_5_31 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_168 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_39_81 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _189_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_50 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_6 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_32_174 vgnd vpwr scs8hd_decap_8
XFILLER_32_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_130 vgnd vpwr scs8hd_decap_4
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
XFILLER_14_185 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_179_ _181_/A _181_/B _137_/C _174_/D _179_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _193_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_100 vgnd vpwr scs8hd_fill_1
X_102_ _102_/A address[2] _102_/C _102_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XFILLER_8_53 vpwr vgnd scs8hd_fill_2
XFILLER_8_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_25_236 vpwr vgnd scs8hd_fill_2
XFILLER_31_217 vgnd vpwr scs8hd_decap_3
XFILLER_16_247 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_50 vgnd vpwr scs8hd_decap_8
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_151 vgnd vpwr scs8hd_decap_3
XANTENNA__104__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_6
XFILLER_30_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_8_210 vgnd vpwr scs8hd_decap_4
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _196_/A _177_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _190_/Y mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_19 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_40 vpwr vgnd scs8hd_fill_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_93 vgnd vpwr scs8hd_decap_8
XFILLER_36_128 vgnd vpwr scs8hd_decap_6
XFILLER_36_117 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_180 vgnd vpwr scs8hd_fill_1
XANTENNA__101__B _157_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XFILLER_2_205 vgnd vpwr scs8hd_decap_8
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_106 vgnd vpwr scs8hd_decap_6
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_32_131 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_131 vpwr vgnd scs8hd_fill_2
XFILLER_23_120 vpwr vgnd scs8hd_fill_2
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _145_/A _181_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_145 vgnd vpwr scs8hd_decap_8
XFILLER_20_167 vpwr vgnd scs8hd_fill_2
XFILLER_20_178 vgnd vpwr scs8hd_decap_6
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_fill_1
XFILLER_11_156 vpwr vgnd scs8hd_fill_2
XFILLER_11_178 vgnd vpwr scs8hd_decap_3
X_101_ _097_/A _157_/A _101_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _192_/A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_201 vgnd vpwr scs8hd_fill_1
XFILLER_19_234 vgnd vpwr scs8hd_decap_8
XFILLER_19_245 vpwr vgnd scs8hd_fill_2
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_229 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_8
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _157_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_22_229 vgnd vpwr scs8hd_decap_3
XFILLER_38_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _186_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 right_top_grid_pin_1_ mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A right_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XFILLER_28_51 vgnd vpwr scs8hd_decap_4
XFILLER_0_166 vpwr vgnd scs8hd_fill_2
XFILLER_0_199 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__115__A _114_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vpwr vgnd scs8hd_fill_2
XFILLER_39_115 vgnd vpwr scs8hd_decap_6
XFILLER_5_77 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _196_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _204_/A _186_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_30_96 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XFILLER_26_173 vgnd vpwr scs8hd_decap_8
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XFILLER_26_195 vpwr vgnd scs8hd_fill_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_32_143 vpwr vgnd scs8hd_fill_2
XFILLER_17_173 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_3
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _183_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_246_ _246_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_177_ _161_/A _145_/B _177_/C _175_/D _177_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__107__B _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_191 vgnd vpwr scs8hd_decap_12
XFILLER_28_202 vpwr vgnd scs8hd_fill_2
XFILLER_28_224 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vpwr vgnd scs8hd_fill_2
X_100_ _100_/A _157_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_97 vgnd vpwr scs8hd_decap_3
XFILLER_19_213 vgnd vpwr scs8hd_decap_6
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_229_ _229_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_20 vgnd vpwr scs8hd_decap_4
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__221__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_156 vgnd vpwr scs8hd_decap_6
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_34 vgnd vpwr scs8hd_fill_1
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _198_/Y mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__131__A _157_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 right_top_grid_pin_11_ mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_76 vpwr vgnd scs8hd_fill_2
XFILLER_30_86 vgnd vpwr scs8hd_decap_6
XFILLER_39_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__A _125_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_270 vgnd vpwr scs8hd_decap_4
XFILLER_35_174 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_5.LATCH_0_.latch data_in _192_/A _173_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_6
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XFILLER_25_97 vpwr vgnd scs8hd_fill_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_177 vpwr vgnd scs8hd_fill_2
XFILLER_23_155 vpwr vgnd scs8hd_fill_2
XFILLER_23_144 vpwr vgnd scs8hd_fill_2
XFILLER_2_6 vgnd vpwr scs8hd_decap_12
XFILLER_11_66 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _187_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_122 vpwr vgnd scs8hd_fill_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_14_166 vpwr vgnd scs8hd_fill_2
XFILLER_14_177 vgnd vpwr scs8hd_decap_8
X_245_ _245_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_14_199 vpwr vgnd scs8hd_fill_2
X_176_ _161_/A _145_/B _177_/C _174_/D _176_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__123__B _121_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_37_203 vgnd vpwr scs8hd_decap_12
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_181 vpwr vgnd scs8hd_fill_2
XFILLER_28_236 vgnd vpwr scs8hd_decap_12
XFILLER_11_114 vgnd vpwr scs8hd_fill_1
XFILLER_22_43 vgnd vpwr scs8hd_decap_12
XFILLER_22_32 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_169 vgnd vpwr scs8hd_decap_3
XANTENNA__224__A _224_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XANTENNA__118__B _121_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
X_159_ _122_/A _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
X_228_ _228_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_8_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__134__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_217 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _147_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _191_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_113 vpwr vgnd scs8hd_fill_2
XFILLER_28_64 vgnd vpwr scs8hd_decap_4
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_55 vpwr vgnd scs8hd_fill_2
XFILLER_14_88 vgnd vpwr scs8hd_decap_4
XFILLER_30_65 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XANTENNA__232__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _121_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_153 vpwr vgnd scs8hd_fill_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XANTENNA__227__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_120 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_54 vgnd vpwr scs8hd_decap_6
XPHY_43 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _205_/HI _188_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmem_bottom_track_13.LATCH_0_.latch data_in _200_/A _182_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_112 vgnd vpwr scs8hd_decap_4
XANTENNA__137__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _219_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
X_244_ _244_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_14_134 vgnd vpwr scs8hd_fill_1
X_175_ _161_/A _174_/B _174_/C _175_/D _175_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_20_104 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_248 vgnd vpwr scs8hd_decap_12
XFILLER_3_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_108 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
X_158_ _121_/A _159_/B _158_/Y vgnd vpwr scs8hd_nor2_4
X_089_ address[3] address[4] _114_/C _089_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_163 vgnd vpwr scs8hd_decap_12
XANTENNA__134__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _190_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_0_91 vpwr vgnd scs8hd_fill_2
XFILLER_21_254 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_4
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_107 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vpwr vgnd scs8hd_fill_2
XFILLER_29_195 vpwr vgnd scs8hd_fill_2
XFILLER_29_151 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _218_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_35_198 vpwr vgnd scs8hd_fill_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _194_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vpwr vgnd scs8hd_fill_2
XFILLER_25_33 vpwr vgnd scs8hd_fill_2
XFILLER_25_11 vgnd vpwr scs8hd_decap_8
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XFILLER_17_154 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XFILLER_32_168 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_198 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _188_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_243_ _243_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_157 vpwr vgnd scs8hd_fill_2
X_174_ _161_/A _174_/B _174_/C _174_/D _174_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__148__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XFILLER_22_12 vgnd vpwr scs8hd_decap_8
XFILLER_22_89 vgnd vpwr scs8hd_fill_1
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XFILLER_34_208 vgnd vpwr scs8hd_decap_6
XFILLER_19_249 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_157_ _157_/A _159_/B _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_131 vpwr vgnd scs8hd_fill_2
XFILLER_6_142 vpwr vgnd scs8hd_fill_2
XFILLER_8_36 vpwr vgnd scs8hd_fill_2
X_226_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
X_088_ enable _114_/C vgnd vpwr scs8hd_inv_8
XFILLER_6_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_241 vgnd vpwr scs8hd_decap_12
XFILLER_17_56 vgnd vpwr scs8hd_decap_3
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vpwr vgnd scs8hd_fill_2
XFILLER_3_101 vgnd vpwr scs8hd_decap_8
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_266 vpwr vgnd scs8hd_fill_2
XFILLER_9_90 vpwr vgnd scs8hd_fill_2
XFILLER_0_137 vgnd vpwr scs8hd_decap_6
XANTENNA__246__A _246_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XFILLER_30_23 vgnd vpwr scs8hd_decap_8
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_30_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_4
XFILLER_26_100 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vpwr vgnd scs8hd_fill_2
XFILLER_25_67 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_32_147 vgnd vpwr scs8hd_decap_6
XFILLER_32_125 vgnd vpwr scs8hd_decap_6
XFILLER_17_177 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _137_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _145_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_15_ mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_114 vgnd vpwr scs8hd_decap_4
XFILLER_23_103 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
X_242_ _242_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_173_ _161_/X _174_/B _145_/C _175_/D _173_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_217 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_173 vpwr vgnd scs8hd_fill_2
XFILLER_13_180 vgnd vpwr scs8hd_fill_1
XFILLER_28_206 vgnd vpwr scs8hd_decap_4
XFILLER_22_57 vpwr vgnd scs8hd_fill_2
XFILLER_11_117 vgnd vpwr scs8hd_decap_3
XFILLER_11_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
X_225_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_156_ _119_/A _159_/B _156_/Y vgnd vpwr scs8hd_nor2_4
X_087_ _087_/A _118_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_187 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_209 vgnd vpwr scs8hd_decap_6
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_34 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_253 vpwr vgnd scs8hd_fill_2
XFILLER_17_24 vgnd vpwr scs8hd_fill_1
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
XFILLER_33_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__C _145_/C vgnd vpwr scs8hd_diode_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
X_139_ _118_/A _139_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_71 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_223 vpwr vgnd scs8hd_fill_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_234 vgnd vpwr scs8hd_decap_12
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_4
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XFILLER_10_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__156__B _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _161_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _189_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _245_/A vgnd vpwr scs8hd_inv_1
XFILLER_30_57 vgnd vpwr scs8hd_decap_6
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_77 vpwr vgnd scs8hd_fill_2
XFILLER_39_66 vgnd vpwr scs8hd_fill_1
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XFILLER_35_134 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _102_/C vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_17_112 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _174_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_159 vpwr vgnd scs8hd_fill_2
XFILLER_23_148 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _195_/A _176_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_126 vpwr vgnd scs8hd_fill_2
XFILLER_14_148 vgnd vpwr scs8hd_decap_4
X_241_ _241_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
X_172_ _161_/X _174_/B _145_/C _174_/D _172_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_229 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_129 vgnd vpwr scs8hd_fill_1
XANTENNA__180__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A _089_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_8_49 vpwr vgnd scs8hd_fill_2
X_224_ _224_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
X_155_ _118_/A _159_/B _155_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_199 vgnd vpwr scs8hd_decap_12
X_086_ address[1] _083_/Y _099_/C _087_/A vgnd vpwr scs8hd_or3_4
XFILLER_12_80 vpwr vgnd scs8hd_fill_2
XFILLER_33_7 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _161_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _105_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_243 vgnd vpwr scs8hd_fill_1
XFILLER_30_224 vgnd vpwr scs8hd_decap_12
X_207_ _207_/HI _207_/LO vgnd vpwr scs8hd_conb_1
X_138_ _137_/X _139_/B vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_83 vgnd vpwr scs8hd_decap_8
XFILLER_0_94 vgnd vpwr scs8hd_decap_12
XFILLER_21_202 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_3
XFILLER_0_117 vgnd vpwr scs8hd_decap_6
XFILLER_28_68 vgnd vpwr scs8hd_fill_1
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_246 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_176 vgnd vpwr scs8hd_decap_12
XFILLER_38_165 vgnd vpwr scs8hd_decap_8
XFILLER_38_154 vpwr vgnd scs8hd_fill_2
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _188_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_34 vgnd vpwr scs8hd_decap_12
XFILLER_29_132 vgnd vpwr scs8hd_decap_4
XFILLER_29_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_179 vpwr vgnd scs8hd_fill_2
XFILLER_35_157 vpwr vgnd scs8hd_fill_2
XANTENNA__183__A _181_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_8
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_127 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_171 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A enable vgnd vpwr scs8hd_diode_2
X_240_ _240_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_105 vpwr vgnd scs8hd_fill_2
X_171_ _161_/X _174_/B _137_/C _175_/D _171_/Y vgnd vpwr scs8hd_nor4_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _192_/Y mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in _203_/A _185_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__180__B _181_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XFILLER_3_72 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_252 vgnd vpwr scs8hd_decap_12
X_223_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
X_154_ _153_/X _159_/B vgnd vpwr scs8hd_buf_1
XFILLER_10_163 vpwr vgnd scs8hd_fill_2
X_085_ _105_/C _099_/C vgnd vpwr scs8hd_buf_1
XFILLER_33_211 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__175__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_222 vpwr vgnd scs8hd_fill_2
XFILLER_15_233 vpwr vgnd scs8hd_fill_2
XFILLER_30_236 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_206_ _206_/HI _206_/LO vgnd vpwr scs8hd_conb_1
X_137_ _145_/A _145_/B _137_/C _137_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_181 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_21_258 vgnd vpwr scs8hd_decap_4
XANTENNA__186__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _220_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_47 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _095_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_258 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_240 vgnd vpwr scs8hd_decap_4
XANTENNA__172__C _145_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_188 vgnd vpwr scs8hd_decap_12
XFILLER_38_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XFILLER_14_49 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_4
XFILLER_39_46 vgnd vpwr scs8hd_decap_12
XFILLER_29_155 vpwr vgnd scs8hd_fill_2
XFILLER_29_199 vgnd vpwr scs8hd_decap_3
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_20_70 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _224_/A vgnd vpwr scs8hd_inv_1
XANTENNA__183__B _112_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_103 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_169 vpwr vgnd scs8hd_fill_2
XFILLER_26_147 vgnd vpwr scs8hd_fill_1
XFILLER_26_125 vgnd vpwr scs8hd_decap_3
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__093__B _097_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_147 vpwr vgnd scs8hd_fill_2
XFILLER_17_158 vpwr vgnd scs8hd_fill_2
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_28 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_194 vpwr vgnd scs8hd_fill_2
XFILLER_22_161 vpwr vgnd scs8hd_fill_2
X_170_ _161_/X _174_/B _137_/C _174_/D _170_/Y vgnd vpwr scs8hd_nor4_4
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_9_143 vpwr vgnd scs8hd_fill_2
XFILLER_9_187 vpwr vgnd scs8hd_fill_2
XFILLER_13_172 vpwr vgnd scs8hd_fill_2
XANTENNA__180__C _137_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_84 vgnd vpwr scs8hd_decap_3
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_264 vgnd vpwr scs8hd_decap_12
X_222_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
Xmem_bottom_track_5.LATCH_1_.latch data_in _191_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
XFILLER_6_135 vgnd vpwr scs8hd_decap_4
XFILLER_10_120 vpwr vgnd scs8hd_fill_2
XFILLER_10_175 vgnd vpwr scs8hd_decap_8
XFILLER_10_186 vpwr vgnd scs8hd_fill_2
X_153_ _145_/A _145_/B _174_/C _153_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_146 vgnd vpwr scs8hd_decap_6
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
X_084_ address[0] _105_/C vgnd vpwr scs8hd_inv_8
XFILLER_19_7 vgnd vpwr scs8hd_decap_3
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
XANTENNA__175__C _174_/C vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_16 vpwr vgnd scs8hd_fill_2
XFILLER_17_27 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_138 vpwr vgnd scs8hd_fill_2
XFILLER_3_127 vgnd vpwr scs8hd_decap_4
XFILLER_15_201 vpwr vgnd scs8hd_fill_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_30_248 vgnd vpwr scs8hd_decap_12
X_205_ _205_/HI _205_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_136_ address[5] _145_/B vgnd vpwr scs8hd_inv_8
XFILLER_2_193 vgnd vpwr scs8hd_decap_12
XANTENNA__186__B _112_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
X_119_ _119_/A _121_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_252 vgnd vpwr scs8hd_decap_3
XANTENNA__172__D _174_/D vgnd vpwr scs8hd_diode_2
XFILLER_38_134 vgnd vpwr scs8hd_fill_1
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A right_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_69 vgnd vpwr scs8hd_decap_4
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_112 vgnd vpwr scs8hd_decap_4
XFILLER_4_211 vgnd vpwr scs8hd_decap_3
XFILLER_29_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__183__C _174_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XFILLER_26_137 vpwr vgnd scs8hd_fill_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _187_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_17_126 vpwr vgnd scs8hd_fill_2
XFILLER_40_140 vgnd vpwr scs8hd_decap_12
XFILLER_25_192 vpwr vgnd scs8hd_fill_2
XFILLER_31_140 vgnd vpwr scs8hd_fill_1
XFILLER_31_195 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_166 vpwr vgnd scs8hd_fill_2
XFILLER_9_177 vpwr vgnd scs8hd_fill_2
XFILLER_13_184 vpwr vgnd scs8hd_fill_2
XFILLER_3_52 vgnd vpwr scs8hd_decap_6
XANTENNA__180__D _175_/D vgnd vpwr scs8hd_diode_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_276 vgnd vpwr scs8hd_fill_1
X_152_ _123_/A _150_/B _152_/Y vgnd vpwr scs8hd_nor2_4
X_221_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_114 vgnd vpwr scs8hd_decap_6
XFILLER_10_143 vpwr vgnd scs8hd_fill_2
XFILLER_12_61 vpwr vgnd scs8hd_fill_2
X_083_ address[2] _083_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A right_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_80 vgnd vpwr scs8hd_fill_1
XFILLER_26_9 vgnd vpwr scs8hd_decap_8
XFILLER_18_254 vgnd vpwr scs8hd_fill_1
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XFILLER_33_224 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _175_/D vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_13.LATCH_1_.latch data_in _199_/A _181_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_224 vpwr vgnd scs8hd_fill_2
XFILLER_33_38 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_82 vgnd vpwr scs8hd_decap_6
X_135_ address[6] _145_/A vgnd vpwr scs8hd_inv_8
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__186__C _177_/C vgnd vpwr scs8hd_diode_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_12_205 vpwr vgnd scs8hd_fill_2
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_34_81 vpwr vgnd scs8hd_fill_2
X_118_ _118_/A _121_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_29_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_138 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vpwr vgnd scs8hd_fill_2
XANTENNA__183__D _099_/C vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 right_top_grid_pin_13_ mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_119 vgnd vpwr scs8hd_decap_4
XFILLER_32_108 vpwr vgnd scs8hd_fill_2
XFILLER_40_152 vgnd vpwr scs8hd_fill_1
XFILLER_15_83 vgnd vpwr scs8hd_decap_3
XFILLER_16_193 vpwr vgnd scs8hd_fill_2
XFILLER_11_19 vgnd vpwr scs8hd_decap_4
XFILLER_39_252 vgnd vpwr scs8hd_decap_4
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_3_31 vgnd vpwr scs8hd_decap_12
XANTENNA__099__C _099_/C vgnd vpwr scs8hd_diode_2
X_220_ _220_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
X_151_ _122_/A _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XFILLER_33_236 vgnd vpwr scs8hd_decap_8
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_181 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _190_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _214_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_206 vgnd vpwr scs8hd_decap_8
XFILLER_23_50 vgnd vpwr scs8hd_decap_4
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_134_ _123_/A _133_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_7 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_1_.latch data_in _187_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__186__D _102_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_117_ _116_/X _121_/B vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_125 vgnd vpwr scs8hd_fill_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_19 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_191 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_8
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_31_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_14_109 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_175 vgnd vpwr scs8hd_decap_8
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_83 vgnd vpwr scs8hd_decap_8
XFILLER_9_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_76 vgnd vpwr scs8hd_decap_8
XFILLER_3_43 vgnd vpwr scs8hd_decap_6
XFILLER_27_223 vpwr vgnd scs8hd_fill_2
X_150_ _121_/A _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_167 vgnd vpwr scs8hd_decap_4
XFILLER_12_41 vpwr vgnd scs8hd_fill_2
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_237 vgnd vpwr scs8hd_decap_6
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
X_133_ _122_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_270 vgnd vpwr scs8hd_decap_6
XFILLER_23_62 vgnd vpwr scs8hd_fill_1
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_14_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_218 vgnd vpwr scs8hd_decap_12
X_116_ _161_/A _112_/X _145_/C _116_/X vgnd vpwr scs8hd_or3_4
XANTENNA__105__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_148 vgnd vpwr scs8hd_decap_4
XFILLER_30_19 vgnd vpwr scs8hd_fill_1
XFILLER_4_258 vgnd vpwr scs8hd_decap_12
XFILLER_20_41 vpwr vgnd scs8hd_fill_2
XFILLER_20_74 vgnd vpwr scs8hd_fill_1
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_6_54 vgnd vpwr scs8hd_decap_3
XFILLER_6_65 vpwr vgnd scs8hd_fill_2
XFILLER_26_107 vpwr vgnd scs8hd_fill_2
XFILLER_25_19 vgnd vpwr scs8hd_decap_3
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_fill_1
XFILLER_31_95 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_fill_1
XFILLER_31_51 vgnd vpwr scs8hd_decap_4
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XFILLER_16_173 vgnd vpwr scs8hd_decap_12
XFILLER_31_154 vpwr vgnd scs8hd_fill_2
XFILLER_31_132 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_221 vpwr vgnd scs8hd_fill_2
XFILLER_39_210 vpwr vgnd scs8hd_fill_2
XFILLER_22_165 vgnd vpwr scs8hd_fill_1
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_198 vpwr vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_51 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vgnd vpwr scs8hd_decap_4
XFILLER_13_132 vgnd vpwr scs8hd_decap_3
XFILLER_13_176 vgnd vpwr scs8hd_decap_4
XANTENNA__113__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_202 vgnd vpwr scs8hd_decap_6
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_106 vgnd vpwr scs8hd_decap_6
XFILLER_10_124 vpwr vgnd scs8hd_fill_2
XFILLER_5_3 vgnd vpwr scs8hd_decap_6
XFILLER_12_97 vgnd vpwr scs8hd_fill_1
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_37_50 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_224 vpwr vgnd scs8hd_fill_2
XFILLER_37_83 vgnd vpwr scs8hd_decap_12
XFILLER_18_235 vgnd vpwr scs8hd_decap_8
XFILLER_18_246 vgnd vpwr scs8hd_decap_8
XFILLER_18_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_33_19 vgnd vpwr scs8hd_decap_8
XFILLER_32_271 vgnd vpwr scs8hd_decap_4
XFILLER_3_109 vpwr vgnd scs8hd_fill_2
XFILLER_15_205 vpwr vgnd scs8hd_fill_2
X_132_ _121_/A _133_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_74 vpwr vgnd scs8hd_fill_2
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _123_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XFILLER_21_219 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_252 vpwr vgnd scs8hd_fill_2
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_52 vpwr vgnd scs8hd_fill_2
X_115_ _114_/X _145_/C vgnd vpwr scs8hd_buf_1
XFILLER_11_252 vgnd vpwr scs8hd_decap_12
XANTENNA__105__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_29_62 vgnd vpwr scs8hd_decap_3
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XFILLER_20_64 vgnd vpwr scs8hd_decap_4
XFILLER_29_95 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_11 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_196 vgnd vpwr scs8hd_decap_12
XFILLER_34_174 vgnd vpwr scs8hd_decap_12
XFILLER_34_163 vpwr vgnd scs8hd_fill_2
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_130 vpwr vgnd scs8hd_fill_2
XFILLER_17_108 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_163 vgnd vpwr scs8hd_decap_3
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__C _102_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_185 vgnd vpwr scs8hd_fill_1
XFILLER_31_199 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
.ends

