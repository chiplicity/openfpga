VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 29.960 120.000 30.560 ;
    END
  END ccff_tail
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 2.400 99.920 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 34.040 120.000 34.640 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 37.440 120.000 38.040 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 40.840 120.000 41.440 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 44.920 120.000 45.520 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 48.320 120.000 48.920 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 51.720 120.000 52.320 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 55.800 120.000 56.400 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 59.200 120.000 59.800 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 62.600 120.000 63.200 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 66.680 120.000 67.280 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 70.080 120.000 70.680 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 73.480 120.000 74.080 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 77.560 120.000 78.160 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 80.960 120.000 81.560 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 84.360 120.000 84.960 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 88.440 120.000 89.040 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 1.400 120.000 2.000 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 91.840 120.000 92.440 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 4.800 120.000 5.400 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 95.240 120.000 95.840 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 8.200 120.000 8.800 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 99.320 120.000 99.920 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 12.280 120.000 12.880 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 102.720 120.000 103.320 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 15.680 120.000 16.280 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 106.120 120.000 106.720 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 19.080 120.000 19.680 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 110.200 120.000 110.800 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 23.160 120.000 23.760 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 113.600 120.000 114.200 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 26.560 120.000 27.160 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 117.000 120.000 117.600 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 117.600 29.810 120.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 117.600 65.230 120.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 117.600 68.450 120.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 117.600 72.130 120.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 117.600 75.810 120.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 117.600 79.030 120.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.430 117.600 82.710 120.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 117.600 33.490 120.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 117.600 36.710 120.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 117.600 86.390 120.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.330 117.600 89.610 120.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 117.600 93.290 120.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.470 117.600 1.750 120.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 117.600 96.970 120.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 117.600 4.970 120.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 117.600 100.190 120.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 117.600 8.650 120.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 117.600 103.870 120.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.050 117.600 12.330 120.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 117.600 107.550 120.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 117.600 15.550 120.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 117.600 110.770 120.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 117.600 19.230 120.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 117.600 40.390 120.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.170 117.600 114.450 120.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 117.600 22.910 120.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 117.600 118.130 120.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 117.600 26.130 120.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 117.600 44.070 120.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 117.600 47.290 120.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 117.600 50.970 120.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 117.600 54.650 120.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 117.600 57.870 120.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 117.600 61.550 120.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.880 10.640 24.480 109.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.040 10.640 42.640 109.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 114.080 110.415 ;
      LAYER met1 ;
        RECT 1.450 10.240 118.150 114.200 ;
      LAYER met2 ;
        RECT 2.030 117.320 4.410 117.600 ;
        RECT 5.250 117.320 8.090 117.600 ;
        RECT 8.930 117.320 11.770 117.600 ;
        RECT 12.610 117.320 14.990 117.600 ;
        RECT 15.830 117.320 18.670 117.600 ;
        RECT 19.510 117.320 22.350 117.600 ;
        RECT 23.190 117.320 25.570 117.600 ;
        RECT 26.410 117.320 29.250 117.600 ;
        RECT 30.090 117.320 32.930 117.600 ;
        RECT 33.770 117.320 36.150 117.600 ;
        RECT 36.990 117.320 39.830 117.600 ;
        RECT 40.670 117.320 43.510 117.600 ;
        RECT 44.350 117.320 46.730 117.600 ;
        RECT 47.570 117.320 50.410 117.600 ;
        RECT 51.250 117.320 54.090 117.600 ;
        RECT 54.930 117.320 57.310 117.600 ;
        RECT 58.150 117.320 60.990 117.600 ;
        RECT 61.830 117.320 64.670 117.600 ;
        RECT 65.510 117.320 67.890 117.600 ;
        RECT 68.730 117.320 71.570 117.600 ;
        RECT 72.410 117.320 75.250 117.600 ;
        RECT 76.090 117.320 78.470 117.600 ;
        RECT 79.310 117.320 82.150 117.600 ;
        RECT 82.990 117.320 85.830 117.600 ;
        RECT 86.670 117.320 89.050 117.600 ;
        RECT 89.890 117.320 92.730 117.600 ;
        RECT 93.570 117.320 96.410 117.600 ;
        RECT 97.250 117.320 99.630 117.600 ;
        RECT 100.470 117.320 103.310 117.600 ;
        RECT 104.150 117.320 106.990 117.600 ;
        RECT 107.830 117.320 110.210 117.600 ;
        RECT 111.050 117.320 113.890 117.600 ;
        RECT 114.730 117.320 117.570 117.600 ;
        RECT 1.480 2.680 118.120 117.320 ;
        RECT 1.480 1.515 19.590 2.680 ;
        RECT 20.430 1.515 59.610 2.680 ;
        RECT 60.450 1.515 99.630 2.680 ;
        RECT 100.470 1.515 118.120 2.680 ;
      LAYER met3 ;
        RECT 2.400 116.600 117.200 117.465 ;
        RECT 2.400 114.600 117.600 116.600 ;
        RECT 2.400 113.200 117.200 114.600 ;
        RECT 2.400 111.200 117.600 113.200 ;
        RECT 2.400 109.800 117.200 111.200 ;
        RECT 2.400 107.120 117.600 109.800 ;
        RECT 2.400 105.720 117.200 107.120 ;
        RECT 2.400 103.720 117.600 105.720 ;
        RECT 2.400 102.320 117.200 103.720 ;
        RECT 2.400 100.320 117.600 102.320 ;
        RECT 2.800 98.920 117.200 100.320 ;
        RECT 2.400 96.240 117.600 98.920 ;
        RECT 2.400 94.840 117.200 96.240 ;
        RECT 2.400 92.840 117.600 94.840 ;
        RECT 2.400 91.440 117.200 92.840 ;
        RECT 2.400 89.440 117.600 91.440 ;
        RECT 2.400 88.040 117.200 89.440 ;
        RECT 2.400 85.360 117.600 88.040 ;
        RECT 2.400 83.960 117.200 85.360 ;
        RECT 2.400 81.960 117.600 83.960 ;
        RECT 2.400 80.560 117.200 81.960 ;
        RECT 2.400 78.560 117.600 80.560 ;
        RECT 2.400 77.160 117.200 78.560 ;
        RECT 2.400 74.480 117.600 77.160 ;
        RECT 2.400 73.080 117.200 74.480 ;
        RECT 2.400 71.080 117.600 73.080 ;
        RECT 2.400 69.680 117.200 71.080 ;
        RECT 2.400 67.680 117.600 69.680 ;
        RECT 2.400 66.280 117.200 67.680 ;
        RECT 2.400 63.600 117.600 66.280 ;
        RECT 2.400 62.200 117.200 63.600 ;
        RECT 2.400 60.200 117.600 62.200 ;
        RECT 2.800 58.800 117.200 60.200 ;
        RECT 2.400 56.800 117.600 58.800 ;
        RECT 2.400 55.400 117.200 56.800 ;
        RECT 2.400 52.720 117.600 55.400 ;
        RECT 2.400 51.320 117.200 52.720 ;
        RECT 2.400 49.320 117.600 51.320 ;
        RECT 2.400 47.920 117.200 49.320 ;
        RECT 2.400 45.920 117.600 47.920 ;
        RECT 2.400 44.520 117.200 45.920 ;
        RECT 2.400 41.840 117.600 44.520 ;
        RECT 2.400 40.440 117.200 41.840 ;
        RECT 2.400 38.440 117.600 40.440 ;
        RECT 2.400 37.040 117.200 38.440 ;
        RECT 2.400 35.040 117.600 37.040 ;
        RECT 2.400 33.640 117.200 35.040 ;
        RECT 2.400 30.960 117.600 33.640 ;
        RECT 2.400 29.560 117.200 30.960 ;
        RECT 2.400 27.560 117.600 29.560 ;
        RECT 2.400 26.160 117.200 27.560 ;
        RECT 2.400 24.160 117.600 26.160 ;
        RECT 2.400 22.760 117.200 24.160 ;
        RECT 2.400 20.760 117.600 22.760 ;
        RECT 2.800 20.080 117.600 20.760 ;
        RECT 2.800 19.360 117.200 20.080 ;
        RECT 2.400 18.680 117.200 19.360 ;
        RECT 2.400 16.680 117.600 18.680 ;
        RECT 2.400 15.280 117.200 16.680 ;
        RECT 2.400 13.280 117.600 15.280 ;
        RECT 2.400 11.880 117.200 13.280 ;
        RECT 2.400 9.200 117.600 11.880 ;
        RECT 2.400 7.800 117.200 9.200 ;
        RECT 2.400 5.800 117.600 7.800 ;
        RECT 2.400 4.400 117.200 5.800 ;
        RECT 2.400 2.400 117.600 4.400 ;
        RECT 2.400 1.535 117.200 2.400 ;
      LAYER met4 ;
        RECT 20.535 10.240 22.480 109.040 ;
        RECT 24.880 10.240 40.640 109.040 ;
        RECT 43.040 10.240 105.505 109.040 ;
        RECT 20.535 8.335 105.505 10.240 ;
  END
END grid_clb
END LIBRARY

