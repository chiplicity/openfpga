magic
tech EFS8A
magscale 1 2
timestamp 1603804015
<< locali >>
rect 6009 18207 6043 18309
rect 8125 18139 8159 18377
rect 8401 12699 8435 12869
<< viali >>
rect 7849 35241 7883 35275
rect 5457 35105 5491 35139
rect 7665 35105 7699 35139
rect 5641 34969 5675 35003
rect 4997 34697 5031 34731
rect 9689 34697 9723 34731
rect 13645 34697 13679 34731
rect 8585 34629 8619 34663
rect 5181 34493 5215 34527
rect 5733 34493 5767 34527
rect 7757 34493 7791 34527
rect 8401 34493 8435 34527
rect 9045 34493 9079 34527
rect 9505 34493 9539 34527
rect 10057 34493 10091 34527
rect 13461 34493 13495 34527
rect 14013 34493 14047 34527
rect 5365 34357 5399 34391
rect 7113 22389 7147 22423
rect 6688 22049 6722 22083
rect 8033 22049 8067 22083
rect 6791 21981 6825 22015
rect 7665 21981 7699 22015
rect 10517 21641 10551 21675
rect 6653 21573 6687 21607
rect 7481 21505 7515 21539
rect 9020 21437 9054 21471
rect 9505 21437 9539 21471
rect 10333 21437 10367 21471
rect 7573 21369 7607 21403
rect 8125 21369 8159 21403
rect 7205 21301 7239 21335
rect 8401 21301 8435 21335
rect 9091 21301 9125 21335
rect 10885 21301 10919 21335
rect 7389 21097 7423 21131
rect 6929 21029 6963 21063
rect 7941 21029 7975 21063
rect 8493 21029 8527 21063
rect 6837 20961 6871 20995
rect 9756 20961 9790 20995
rect 7849 20893 7883 20927
rect 9827 20757 9861 20791
rect 7665 20553 7699 20587
rect 8861 20553 8895 20587
rect 8401 20485 8435 20519
rect 7849 20417 7883 20451
rect 7941 20281 7975 20315
rect 9137 20281 9171 20315
rect 6285 20213 6319 20247
rect 7297 20213 7331 20247
rect 9781 20213 9815 20247
rect 7941 19941 7975 19975
rect 8033 19941 8067 19975
rect 8309 19805 8343 19839
rect 8217 19465 8251 19499
rect 6653 19261 6687 19295
rect 6929 19261 6963 19295
rect 6837 19193 6871 19227
rect 7941 19125 7975 19159
rect 11299 18921 11333 18955
rect 6745 18853 6779 18887
rect 5616 18785 5650 18819
rect 11196 18785 11230 18819
rect 6653 18717 6687 18751
rect 7205 18649 7239 18683
rect 5687 18581 5721 18615
rect 8401 18581 8435 18615
rect 4859 18377 4893 18411
rect 5641 18377 5675 18411
rect 6653 18377 6687 18411
rect 8125 18377 8159 18411
rect 8217 18377 8251 18411
rect 6009 18309 6043 18343
rect 6193 18309 6227 18343
rect 5273 18241 5307 18275
rect 7297 18241 7331 18275
rect 4788 18173 4822 18207
rect 5784 18173 5818 18207
rect 6009 18173 6043 18207
rect 8493 18241 8527 18275
rect 8769 18241 8803 18275
rect 9873 18173 9907 18207
rect 10149 18173 10183 18207
rect 5871 18105 5905 18139
rect 6929 18105 6963 18139
rect 7021 18105 7055 18139
rect 8125 18105 8159 18139
rect 8585 18105 8619 18139
rect 7849 18037 7883 18071
rect 10241 18037 10275 18071
rect 11161 18037 11195 18071
rect 5457 17833 5491 17867
rect 6469 17833 6503 17867
rect 8493 17833 8527 17867
rect 6745 17765 6779 17799
rect 7297 17765 7331 17799
rect 10333 17765 10367 17799
rect 5641 17697 5675 17731
rect 8309 17697 8343 17731
rect 6653 17629 6687 17663
rect 10241 17629 10275 17663
rect 10609 17629 10643 17663
rect 7573 17493 7607 17527
rect 10057 17493 10091 17527
rect 5089 17289 5123 17323
rect 6285 17289 6319 17323
rect 7757 17289 7791 17323
rect 9873 17289 9907 17323
rect 10977 17289 11011 17323
rect 5641 17221 5675 17255
rect 10609 17221 10643 17255
rect 5733 17153 5767 17187
rect 8953 17153 8987 17187
rect 6837 17085 6871 17119
rect 7158 17017 7192 17051
rect 8309 17017 8343 17051
rect 9505 17017 9539 17051
rect 10057 17017 10091 17051
rect 10149 17017 10183 17051
rect 6561 16949 6595 16983
rect 8125 16745 8159 16779
rect 10609 16745 10643 16779
rect 7567 16677 7601 16711
rect 10010 16677 10044 16711
rect 11621 16677 11655 16711
rect 6228 16609 6262 16643
rect 6331 16609 6365 16643
rect 8401 16609 8435 16643
rect 9689 16609 9723 16643
rect 7205 16541 7239 16575
rect 11529 16541 11563 16575
rect 11805 16541 11839 16575
rect 6837 16405 6871 16439
rect 9413 16405 9447 16439
rect 8585 16201 8619 16235
rect 11069 16201 11103 16235
rect 7113 15997 7147 16031
rect 7481 15997 7515 16031
rect 7665 15997 7699 16031
rect 9413 15997 9447 16031
rect 11196 15997 11230 16031
rect 11621 15997 11655 16031
rect 7986 15929 8020 15963
rect 8953 15929 8987 15963
rect 9775 15929 9809 15963
rect 11299 15929 11333 15963
rect 11989 15929 12023 15963
rect 6193 15861 6227 15895
rect 9229 15861 9263 15895
rect 10333 15861 10367 15895
rect 8401 15657 8435 15691
rect 9413 15657 9447 15691
rect 6653 15589 6687 15623
rect 7843 15589 7877 15623
rect 9873 15589 9907 15623
rect 10425 15589 10459 15623
rect 6009 15521 6043 15555
rect 6469 15521 6503 15555
rect 7481 15453 7515 15487
rect 9781 15453 9815 15487
rect 7297 15317 7331 15351
rect 6009 15113 6043 15147
rect 8217 15113 8251 15147
rect 10333 15113 10367 15147
rect 9597 14977 9631 15011
rect 9873 14977 9907 15011
rect 7113 14909 7147 14943
rect 7481 14909 7515 14943
rect 7665 14909 7699 14943
rect 8769 14909 8803 14943
rect 8953 14909 8987 14943
rect 6377 14773 6411 14807
rect 7297 14773 7331 14807
rect 9781 14569 9815 14603
rect 6187 14501 6221 14535
rect 8769 14501 8803 14535
rect 8125 14433 8159 14467
rect 8493 14433 8527 14467
rect 9689 14433 9723 14467
rect 10241 14433 10275 14467
rect 5825 14365 5859 14399
rect 7205 14365 7239 14399
rect 5273 14229 5307 14263
rect 6745 14229 6779 14263
rect 7573 14229 7607 14263
rect 7757 14025 7791 14059
rect 9873 14025 9907 14059
rect 8493 13957 8527 13991
rect 5089 13889 5123 13923
rect 5273 13889 5307 13923
rect 6653 13821 6687 13855
rect 8677 13821 8711 13855
rect 10333 13821 10367 13855
rect 5365 13753 5399 13787
rect 5917 13753 5951 13787
rect 7113 13753 7147 13787
rect 8998 13753 9032 13787
rect 6193 13685 6227 13719
rect 8125 13685 8159 13719
rect 9597 13685 9631 13719
rect 6469 13481 6503 13515
rect 6929 13481 6963 13515
rect 5226 13413 5260 13447
rect 6837 13345 6871 13379
rect 7389 13345 7423 13379
rect 7481 13345 7515 13379
rect 7849 13345 7883 13379
rect 4905 13277 4939 13311
rect 9689 13277 9723 13311
rect 5825 13141 5859 13175
rect 8677 13141 8711 13175
rect 9137 13141 9171 13175
rect 8401 12869 8435 12903
rect 8677 12869 8711 12903
rect 5917 12801 5951 12835
rect 4629 12733 4663 12767
rect 6285 12733 6319 12767
rect 6653 12733 6687 12767
rect 7113 12733 7147 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 8033 12733 8067 12767
rect 10885 12801 10919 12835
rect 9045 12733 9079 12767
rect 9137 12733 9171 12767
rect 9689 12733 9723 12767
rect 10149 12733 10183 12767
rect 10333 12733 10367 12767
rect 5273 12665 5307 12699
rect 5365 12665 5399 12699
rect 8401 12665 8435 12699
rect 4997 12597 5031 12631
rect 6929 12597 6963 12631
rect 9413 12597 9447 12631
rect 5273 12393 5307 12427
rect 5549 12393 5583 12427
rect 8677 12393 8711 12427
rect 6561 12325 6595 12359
rect 6929 12325 6963 12359
rect 9873 12325 9907 12359
rect 7389 12257 7423 12291
rect 7941 12257 7975 12291
rect 8125 12257 8159 12291
rect 8677 12257 8711 12291
rect 9229 12257 9263 12291
rect 9781 12189 9815 12223
rect 10425 12189 10459 12223
rect 4905 12053 4939 12087
rect 6101 12053 6135 12087
rect 10701 12053 10735 12087
rect 7941 11849 7975 11883
rect 8585 11849 8619 11883
rect 9965 11849 9999 11883
rect 7665 11713 7699 11747
rect 8769 11713 8803 11747
rect 10885 11713 10919 11747
rect 6653 11645 6687 11679
rect 7389 11645 7423 11679
rect 9090 11577 9124 11611
rect 10609 11577 10643 11611
rect 10701 11577 10735 11611
rect 9689 11509 9723 11543
rect 10333 11509 10367 11543
rect 7389 11305 7423 11339
rect 9045 11305 9079 11339
rect 9505 11305 9539 11339
rect 9873 11237 9907 11271
rect 8160 11169 8194 11203
rect 10425 11169 10459 11203
rect 11288 11169 11322 11203
rect 9781 11101 9815 11135
rect 10793 11033 10827 11067
rect 11391 11033 11425 11067
rect 7021 10965 7055 10999
rect 7757 10965 7791 10999
rect 8263 10965 8297 10999
rect 8585 10965 8619 10999
rect 11253 10761 11287 10795
rect 8125 10693 8159 10727
rect 10241 10625 10275 10659
rect 6837 10557 6871 10591
rect 8401 10557 8435 10591
rect 7849 10489 7883 10523
rect 8722 10489 8756 10523
rect 10333 10489 10367 10523
rect 10885 10489 10919 10523
rect 5365 10421 5399 10455
rect 7021 10421 7055 10455
rect 7389 10421 7423 10455
rect 9321 10421 9355 10455
rect 9689 10421 9723 10455
rect 9965 10421 9999 10455
rect 5457 10149 5491 10183
rect 10010 10149 10044 10183
rect 11621 10149 11655 10183
rect 7481 10081 7515 10115
rect 7757 10081 7791 10115
rect 8125 10081 8159 10115
rect 8493 10081 8527 10115
rect 9137 10081 9171 10115
rect 5365 10013 5399 10047
rect 5641 10013 5675 10047
rect 8769 10013 8803 10047
rect 9689 10013 9723 10047
rect 11529 10013 11563 10047
rect 11989 10013 12023 10047
rect 10609 9945 10643 9979
rect 4721 9877 4755 9911
rect 5181 9877 5215 9911
rect 6469 9877 6503 9911
rect 6837 9877 6871 9911
rect 7205 9877 7239 9911
rect 10977 9877 11011 9911
rect 5825 9605 5859 9639
rect 8585 9605 8619 9639
rect 11253 9605 11287 9639
rect 4721 9537 4755 9571
rect 6653 9537 6687 9571
rect 10885 9537 10919 9571
rect 4220 9469 4254 9503
rect 6285 9469 6319 9503
rect 7113 9469 7147 9503
rect 7573 9469 7607 9503
rect 7665 9469 7699 9503
rect 8033 9469 8067 9503
rect 9137 9469 9171 9503
rect 9597 9469 9631 9503
rect 9965 9469 9999 9503
rect 10333 9469 10367 9503
rect 12484 9469 12518 9503
rect 12909 9469 12943 9503
rect 13496 9469 13530 9503
rect 13921 9469 13955 9503
rect 4077 9401 4111 9435
rect 4307 9401 4341 9435
rect 5273 9401 5307 9435
rect 5365 9401 5399 9435
rect 12587 9401 12621 9435
rect 5089 9333 5123 9367
rect 6929 9333 6963 9367
rect 8953 9333 8987 9367
rect 9413 9333 9447 9367
rect 11621 9333 11655 9367
rect 11989 9333 12023 9367
rect 13599 9333 13633 9367
rect 5549 9129 5583 9163
rect 6653 9129 6687 9163
rect 9137 9129 9171 9163
rect 9781 9129 9815 9163
rect 4991 9061 5025 9095
rect 6285 9061 6319 9095
rect 12173 9061 12207 9095
rect 4629 8993 4663 9027
rect 6653 8993 6687 9027
rect 7021 8993 7055 9027
rect 7205 8993 7239 9027
rect 7757 8993 7791 9027
rect 9965 8993 9999 9027
rect 10149 8993 10183 9027
rect 10517 8993 10551 9027
rect 10885 8993 10919 9027
rect 13588 8993 13622 9027
rect 12081 8925 12115 8959
rect 12357 8925 12391 8959
rect 5917 8789 5951 8823
rect 8125 8789 8159 8823
rect 8769 8789 8803 8823
rect 13691 8789 13725 8823
rect 4307 8585 4341 8619
rect 6469 8585 6503 8619
rect 9137 8585 9171 8619
rect 11253 8585 11287 8619
rect 12081 8585 12115 8619
rect 7297 8517 7331 8551
rect 10885 8517 10919 8551
rect 13553 8517 13587 8551
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 4220 8381 4254 8415
rect 7665 8381 7699 8415
rect 8125 8381 8159 8415
rect 8309 8381 8343 8415
rect 8585 8381 8619 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 12484 8381 12518 8415
rect 12909 8381 12943 8415
rect 5365 8313 5399 8347
rect 10010 8313 10044 8347
rect 11621 8313 11655 8347
rect 12587 8313 12621 8347
rect 4629 8245 4663 8279
rect 5089 8245 5123 8279
rect 8769 8245 8803 8279
rect 10609 8245 10643 8279
rect 4629 8041 4663 8075
rect 7665 8041 7699 8075
rect 8033 8041 8067 8075
rect 8677 8041 8711 8075
rect 9045 8041 9079 8075
rect 6054 7973 6088 8007
rect 8401 7973 8435 8007
rect 9413 7973 9447 8007
rect 9873 7973 9907 8007
rect 11437 7973 11471 8007
rect 5273 7905 5307 7939
rect 6653 7905 6687 7939
rect 7481 7905 7515 7939
rect 8493 7905 8527 7939
rect 5733 7837 5767 7871
rect 7021 7837 7055 7871
rect 7389 7837 7423 7871
rect 9781 7837 9815 7871
rect 10425 7837 10459 7871
rect 11345 7837 11379 7871
rect 11897 7769 11931 7803
rect 5641 7701 5675 7735
rect 6193 7497 6227 7531
rect 9597 7497 9631 7531
rect 9873 7497 9907 7531
rect 11897 7497 11931 7531
rect 7573 7361 7607 7395
rect 10517 7361 10551 7395
rect 10793 7361 10827 7395
rect 6929 7293 6963 7327
rect 8677 7293 8711 7327
rect 7849 7225 7883 7259
rect 8998 7225 9032 7259
rect 10609 7225 10643 7259
rect 5733 7157 5767 7191
rect 6653 7157 6687 7191
rect 8493 7157 8527 7191
rect 10333 7157 10367 7191
rect 11437 7157 11471 7191
rect 9137 6953 9171 6987
rect 10149 6953 10183 6987
rect 10517 6953 10551 6987
rect 4972 6817 5006 6851
rect 7297 6817 7331 6851
rect 9724 6817 9758 6851
rect 9827 6817 9861 6851
rect 5043 6681 5077 6715
rect 7481 6681 7515 6715
rect 8677 6613 8711 6647
rect 4353 6409 4387 6443
rect 7205 6409 7239 6443
rect 7941 6409 7975 6443
rect 8677 6409 8711 6443
rect 7021 6205 7055 6239
rect 8493 6205 8527 6239
rect 4721 6137 4755 6171
rect 5273 6137 5307 6171
rect 5365 6137 5399 6171
rect 5917 6137 5951 6171
rect 9689 6137 9723 6171
rect 5089 6069 5123 6103
rect 6561 6069 6595 6103
rect 9045 6069 9079 6103
rect 4399 5865 4433 5899
rect 6929 5865 6963 5899
rect 7297 5865 7331 5899
rect 5181 5797 5215 5831
rect 5457 5797 5491 5831
rect 4296 5729 4330 5763
rect 6561 5729 6595 5763
rect 7297 5729 7331 5763
rect 7573 5729 7607 5763
rect 7849 5729 7883 5763
rect 8217 5729 8251 5763
rect 5365 5661 5399 5695
rect 5825 5661 5859 5695
rect 4813 5525 4847 5559
rect 3111 5321 3145 5355
rect 3893 5321 3927 5355
rect 4445 5321 4479 5355
rect 5917 5321 5951 5355
rect 3525 5253 3559 5287
rect 9965 5253 9999 5287
rect 8585 5185 8619 5219
rect 3040 5117 3074 5151
rect 4036 5117 4070 5151
rect 4997 5117 5031 5151
rect 6653 5117 6687 5151
rect 7021 5117 7055 5151
rect 7389 5117 7423 5151
rect 7665 5117 7699 5151
rect 8217 5117 8251 5151
rect 9781 5117 9815 5151
rect 10333 5117 10367 5151
rect 5359 5049 5393 5083
rect 4123 4981 4157 5015
rect 4905 4981 4939 5015
rect 6285 4981 6319 5015
rect 6929 4981 6963 5015
rect 8953 4981 8987 5015
rect 8217 4777 8251 4811
rect 5641 4709 5675 4743
rect 4480 4641 4514 4675
rect 7297 4641 7331 4675
rect 7665 4641 7699 4675
rect 7849 4641 7883 4675
rect 8309 4641 8343 4675
rect 5549 4573 5583 4607
rect 5825 4573 5859 4607
rect 5089 4505 5123 4539
rect 4353 4437 4387 4471
rect 4583 4437 4617 4471
rect 6469 4437 6503 4471
rect 6929 4437 6963 4471
rect 8769 4437 8803 4471
rect 3801 4233 3835 4267
rect 4445 4233 4479 4267
rect 8125 4233 8159 4267
rect 8861 4165 8895 4199
rect 5273 4097 5307 4131
rect 5917 4097 5951 4131
rect 6285 4097 6319 4131
rect 8732 4097 8766 4131
rect 8953 4097 8987 4131
rect 9321 4097 9355 4131
rect 10609 4097 10643 4131
rect 5089 4029 5123 4063
rect 7205 4029 7239 4063
rect 7757 4029 7791 4063
rect 9689 4029 9723 4063
rect 10333 4029 10367 4063
rect 10977 4029 11011 4063
rect 13461 4029 13495 4063
rect 14013 4029 14047 4063
rect 4169 3961 4203 3995
rect 5365 3961 5399 3995
rect 8585 3961 8619 3995
rect 10149 3961 10183 3995
rect 6653 3893 6687 3927
rect 8493 3893 8527 3927
rect 9965 3893 9999 3927
rect 13645 3893 13679 3927
rect 4905 3689 4939 3723
rect 6745 3689 6779 3723
rect 10333 3689 10367 3723
rect 11437 3689 11471 3723
rect 6187 3621 6221 3655
rect 7113 3621 7147 3655
rect 7573 3553 7607 3587
rect 8953 3553 8987 3587
rect 9689 3553 9723 3587
rect 11253 3553 11287 3587
rect 13461 3553 13495 3587
rect 4537 3485 4571 3519
rect 5825 3485 5859 3519
rect 7941 3485 7975 3519
rect 10057 3485 10091 3519
rect 7389 3417 7423 3451
rect 7738 3417 7772 3451
rect 5273 3349 5307 3383
rect 5549 3349 5583 3383
rect 7849 3349 7883 3383
rect 8033 3349 8067 3383
rect 8677 3349 8711 3383
rect 9413 3349 9447 3383
rect 9827 3349 9861 3383
rect 9965 3349 9999 3383
rect 13645 3349 13679 3383
rect 4077 3145 4111 3179
rect 5346 3145 5380 3179
rect 5825 3145 5859 3179
rect 7757 3145 7791 3179
rect 8585 3145 8619 3179
rect 8861 3145 8895 3179
rect 10425 3145 10459 3179
rect 10793 3145 10827 3179
rect 11529 3145 11563 3179
rect 13001 3145 13035 3179
rect 13461 3145 13495 3179
rect 4721 3077 4755 3111
rect 5457 3077 5491 3111
rect 10057 3077 10091 3111
rect 11161 3077 11195 3111
rect 12633 3077 12667 3111
rect 5089 3009 5123 3043
rect 5549 3009 5583 3043
rect 6653 3009 6687 3043
rect 7389 3009 7423 3043
rect 9045 3009 9079 3043
rect 4169 2941 4203 2975
rect 8125 2941 8159 2975
rect 9137 2941 9171 2975
rect 10977 2941 11011 2975
rect 12449 2941 12483 2975
rect 5181 2873 5215 2907
rect 4353 2805 4387 2839
rect 6285 2805 6319 2839
rect 4813 2601 4847 2635
rect 7021 2601 7055 2635
rect 9505 2601 9539 2635
rect 13277 2601 13311 2635
rect 5273 2533 5307 2567
rect 4169 2465 4203 2499
rect 5181 2465 5215 2499
rect 5825 2465 5859 2499
rect 6377 2465 6411 2499
rect 7021 2465 7055 2499
rect 7665 2465 7699 2499
rect 7757 2465 7791 2499
rect 8309 2465 8343 2499
rect 9045 2465 9079 2499
rect 9781 2465 9815 2499
rect 10333 2465 10367 2499
rect 10885 2465 10919 2499
rect 11437 2465 11471 2499
rect 13093 2465 13127 2499
rect 13645 2465 13679 2499
rect 8677 2397 8711 2431
rect 4353 2329 4387 2363
rect 9965 2329 9999 2363
rect 11069 2329 11103 2363
rect 6653 2261 6687 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 8478 35640 8484 35692
rect 8536 35680 8542 35692
rect 9306 35680 9312 35692
rect 8536 35652 9312 35680
rect 8536 35640 8542 35652
rect 9306 35640 9312 35652
rect 9364 35640 9370 35692
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 7837 35275 7895 35281
rect 7837 35241 7849 35275
rect 7883 35272 7895 35275
rect 8202 35272 8208 35284
rect 7883 35244 8208 35272
rect 7883 35241 7895 35244
rect 7837 35235 7895 35241
rect 8202 35232 8208 35244
rect 8260 35232 8266 35284
rect 5445 35139 5503 35145
rect 5445 35105 5457 35139
rect 5491 35136 5503 35139
rect 5534 35136 5540 35148
rect 5491 35108 5540 35136
rect 5491 35105 5503 35108
rect 5445 35099 5503 35105
rect 5534 35096 5540 35108
rect 5592 35096 5598 35148
rect 5626 35096 5632 35148
rect 5684 35136 5690 35148
rect 5810 35136 5816 35148
rect 5684 35108 5816 35136
rect 5684 35096 5690 35108
rect 5810 35096 5816 35108
rect 5868 35096 5874 35148
rect 7650 35136 7656 35148
rect 7611 35108 7656 35136
rect 7650 35096 7656 35108
rect 7708 35096 7714 35148
rect 5626 35000 5632 35012
rect 5587 34972 5632 35000
rect 5626 34960 5632 34972
rect 5684 34960 5690 35012
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 4798 34688 4804 34740
rect 4856 34728 4862 34740
rect 4985 34731 5043 34737
rect 4985 34728 4997 34731
rect 4856 34700 4997 34728
rect 4856 34688 4862 34700
rect 4985 34697 4997 34700
rect 5031 34697 5043 34731
rect 4985 34691 5043 34697
rect 9677 34731 9735 34737
rect 9677 34697 9689 34731
rect 9723 34728 9735 34731
rect 10962 34728 10968 34740
rect 9723 34700 10968 34728
rect 9723 34697 9735 34700
rect 9677 34691 9735 34697
rect 5000 34524 5028 34691
rect 10962 34688 10968 34700
rect 11020 34688 11026 34740
rect 13630 34728 13636 34740
rect 13591 34700 13636 34728
rect 13630 34688 13636 34700
rect 13688 34688 13694 34740
rect 8573 34663 8631 34669
rect 8573 34629 8585 34663
rect 8619 34660 8631 34663
rect 10134 34660 10140 34672
rect 8619 34632 10140 34660
rect 8619 34629 8631 34632
rect 8573 34623 8631 34629
rect 10134 34620 10140 34632
rect 10192 34620 10198 34672
rect 5169 34527 5227 34533
rect 5169 34524 5181 34527
rect 5000 34496 5181 34524
rect 5169 34493 5181 34496
rect 5215 34493 5227 34527
rect 5169 34487 5227 34493
rect 5534 34484 5540 34536
rect 5592 34524 5598 34536
rect 5721 34527 5779 34533
rect 5721 34524 5733 34527
rect 5592 34496 5733 34524
rect 5592 34484 5598 34496
rect 5721 34493 5733 34496
rect 5767 34493 5779 34527
rect 5721 34487 5779 34493
rect 7650 34484 7656 34536
rect 7708 34524 7714 34536
rect 7745 34527 7803 34533
rect 7745 34524 7757 34527
rect 7708 34496 7757 34524
rect 7708 34484 7714 34496
rect 7745 34493 7757 34496
rect 7791 34524 7803 34527
rect 8202 34524 8208 34536
rect 7791 34496 8208 34524
rect 7791 34493 7803 34496
rect 7745 34487 7803 34493
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 8389 34527 8447 34533
rect 8389 34493 8401 34527
rect 8435 34524 8447 34527
rect 9033 34527 9091 34533
rect 9033 34524 9045 34527
rect 8435 34496 9045 34524
rect 8435 34493 8447 34496
rect 8389 34487 8447 34493
rect 9033 34493 9045 34496
rect 9079 34524 9091 34527
rect 9306 34524 9312 34536
rect 9079 34496 9312 34524
rect 9079 34493 9091 34496
rect 9033 34487 9091 34493
rect 9306 34484 9312 34496
rect 9364 34484 9370 34536
rect 9490 34524 9496 34536
rect 9451 34496 9496 34524
rect 9490 34484 9496 34496
rect 9548 34524 9554 34536
rect 10045 34527 10103 34533
rect 10045 34524 10057 34527
rect 9548 34496 10057 34524
rect 9548 34484 9554 34496
rect 10045 34493 10057 34496
rect 10091 34493 10103 34527
rect 10045 34487 10103 34493
rect 12526 34484 12532 34536
rect 12584 34524 12590 34536
rect 13449 34527 13507 34533
rect 13449 34524 13461 34527
rect 12584 34496 13461 34524
rect 12584 34484 12590 34496
rect 13449 34493 13461 34496
rect 13495 34524 13507 34527
rect 14001 34527 14059 34533
rect 14001 34524 14013 34527
rect 13495 34496 14013 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 14001 34493 14013 34496
rect 14047 34493 14059 34527
rect 14001 34487 14059 34493
rect 5350 34388 5356 34400
rect 5311 34360 5356 34388
rect 5350 34348 5356 34360
rect 5408 34348 5414 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 2130 31696 2136 31748
rect 2188 31736 2194 31748
rect 3970 31736 3976 31748
rect 2188 31708 3976 31736
rect 2188 31696 2194 31708
rect 3970 31696 3976 31708
rect 4028 31696 4034 31748
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 5718 29044 5724 29096
rect 5776 29084 5782 29096
rect 5810 29084 5816 29096
rect 5776 29056 5816 29084
rect 5776 29044 5782 29056
rect 5810 29044 5816 29056
rect 5868 29044 5874 29096
rect 3142 28976 3148 29028
rect 3200 29016 3206 29028
rect 3510 29016 3516 29028
rect 3200 28988 3516 29016
rect 3200 28976 3206 28988
rect 3510 28976 3516 28988
rect 3568 28976 3574 29028
rect 12710 28976 12716 29028
rect 12768 29016 12774 29028
rect 12802 29016 12808 29028
rect 12768 28988 12808 29016
rect 12768 28976 12774 28988
rect 12802 28976 12808 28988
rect 12860 28976 12866 29028
rect 3970 28908 3976 28960
rect 4028 28948 4034 28960
rect 4338 28948 4344 28960
rect 4028 28920 4344 28948
rect 4028 28908 4034 28920
rect 4338 28908 4344 28920
rect 4396 28908 4402 28960
rect 8662 28908 8668 28960
rect 8720 28948 8726 28960
rect 9306 28948 9312 28960
rect 8720 28920 9312 28948
rect 8720 28908 8726 28920
rect 9306 28908 9312 28920
rect 9364 28908 9370 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 5258 27548 5264 27600
rect 5316 27588 5322 27600
rect 5718 27588 5724 27600
rect 5316 27560 5724 27588
rect 5316 27548 5322 27560
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 106 26868 112 26920
rect 164 26908 170 26920
rect 1302 26908 1308 26920
rect 164 26880 1308 26908
rect 164 26868 170 26880
rect 1302 26868 1308 26880
rect 1360 26868 1366 26920
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 7098 22420 7104 22432
rect 7059 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 14 22108 20 22160
rect 72 22148 78 22160
rect 382 22148 388 22160
rect 72 22120 388 22148
rect 72 22108 78 22120
rect 382 22108 388 22120
rect 440 22108 446 22160
rect 6638 22040 6644 22092
rect 6696 22089 6702 22092
rect 6696 22083 6734 22089
rect 6722 22049 6734 22083
rect 8018 22080 8024 22092
rect 7979 22052 8024 22080
rect 6696 22043 6734 22049
rect 6696 22040 6702 22043
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 6779 22015 6837 22021
rect 6779 22012 6791 22015
rect 6604 21984 6791 22012
rect 6604 21972 6610 21984
rect 6779 21981 6791 21984
rect 6825 21981 6837 22015
rect 7650 22012 7656 22024
rect 7611 21984 7656 22012
rect 6779 21975 6837 21981
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 10502 21672 10508 21684
rect 10463 21644 10508 21672
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 6638 21604 6644 21616
rect 6551 21576 6644 21604
rect 6638 21564 6644 21576
rect 6696 21604 6702 21616
rect 8110 21604 8116 21616
rect 6696 21576 8116 21604
rect 6696 21564 6702 21576
rect 8110 21564 8116 21576
rect 8168 21564 8174 21616
rect 7098 21496 7104 21548
rect 7156 21536 7162 21548
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 7156 21508 7481 21536
rect 7156 21496 7162 21508
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 9008 21471 9066 21477
rect 9008 21437 9020 21471
rect 9054 21468 9066 21471
rect 9493 21471 9551 21477
rect 9493 21468 9505 21471
rect 9054 21440 9505 21468
rect 9054 21437 9066 21440
rect 9008 21431 9066 21437
rect 9493 21437 9505 21440
rect 9539 21468 9551 21471
rect 10321 21471 10379 21477
rect 10321 21468 10333 21471
rect 9539 21440 10333 21468
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 10321 21437 10333 21440
rect 10367 21468 10379 21471
rect 10367 21440 10824 21468
rect 10367 21437 10379 21440
rect 10321 21431 10379 21437
rect 7561 21403 7619 21409
rect 7561 21369 7573 21403
rect 7607 21369 7619 21403
rect 8110 21400 8116 21412
rect 8071 21372 8116 21400
rect 7561 21363 7619 21369
rect 7190 21332 7196 21344
rect 7151 21304 7196 21332
rect 7190 21292 7196 21304
rect 7248 21332 7254 21344
rect 7576 21332 7604 21363
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 10796 21344 10824 21440
rect 7248 21304 7604 21332
rect 7248 21292 7254 21304
rect 8018 21292 8024 21344
rect 8076 21332 8082 21344
rect 8389 21335 8447 21341
rect 8389 21332 8401 21335
rect 8076 21304 8401 21332
rect 8076 21292 8082 21304
rect 8389 21301 8401 21304
rect 8435 21301 8447 21335
rect 8389 21295 8447 21301
rect 8570 21292 8576 21344
rect 8628 21332 8634 21344
rect 9079 21335 9137 21341
rect 9079 21332 9091 21335
rect 8628 21304 9091 21332
rect 8628 21292 8634 21304
rect 9079 21301 9091 21304
rect 9125 21301 9137 21335
rect 9079 21295 9137 21301
rect 10778 21292 10784 21344
rect 10836 21332 10842 21344
rect 10873 21335 10931 21341
rect 10873 21332 10885 21335
rect 10836 21304 10885 21332
rect 10836 21292 10842 21304
rect 10873 21301 10885 21304
rect 10919 21301 10931 21335
rect 10873 21295 10931 21301
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 7098 21088 7104 21140
rect 7156 21128 7162 21140
rect 7377 21131 7435 21137
rect 7377 21128 7389 21131
rect 7156 21100 7389 21128
rect 7156 21088 7162 21100
rect 7377 21097 7389 21100
rect 7423 21097 7435 21131
rect 7377 21091 7435 21097
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21060 6975 21063
rect 7190 21060 7196 21072
rect 6963 21032 7196 21060
rect 6963 21029 6975 21032
rect 6917 21023 6975 21029
rect 7190 21020 7196 21032
rect 7248 21020 7254 21072
rect 7926 21060 7932 21072
rect 7300 21032 7932 21060
rect 6825 20995 6883 21001
rect 6825 20961 6837 20995
rect 6871 20992 6883 20995
rect 7300 20992 7328 21032
rect 7926 21020 7932 21032
rect 7984 21020 7990 21072
rect 8110 21020 8116 21072
rect 8168 21060 8174 21072
rect 8481 21063 8539 21069
rect 8481 21060 8493 21063
rect 8168 21032 8493 21060
rect 8168 21020 8174 21032
rect 8481 21029 8493 21032
rect 8527 21029 8539 21063
rect 8481 21023 8539 21029
rect 9766 21001 9772 21004
rect 6871 20964 7328 20992
rect 9744 20995 9772 21001
rect 6871 20961 6883 20964
rect 6825 20955 6883 20961
rect 9744 20961 9756 20995
rect 9744 20955 9772 20961
rect 9766 20952 9772 20955
rect 9824 20952 9830 21004
rect 7837 20927 7895 20933
rect 7837 20893 7849 20927
rect 7883 20924 7895 20927
rect 8294 20924 8300 20936
rect 7883 20896 8300 20924
rect 7883 20893 7895 20896
rect 7837 20887 7895 20893
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9815 20791 9873 20797
rect 9815 20788 9827 20791
rect 9732 20760 9827 20788
rect 9732 20748 9738 20760
rect 9815 20757 9827 20760
rect 9861 20757 9873 20791
rect 9815 20751 9873 20757
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 7650 20584 7656 20596
rect 7611 20556 7656 20584
rect 7650 20544 7656 20556
rect 7708 20544 7714 20596
rect 8849 20587 8907 20593
rect 8849 20553 8861 20587
rect 8895 20584 8907 20587
rect 9582 20584 9588 20596
rect 8895 20556 9588 20584
rect 8895 20553 8907 20556
rect 8849 20547 8907 20553
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8389 20519 8447 20525
rect 8389 20516 8401 20519
rect 8352 20488 8401 20516
rect 8352 20476 8358 20488
rect 8389 20485 8401 20488
rect 8435 20485 8447 20519
rect 8389 20479 8447 20485
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20448 7895 20451
rect 8864 20448 8892 20547
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 7883 20420 8892 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20281 7987 20315
rect 7929 20275 7987 20281
rect 6273 20247 6331 20253
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 7282 20244 7288 20256
rect 6319 20216 7288 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 7944 20244 7972 20275
rect 8294 20272 8300 20324
rect 8352 20312 8358 20324
rect 9125 20315 9183 20321
rect 9125 20312 9137 20315
rect 8352 20284 9137 20312
rect 8352 20272 8358 20284
rect 9125 20281 9137 20284
rect 9171 20281 9183 20315
rect 9125 20275 9183 20281
rect 9766 20244 9772 20256
rect 7708 20216 7972 20244
rect 9679 20216 9772 20244
rect 7708 20204 7714 20216
rect 9766 20204 9772 20216
rect 9824 20244 9830 20256
rect 10962 20244 10968 20256
rect 9824 20216 10968 20244
rect 9824 20204 9830 20216
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 8110 20040 8116 20052
rect 7944 20012 8116 20040
rect 7944 19981 7972 20012
rect 8110 20000 8116 20012
rect 8168 20040 8174 20052
rect 8570 20040 8576 20052
rect 8168 20012 8576 20040
rect 8168 20000 8174 20012
rect 8570 20000 8576 20012
rect 8628 20000 8634 20052
rect 7929 19975 7987 19981
rect 7929 19941 7941 19975
rect 7975 19941 7987 19975
rect 7929 19935 7987 19941
rect 8018 19932 8024 19984
rect 8076 19972 8082 19984
rect 8076 19944 8121 19972
rect 8076 19932 8082 19944
rect 8294 19836 8300 19848
rect 8255 19808 8300 19836
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 8205 19499 8263 19505
rect 8205 19496 8217 19499
rect 8168 19468 8217 19496
rect 8168 19456 8174 19468
rect 8205 19465 8217 19468
rect 8251 19465 8263 19499
rect 8205 19459 8263 19465
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4338 19360 4344 19372
rect 4120 19332 4344 19360
rect 4120 19320 4126 19332
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 8754 19360 8760 19372
rect 8720 19332 8760 19360
rect 8720 19320 8726 19332
rect 8754 19320 8760 19332
rect 8812 19320 8818 19372
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 12894 19360 12900 19372
rect 12676 19332 12900 19360
rect 12676 19320 12682 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6914 19292 6920 19304
rect 6687 19264 6920 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 12526 19292 12532 19304
rect 12400 19264 12532 19292
rect 12400 19252 12406 19264
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 6822 19224 6828 19236
rect 6783 19196 6828 19224
rect 6822 19184 6828 19196
rect 6880 19184 6886 19236
rect 7929 19159 7987 19165
rect 7929 19125 7941 19159
rect 7975 19156 7987 19159
rect 8018 19156 8024 19168
rect 7975 19128 8024 19156
rect 7975 19125 7987 19128
rect 7929 19119 7987 19125
rect 8018 19116 8024 19128
rect 8076 19156 8082 19168
rect 8386 19156 8392 19168
rect 8076 19128 8392 19156
rect 8076 19116 8082 19128
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 9490 18952 9496 18964
rect 6288 18924 9496 18952
rect 5626 18825 5632 18828
rect 5604 18819 5632 18825
rect 5604 18816 5616 18819
rect 5539 18788 5616 18816
rect 5604 18785 5616 18788
rect 5684 18816 5690 18828
rect 6288 18816 6316 18924
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 11330 18961 11336 18964
rect 11287 18955 11336 18961
rect 11287 18921 11299 18955
rect 11333 18921 11336 18955
rect 11287 18915 11336 18921
rect 11330 18912 11336 18915
rect 11388 18912 11394 18964
rect 6733 18887 6791 18893
rect 6733 18853 6745 18887
rect 6779 18884 6791 18887
rect 6822 18884 6828 18896
rect 6779 18856 6828 18884
rect 6779 18853 6791 18856
rect 6733 18847 6791 18853
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 5684 18788 6316 18816
rect 5604 18779 5632 18785
rect 5626 18776 5632 18779
rect 5684 18776 5690 18788
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11184 18819 11242 18825
rect 11184 18816 11196 18819
rect 11112 18788 11196 18816
rect 11112 18776 11118 18788
rect 11184 18785 11196 18788
rect 11230 18785 11242 18819
rect 11184 18779 11242 18785
rect 6638 18748 6644 18760
rect 6599 18720 6644 18748
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 7190 18680 7196 18692
rect 7151 18652 7196 18680
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 5675 18615 5733 18621
rect 5675 18581 5687 18615
rect 5721 18612 5733 18615
rect 8294 18612 8300 18624
rect 5721 18584 8300 18612
rect 5721 18581 5733 18584
rect 5675 18575 5733 18581
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 8389 18615 8447 18621
rect 8389 18612 8401 18615
rect 8352 18584 8401 18612
rect 8352 18572 8358 18584
rect 8389 18581 8401 18584
rect 8435 18581 8447 18615
rect 8389 18575 8447 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4847 18411 4905 18417
rect 4847 18408 4859 18411
rect 4212 18380 4859 18408
rect 4212 18368 4218 18380
rect 4847 18377 4859 18380
rect 4893 18377 4905 18411
rect 5626 18408 5632 18420
rect 5587 18380 5632 18408
rect 4847 18371 4905 18377
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 6822 18408 6828 18420
rect 6687 18380 6828 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 6972 18380 8125 18408
rect 6972 18368 6978 18380
rect 8113 18377 8125 18380
rect 8159 18408 8171 18411
rect 8205 18411 8263 18417
rect 8205 18408 8217 18411
rect 8159 18380 8217 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 8205 18377 8217 18380
rect 8251 18377 8263 18411
rect 8205 18371 8263 18377
rect 3050 18300 3056 18352
rect 3108 18340 3114 18352
rect 5810 18340 5816 18352
rect 3108 18312 5816 18340
rect 3108 18300 3114 18312
rect 5810 18300 5816 18312
rect 5868 18340 5874 18352
rect 5997 18343 6055 18349
rect 5997 18340 6009 18343
rect 5868 18312 6009 18340
rect 5868 18300 5874 18312
rect 5997 18309 6009 18312
rect 6043 18340 6055 18343
rect 6181 18343 6239 18349
rect 6181 18340 6193 18343
rect 6043 18312 6193 18340
rect 6043 18309 6055 18312
rect 5997 18303 6055 18309
rect 6181 18309 6193 18312
rect 6227 18309 6239 18343
rect 6181 18303 6239 18309
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7248 18312 8800 18340
rect 7248 18300 7254 18312
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18272 5319 18275
rect 7282 18272 7288 18284
rect 5307 18244 7288 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 4776 18207 4834 18213
rect 4776 18173 4788 18207
rect 4822 18204 4834 18207
rect 5276 18204 5304 18235
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8772 18281 8800 18312
rect 8481 18275 8539 18281
rect 8481 18272 8493 18275
rect 8352 18244 8493 18272
rect 8352 18232 8358 18244
rect 8481 18241 8493 18244
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18241 8815 18275
rect 8757 18235 8815 18241
rect 4822 18176 5304 18204
rect 5772 18207 5830 18213
rect 4822 18173 4834 18176
rect 4776 18167 4834 18173
rect 5772 18173 5784 18207
rect 5818 18204 5830 18207
rect 5997 18207 6055 18213
rect 5997 18204 6009 18207
rect 5818 18176 6009 18204
rect 5818 18173 5830 18176
rect 5772 18167 5830 18173
rect 5997 18173 6009 18176
rect 6043 18173 6055 18207
rect 5997 18167 6055 18173
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18204 9919 18207
rect 10134 18204 10140 18216
rect 9907 18176 10140 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 5859 18139 5917 18145
rect 5859 18105 5871 18139
rect 5905 18136 5917 18139
rect 6638 18136 6644 18148
rect 5905 18108 6644 18136
rect 5905 18105 5917 18108
rect 5859 18099 5917 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 6914 18136 6920 18148
rect 6875 18108 6920 18136
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 7098 18136 7104 18148
rect 7055 18108 7104 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 8110 18136 8116 18148
rect 8023 18108 8116 18136
rect 8110 18096 8116 18108
rect 8168 18136 8174 18148
rect 8573 18139 8631 18145
rect 8573 18136 8585 18139
rect 8168 18108 8585 18136
rect 8168 18096 8174 18108
rect 8573 18105 8585 18108
rect 8619 18105 8631 18139
rect 8573 18099 8631 18105
rect 7116 18068 7144 18096
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7116 18040 7849 18068
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 10226 18068 10232 18080
rect 10187 18040 10232 18068
rect 7837 18031 7895 18037
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 11112 18040 11161 18068
rect 11112 18028 11118 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 5442 17864 5448 17876
rect 5403 17836 5448 17864
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 6457 17867 6515 17873
rect 6457 17833 6469 17867
rect 6503 17864 6515 17867
rect 6638 17864 6644 17876
rect 6503 17836 6644 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 6733 17799 6791 17805
rect 6733 17796 6745 17799
rect 5644 17768 6745 17796
rect 5644 17737 5672 17768
rect 6733 17765 6745 17768
rect 6779 17796 6791 17799
rect 6822 17796 6828 17808
rect 6779 17768 6828 17796
rect 6779 17765 6791 17768
rect 6733 17759 6791 17765
rect 6822 17756 6828 17768
rect 6880 17756 6886 17808
rect 7282 17796 7288 17808
rect 7243 17768 7288 17796
rect 7282 17756 7288 17768
rect 7340 17756 7346 17808
rect 10226 17756 10232 17808
rect 10284 17796 10290 17808
rect 10321 17799 10379 17805
rect 10321 17796 10333 17799
rect 10284 17768 10333 17796
rect 10284 17756 10290 17768
rect 10321 17765 10333 17768
rect 10367 17765 10379 17799
rect 10321 17759 10379 17765
rect 5629 17731 5687 17737
rect 5629 17697 5641 17731
rect 5675 17697 5687 17731
rect 8294 17728 8300 17740
rect 8255 17700 8300 17728
rect 5629 17691 5687 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 6638 17660 6644 17672
rect 6599 17632 6644 17660
rect 6638 17620 6644 17632
rect 6696 17660 6702 17672
rect 7098 17660 7104 17672
rect 6696 17632 7104 17660
rect 6696 17620 6702 17632
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 9916 17632 10241 17660
rect 9916 17620 9922 17632
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 10229 17623 10287 17629
rect 10594 17620 10600 17632
rect 10652 17660 10658 17672
rect 11054 17660 11060 17672
rect 10652 17632 11060 17660
rect 10652 17620 10658 17632
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7561 17527 7619 17533
rect 7561 17524 7573 17527
rect 6972 17496 7573 17524
rect 6972 17484 6978 17496
rect 7561 17493 7573 17496
rect 7607 17493 7619 17527
rect 7561 17487 7619 17493
rect 10045 17527 10103 17533
rect 10045 17493 10057 17527
rect 10091 17524 10103 17527
rect 10134 17524 10140 17536
rect 10091 17496 10140 17524
rect 10091 17493 10103 17496
rect 10045 17487 10103 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 6273 17323 6331 17329
rect 6273 17320 6285 17323
rect 5123 17292 6285 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 6273 17289 6285 17292
rect 6319 17320 6331 17323
rect 6822 17320 6828 17332
rect 6319 17292 6828 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6822 17280 6828 17292
rect 6880 17320 6886 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 6880 17292 7757 17320
rect 6880 17280 6886 17292
rect 7745 17289 7757 17292
rect 7791 17289 7803 17323
rect 9858 17320 9864 17332
rect 7745 17283 7803 17289
rect 8956 17292 9864 17320
rect 5629 17255 5687 17261
rect 5629 17221 5641 17255
rect 5675 17252 5687 17255
rect 6638 17252 6644 17264
rect 5675 17224 6644 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 5721 17187 5779 17193
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 6914 17184 6920 17196
rect 5767 17156 6920 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 8956 17193 8984 17292
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10284 17292 10977 17320
rect 10284 17280 10290 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 10965 17283 11023 17289
rect 10594 17252 10600 17264
rect 10555 17224 10600 17252
rect 10594 17212 10600 17224
rect 10652 17212 10658 17264
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6696 17088 6837 17116
rect 6696 17076 6702 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7146 17051 7204 17057
rect 7146 17048 7158 17051
rect 6564 17020 7158 17048
rect 6178 16940 6184 16992
rect 6236 16980 6242 16992
rect 6564 16989 6592 17020
rect 7146 17017 7158 17020
rect 7192 17017 7204 17051
rect 8294 17048 8300 17060
rect 8255 17020 8300 17048
rect 7146 17011 7204 17017
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 9493 17051 9551 17057
rect 9493 17017 9505 17051
rect 9539 17048 9551 17051
rect 10042 17048 10048 17060
rect 9539 17020 10048 17048
rect 9539 17017 9551 17020
rect 9493 17011 9551 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10134 17008 10140 17060
rect 10192 17048 10198 17060
rect 10192 17020 10237 17048
rect 10192 17008 10198 17020
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6236 16952 6561 16980
rect 6236 16940 6242 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 8110 16776 8116 16788
rect 8071 16748 8116 16776
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10597 16779 10655 16785
rect 10597 16776 10609 16779
rect 10192 16748 10609 16776
rect 10192 16736 10198 16748
rect 10597 16745 10609 16748
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 7555 16711 7613 16717
rect 7555 16677 7567 16711
rect 7601 16708 7613 16711
rect 7834 16708 7840 16720
rect 7601 16680 7840 16708
rect 7601 16677 7613 16680
rect 7555 16671 7613 16677
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 9998 16711 10056 16717
rect 9998 16708 10010 16711
rect 9824 16680 10010 16708
rect 9824 16668 9830 16680
rect 9998 16677 10010 16680
rect 10044 16677 10056 16711
rect 9998 16671 10056 16677
rect 11609 16711 11667 16717
rect 11609 16677 11621 16711
rect 11655 16708 11667 16711
rect 11698 16708 11704 16720
rect 11655 16680 11704 16708
rect 11655 16677 11667 16680
rect 11609 16671 11667 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6216 16643 6274 16649
rect 6216 16640 6228 16643
rect 6144 16612 6228 16640
rect 6144 16600 6150 16612
rect 6216 16609 6228 16612
rect 6262 16609 6274 16643
rect 6216 16603 6274 16609
rect 6319 16643 6377 16649
rect 6319 16609 6331 16643
rect 6365 16640 6377 16643
rect 6822 16640 6828 16652
rect 6365 16612 6828 16640
rect 6365 16609 6377 16612
rect 6319 16603 6377 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 8220 16612 8401 16640
rect 7193 16575 7251 16581
rect 7193 16541 7205 16575
rect 7239 16572 7251 16575
rect 7282 16572 7288 16584
rect 7239 16544 7288 16572
rect 7239 16541 7251 16544
rect 7193 16535 7251 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 8220 16572 8248 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 8389 16603 8447 16609
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 7800 16544 8248 16572
rect 7800 16532 7806 16544
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11112 16544 11529 16572
rect 11112 16532 11118 16544
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 11808 16504 11836 16535
rect 10100 16476 11836 16504
rect 10100 16464 10106 16476
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 6825 16439 6883 16445
rect 6825 16436 6837 16439
rect 6696 16408 6837 16436
rect 6696 16396 6702 16408
rect 6825 16405 6837 16408
rect 6871 16405 6883 16439
rect 9398 16436 9404 16448
rect 9359 16408 9404 16436
rect 6825 16399 6883 16405
rect 9398 16396 9404 16408
rect 9456 16396 9462 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 8573 16235 8631 16241
rect 8573 16232 8585 16235
rect 8444 16204 8585 16232
rect 8444 16192 8450 16204
rect 8573 16201 8585 16204
rect 8619 16201 8631 16235
rect 11054 16232 11060 16244
rect 11015 16204 11060 16232
rect 8573 16195 8631 16201
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6236 16000 7113 16028
rect 6236 15988 6242 16000
rect 7101 15997 7113 16000
rect 7147 16028 7159 16031
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7147 16000 7481 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 7742 16028 7748 16040
rect 7699 16000 7748 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 7484 15960 7512 15991
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 8754 15988 8760 16040
rect 8812 16028 8818 16040
rect 9398 16028 9404 16040
rect 8812 16000 9404 16028
rect 8812 15988 8818 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 11146 15988 11152 16040
rect 11204 16037 11210 16040
rect 11204 16031 11242 16037
rect 11230 16028 11242 16031
rect 11609 16031 11667 16037
rect 11609 16028 11621 16031
rect 11230 16000 11621 16028
rect 11230 15997 11242 16000
rect 11204 15991 11242 15997
rect 11609 15997 11621 16000
rect 11655 15997 11667 16031
rect 11609 15991 11667 15997
rect 11204 15988 11210 15991
rect 7834 15960 7840 15972
rect 7484 15932 7840 15960
rect 7834 15920 7840 15932
rect 7892 15960 7898 15972
rect 7974 15963 8032 15969
rect 7974 15960 7986 15963
rect 7892 15932 7986 15960
rect 7892 15920 7898 15932
rect 7974 15929 7986 15932
rect 8020 15929 8032 15963
rect 7974 15923 8032 15929
rect 8941 15963 8999 15969
rect 8941 15929 8953 15963
rect 8987 15960 8999 15963
rect 9582 15960 9588 15972
rect 8987 15932 9588 15960
rect 8987 15929 8999 15932
rect 8941 15923 8999 15929
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 6181 15895 6239 15901
rect 6181 15892 6193 15895
rect 6144 15864 6193 15892
rect 6144 15852 6150 15864
rect 6181 15861 6193 15864
rect 6227 15861 6239 15895
rect 7989 15892 8017 15923
rect 9582 15920 9588 15932
rect 9640 15920 9646 15972
rect 9766 15969 9772 15972
rect 9763 15960 9772 15969
rect 9727 15932 9772 15960
rect 9763 15923 9772 15932
rect 9766 15920 9772 15923
rect 9824 15920 9830 15972
rect 10410 15920 10416 15972
rect 10468 15960 10474 15972
rect 11287 15963 11345 15969
rect 11287 15960 11299 15963
rect 10468 15932 11299 15960
rect 10468 15920 10474 15932
rect 11287 15929 11299 15932
rect 11333 15929 11345 15963
rect 11698 15960 11704 15972
rect 11287 15923 11345 15929
rect 11532 15932 11704 15960
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 7989 15864 9229 15892
rect 6181 15855 6239 15861
rect 9217 15861 9229 15864
rect 9263 15892 9275 15895
rect 9398 15892 9404 15904
rect 9263 15864 9404 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 10321 15895 10379 15901
rect 10321 15892 10333 15895
rect 9548 15864 10333 15892
rect 9548 15852 9554 15864
rect 10321 15861 10333 15864
rect 10367 15892 10379 15895
rect 11532 15892 11560 15932
rect 11698 15920 11704 15932
rect 11756 15960 11762 15972
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 11756 15932 11989 15960
rect 11756 15920 11762 15932
rect 11977 15929 11989 15932
rect 12023 15929 12035 15963
rect 11977 15923 12035 15929
rect 10367 15864 11560 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 8846 15688 8852 15700
rect 8435 15660 8852 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 9398 15648 9404 15660
rect 9456 15688 9462 15700
rect 9766 15688 9772 15700
rect 9456 15660 9772 15688
rect 9456 15648 9462 15660
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 6638 15620 6644 15632
rect 6599 15592 6644 15620
rect 6638 15580 6644 15592
rect 6696 15580 6702 15632
rect 7834 15629 7840 15632
rect 7831 15620 7840 15629
rect 7795 15592 7840 15620
rect 7831 15583 7840 15592
rect 7834 15580 7840 15583
rect 7892 15580 7898 15632
rect 9858 15620 9864 15632
rect 9819 15592 9864 15620
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 10042 15580 10048 15632
rect 10100 15620 10106 15632
rect 10413 15623 10471 15629
rect 10413 15620 10425 15623
rect 10100 15592 10425 15620
rect 10100 15580 10106 15592
rect 10413 15589 10425 15592
rect 10459 15589 10471 15623
rect 10413 15583 10471 15589
rect 5994 15552 6000 15564
rect 5955 15524 6000 15552
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15552 6515 15555
rect 6914 15552 6920 15564
rect 6503 15524 6920 15552
rect 6503 15521 6515 15524
rect 6457 15515 6515 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7558 15484 7564 15496
rect 7515 15456 7564 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 10410 15484 10416 15496
rect 9815 15456 10416 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 7282 15348 7288 15360
rect 7243 15320 7288 15348
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 5994 15144 6000 15156
rect 5955 15116 6000 15144
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7892 15116 8217 15144
rect 7892 15104 7898 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10410 15144 10416 15156
rect 10367 15116 10416 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 8110 15008 8116 15020
rect 7484 14980 8116 15008
rect 7484 14949 7512 14980
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9858 15008 9864 15020
rect 9631 14980 9864 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7147 14912 7481 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 7653 14903 7711 14909
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14940 8815 14943
rect 8941 14943 8999 14949
rect 8941 14940 8953 14943
rect 8803 14912 8953 14940
rect 8803 14909 8815 14912
rect 8757 14903 8815 14909
rect 8941 14909 8953 14912
rect 8987 14940 8999 14943
rect 9490 14940 9496 14952
rect 8987 14912 9496 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 7668 14872 7696 14903
rect 9490 14900 9496 14912
rect 9548 14900 9554 14952
rect 6932 14844 7696 14872
rect 6932 14816 6960 14844
rect 6365 14807 6423 14813
rect 6365 14773 6377 14807
rect 6411 14804 6423 14807
rect 6914 14804 6920 14816
rect 6411 14776 6920 14804
rect 6411 14773 6423 14776
rect 6365 14767 6423 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 9769 14603 9827 14609
rect 9769 14600 9781 14603
rect 9732 14572 9781 14600
rect 9732 14560 9738 14572
rect 9769 14569 9781 14572
rect 9815 14569 9827 14603
rect 9769 14563 9827 14569
rect 6178 14541 6184 14544
rect 6175 14532 6184 14541
rect 6139 14504 6184 14532
rect 6175 14495 6184 14504
rect 6178 14492 6184 14495
rect 6236 14492 6242 14544
rect 8754 14532 8760 14544
rect 8715 14504 8760 14532
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 8481 14467 8539 14473
rect 8481 14464 8493 14467
rect 8444 14436 8493 14464
rect 8444 14424 8450 14436
rect 8481 14433 8493 14436
rect 8527 14433 8539 14467
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 8481 14427 8539 14433
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 6638 14396 6644 14408
rect 5859 14368 6644 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6914 14396 6920 14408
rect 6788 14368 6920 14396
rect 6788 14356 6794 14368
rect 6914 14356 6920 14368
rect 6972 14396 6978 14408
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 6972 14368 7205 14396
rect 6972 14356 6978 14368
rect 7193 14365 7205 14368
rect 7239 14365 7251 14399
rect 8496 14396 8524 14427
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10318 14464 10324 14476
rect 10275 14436 10324 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10244 14396 10272 14427
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 8496 14368 10272 14396
rect 7193 14359 7251 14365
rect 5261 14263 5319 14269
rect 5261 14229 5273 14263
rect 5307 14260 5319 14263
rect 5350 14260 5356 14272
rect 5307 14232 5356 14260
rect 5307 14229 5319 14232
rect 5261 14223 5319 14229
rect 5350 14220 5356 14232
rect 5408 14260 5414 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 5408 14232 6745 14260
rect 5408 14220 5414 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 7558 14260 7564 14272
rect 7519 14232 7564 14260
rect 6733 14223 6791 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 7745 14059 7803 14065
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 8386 14056 8392 14068
rect 7791 14028 8392 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 9732 14028 9873 14056
rect 9732 14016 9738 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 9861 14019 9919 14025
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 7892 13960 8493 13988
rect 7892 13948 7898 13960
rect 8481 13957 8493 13960
rect 8527 13988 8539 13991
rect 8570 13988 8576 14000
rect 8527 13960 8576 13988
rect 8527 13957 8539 13960
rect 8481 13951 8539 13957
rect 8570 13948 8576 13960
rect 8628 13948 8634 14000
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5123 13892 5273 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5261 13889 5273 13892
rect 5307 13920 5319 13923
rect 5442 13920 5448 13932
rect 5307 13892 5448 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 6638 13852 6644 13864
rect 6551 13824 6644 13852
rect 6638 13812 6644 13824
rect 6696 13852 6702 13864
rect 8662 13852 8668 13864
rect 6696 13824 6868 13852
rect 8623 13824 8668 13852
rect 6696 13812 6702 13824
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5902 13784 5908 13796
rect 5408 13756 5453 13784
rect 5863 13756 5908 13784
rect 5408 13744 5414 13756
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 6840 13784 6868 13824
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 10318 13852 10324 13864
rect 10279 13824 10324 13852
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 6914 13784 6920 13796
rect 6840 13756 6920 13784
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 7101 13787 7159 13793
rect 7101 13753 7113 13787
rect 7147 13784 7159 13787
rect 7834 13784 7840 13796
rect 7147 13756 7840 13784
rect 7147 13753 7159 13756
rect 7101 13747 7159 13753
rect 7834 13744 7840 13756
rect 7892 13744 7898 13796
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 8986 13787 9044 13793
rect 8986 13784 8998 13787
rect 8628 13756 8998 13784
rect 8628 13744 8634 13756
rect 8986 13753 8998 13756
rect 9032 13753 9044 13787
rect 8986 13747 9044 13753
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 6178 13716 6184 13728
rect 5224 13688 6184 13716
rect 5224 13676 5230 13688
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 8110 13716 8116 13728
rect 8071 13688 8116 13716
rect 8110 13676 8116 13688
rect 8168 13676 8174 13728
rect 9582 13716 9588 13728
rect 9543 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 6052 13484 6469 13512
rect 6052 13472 6058 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6457 13475 6515 13481
rect 5166 13404 5172 13456
rect 5224 13453 5230 13456
rect 5224 13447 5272 13453
rect 5224 13413 5226 13447
rect 5260 13413 5272 13447
rect 5224 13407 5272 13413
rect 5224 13404 5230 13407
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 6086 13444 6092 13456
rect 5868 13416 6092 13444
rect 5868 13404 5874 13416
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 6472 13444 6500 13475
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8018 13444 8024 13456
rect 6472 13416 8024 13444
rect 6822 13376 6828 13388
rect 6783 13348 6828 13376
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7484 13385 7512 13416
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13345 7527 13379
rect 7834 13376 7840 13388
rect 7795 13348 7840 13376
rect 7469 13339 7527 13345
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4672 13280 4905 13308
rect 4672 13268 4678 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 7392 13308 7420 13339
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 7650 13308 7656 13320
rect 7392 13280 7656 13308
rect 4893 13271 4951 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9766 13308 9772 13320
rect 9723 13280 9772 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5408 13144 5825 13172
rect 5408 13132 5414 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 5813 13135 5871 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8812 13144 9137 13172
rect 8812 13132 8818 13144
rect 9125 13141 9137 13144
rect 9171 13141 9183 13175
rect 9125 13135 9183 13141
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 8389 12903 8447 12909
rect 8389 12869 8401 12903
rect 8435 12900 8447 12903
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 8435 12872 8677 12900
rect 8435 12869 8447 12872
rect 8389 12863 8447 12869
rect 8665 12869 8677 12872
rect 8711 12900 8723 12903
rect 8711 12872 9352 12900
rect 8711 12869 8723 12872
rect 8665 12863 8723 12869
rect 9324 12844 9352 12872
rect 5902 12832 5908 12844
rect 5863 12804 5908 12832
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 7374 12832 7380 12844
rect 7116 12804 7380 12832
rect 4614 12764 4620 12776
rect 4575 12736 4620 12764
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 6273 12767 6331 12773
rect 6273 12733 6285 12767
rect 6319 12764 6331 12767
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6319 12736 6653 12764
rect 6319 12733 6331 12736
rect 6273 12727 6331 12733
rect 6641 12733 6653 12736
rect 6687 12764 6699 12767
rect 6822 12764 6828 12776
rect 6687 12736 6828 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 6822 12724 6828 12736
rect 6880 12764 6886 12776
rect 7116 12773 7144 12804
rect 7374 12792 7380 12804
rect 7432 12832 7438 12844
rect 7432 12804 9076 12832
rect 7432 12792 7438 12804
rect 7101 12767 7159 12773
rect 7101 12764 7113 12767
rect 6880 12736 7113 12764
rect 6880 12724 6886 12736
rect 7101 12733 7113 12736
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 5074 12656 5080 12708
rect 5132 12696 5138 12708
rect 5261 12699 5319 12705
rect 5261 12696 5273 12699
rect 5132 12668 5273 12696
rect 5132 12656 5138 12668
rect 5261 12665 5273 12668
rect 5307 12665 5319 12699
rect 5261 12659 5319 12665
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 7576 12696 7604 12727
rect 7760 12696 7788 12727
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 9048 12773 9076 12804
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 9364 12804 10885 12832
rect 9364 12792 9370 12804
rect 8021 12767 8079 12773
rect 8021 12764 8033 12767
rect 7892 12736 8033 12764
rect 7892 12724 7898 12736
rect 8021 12733 8033 12736
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 9125 12767 9183 12773
rect 9125 12764 9137 12767
rect 9079 12736 9137 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 9125 12733 9137 12736
rect 9171 12733 9183 12767
rect 9674 12764 9680 12776
rect 9635 12736 9680 12764
rect 9125 12727 9183 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10152 12773 10180 12804
rect 10873 12801 10885 12804
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12733 10195 12767
rect 10137 12727 10195 12733
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 8110 12696 8116 12708
rect 5408 12668 5453 12696
rect 7576 12668 7696 12696
rect 7760 12668 8116 12696
rect 5408 12656 5414 12668
rect 7668 12640 7696 12668
rect 8110 12656 8116 12668
rect 8168 12696 8174 12708
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 8168 12668 8401 12696
rect 8168 12656 8174 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 8389 12659 8447 12665
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 10336 12696 10364 12727
rect 8812 12668 10364 12696
rect 8812 12656 8818 12668
rect 4985 12631 5043 12637
rect 4985 12597 4997 12631
rect 5031 12628 5043 12631
rect 5166 12628 5172 12640
rect 5031 12600 5172 12628
rect 5031 12597 5043 12600
rect 4985 12591 5043 12597
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 6914 12628 6920 12640
rect 6875 12600 6920 12628
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7650 12588 7656 12640
rect 7708 12588 7714 12640
rect 9398 12628 9404 12640
rect 9359 12600 9404 12628
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 5261 12427 5319 12433
rect 5261 12393 5273 12427
rect 5307 12424 5319 12427
rect 5350 12424 5356 12436
rect 5307 12396 5356 12424
rect 5307 12393 5319 12396
rect 5261 12387 5319 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 5537 12427 5595 12433
rect 5537 12424 5549 12427
rect 5500 12396 5549 12424
rect 5500 12384 5506 12396
rect 5537 12393 5549 12396
rect 5583 12393 5595 12427
rect 8662 12424 8668 12436
rect 8623 12396 8668 12424
rect 5537 12387 5595 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9582 12384 9588 12436
rect 9640 12384 9646 12436
rect 6549 12359 6607 12365
rect 6549 12325 6561 12359
rect 6595 12356 6607 12359
rect 6917 12359 6975 12365
rect 6917 12356 6929 12359
rect 6595 12328 6929 12356
rect 6595 12325 6607 12328
rect 6549 12319 6607 12325
rect 6917 12325 6929 12328
rect 6963 12356 6975 12359
rect 7650 12356 7656 12368
rect 6963 12328 7656 12356
rect 6963 12325 6975 12328
rect 6917 12319 6975 12325
rect 7650 12316 7656 12328
rect 7708 12356 7714 12368
rect 9600 12356 9628 12384
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 7708 12328 9260 12356
rect 9600 12328 9873 12356
rect 7708 12316 7714 12328
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7944 12297 7972 12328
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 7929 12251 7987 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8662 12288 8668 12300
rect 8623 12260 8668 12288
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 9232 12297 9260 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9582 12288 9588 12300
rect 9263 12260 9588 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10870 12220 10876 12232
rect 10459 12192 10876 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12084 4951 12087
rect 5074 12084 5080 12096
rect 4939 12056 5080 12084
rect 4939 12053 4951 12056
rect 4893 12047 4951 12053
rect 5074 12044 5080 12056
rect 5132 12084 5138 12096
rect 5442 12084 5448 12096
rect 5132 12056 5448 12084
rect 5132 12044 5138 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 6052 12056 6101 12084
rect 6052 12044 6058 12056
rect 6089 12053 6101 12056
rect 6135 12084 6147 12087
rect 7834 12084 7840 12096
rect 6135 12056 7840 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10652 12056 10701 12084
rect 10652 12044 10658 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 7432 11852 7941 11880
rect 7432 11840 7438 11852
rect 7929 11849 7941 11852
rect 7975 11849 7987 11883
rect 8570 11880 8576 11892
rect 8531 11852 8576 11880
rect 7929 11843 7987 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9824 11852 9965 11880
rect 9824 11840 9830 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 7650 11744 7656 11756
rect 7611 11716 7656 11744
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 9030 11744 9036 11756
rect 8803 11716 9036 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 9030 11704 9036 11716
rect 9088 11744 9094 11756
rect 9398 11744 9404 11756
rect 9088 11716 9404 11744
rect 9088 11704 9094 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 10870 11744 10876 11756
rect 10831 11716 10876 11744
rect 10870 11704 10876 11716
rect 10928 11744 10934 11756
rect 11974 11744 11980 11756
rect 10928 11716 11980 11744
rect 10928 11704 10934 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 7374 11676 7380 11688
rect 6687 11648 7380 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 9078 11611 9136 11617
rect 9078 11608 9090 11611
rect 8628 11580 9090 11608
rect 8628 11568 8634 11580
rect 9078 11577 9090 11580
rect 9124 11577 9136 11611
rect 10594 11608 10600 11620
rect 10555 11580 10600 11608
rect 9078 11571 9136 11577
rect 10594 11568 10600 11580
rect 10652 11568 10658 11620
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11577 10747 11611
rect 10689 11571 10747 11577
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9723 11512 10333 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 10321 11509 10333 11512
rect 10367 11540 10379 11543
rect 10704 11540 10732 11571
rect 10367 11512 10732 11540
rect 10367 11509 10379 11512
rect 10321 11503 10379 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 7377 11339 7435 11345
rect 7377 11305 7389 11339
rect 7423 11336 7435 11339
rect 7650 11336 7656 11348
rect 7423 11308 7656 11336
rect 7423 11305 7435 11308
rect 7377 11299 7435 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 9030 11336 9036 11348
rect 8991 11308 9036 11336
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9490 11336 9496 11348
rect 9451 11308 9496 11336
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9824 11240 9873 11268
rect 9824 11228 9830 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 8110 11160 8116 11212
rect 8168 11209 8174 11212
rect 8168 11203 8206 11209
rect 8194 11169 8206 11203
rect 8168 11163 8206 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10594 11200 10600 11212
rect 10459 11172 10600 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 8168 11160 8174 11163
rect 10594 11160 10600 11172
rect 10652 11200 10658 11212
rect 10870 11200 10876 11212
rect 10652 11172 10876 11200
rect 10652 11160 10658 11172
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11276 11203 11334 11209
rect 11276 11200 11288 11203
rect 11112 11172 11288 11200
rect 11112 11160 11118 11172
rect 11276 11169 11288 11172
rect 11322 11169 11334 11203
rect 11276 11163 11334 11169
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 10962 11132 10968 11144
rect 9815 11104 10968 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 10410 11024 10416 11076
rect 10468 11064 10474 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 10468 11036 10793 11064
rect 10468 11024 10474 11036
rect 10781 11033 10793 11036
rect 10827 11064 10839 11067
rect 11379 11067 11437 11073
rect 11379 11064 11391 11067
rect 10827 11036 11391 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11379 11033 11391 11036
rect 11425 11033 11437 11067
rect 11379 11027 11437 11033
rect 7009 10999 7067 11005
rect 7009 10965 7021 10999
rect 7055 10996 7067 10999
rect 7098 10996 7104 11008
rect 7055 10968 7104 10996
rect 7055 10965 7067 10968
rect 7009 10959 7067 10965
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7745 10999 7803 11005
rect 7745 10965 7757 10999
rect 7791 10996 7803 10999
rect 8018 10996 8024 11008
rect 7791 10968 8024 10996
rect 7791 10965 7803 10968
rect 7745 10959 7803 10965
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 8202 10956 8208 11008
rect 8260 11005 8266 11008
rect 8260 10999 8309 11005
rect 8260 10965 8263 10999
rect 8297 10965 8309 10999
rect 8570 10996 8576 11008
rect 8531 10968 8576 10996
rect 8260 10959 8309 10965
rect 8260 10956 8266 10959
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 11112 10764 11253 10792
rect 11112 10752 11118 10764
rect 11241 10761 11253 10764
rect 11287 10792 11299 10795
rect 12710 10792 12716 10804
rect 11287 10764 12716 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 8110 10724 8116 10736
rect 8071 10696 8116 10724
rect 8110 10684 8116 10696
rect 8168 10684 8174 10736
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10410 10656 10416 10668
rect 10275 10628 10416 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 8389 10591 8447 10597
rect 6871 10560 7420 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 7392 10464 7420 10560
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8570 10588 8576 10600
rect 8435 10560 8576 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8570 10548 8576 10560
rect 8628 10588 8634 10600
rect 9398 10588 9404 10600
rect 8628 10560 9404 10588
rect 8628 10548 8634 10560
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 8710 10523 8768 10529
rect 8710 10520 8722 10523
rect 7883 10492 8722 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8710 10489 8722 10492
rect 8756 10520 8768 10523
rect 8846 10520 8852 10532
rect 8756 10492 8852 10520
rect 8756 10489 8768 10492
rect 8710 10483 8768 10489
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 10321 10523 10379 10529
rect 9324 10492 9904 10520
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 7006 10452 7012 10464
rect 6967 10424 7012 10452
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 9324 10461 9352 10492
rect 9876 10464 9904 10492
rect 10321 10489 10333 10523
rect 10367 10489 10379 10523
rect 10870 10520 10876 10532
rect 10831 10492 10876 10520
rect 10321 10483 10379 10489
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10421 9367 10455
rect 9309 10415 9367 10421
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9766 10452 9772 10464
rect 9723 10424 9772 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 9953 10455 10011 10461
rect 9953 10452 9965 10455
rect 9916 10424 9965 10452
rect 9916 10412 9922 10424
rect 9953 10421 9965 10424
rect 9999 10452 10011 10455
rect 10336 10452 10364 10483
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 9999 10424 10364 10452
rect 9999 10421 10011 10424
rect 9953 10415 10011 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 5445 10183 5503 10189
rect 5445 10180 5457 10183
rect 5408 10152 5457 10180
rect 5408 10140 5414 10152
rect 5445 10149 5457 10152
rect 5491 10149 5503 10183
rect 5445 10143 5503 10149
rect 8846 10140 8852 10192
rect 8904 10180 8910 10192
rect 9998 10183 10056 10189
rect 9998 10180 10010 10183
rect 8904 10152 10010 10180
rect 8904 10140 8910 10152
rect 9998 10149 10010 10152
rect 10044 10149 10056 10183
rect 9998 10143 10056 10149
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 11609 10183 11667 10189
rect 11609 10180 11621 10183
rect 11572 10152 11621 10180
rect 11572 10140 11578 10152
rect 11609 10149 11621 10152
rect 11655 10149 11667 10183
rect 11609 10143 11667 10149
rect 7466 10112 7472 10124
rect 7427 10084 7472 10112
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10081 7803 10115
rect 8110 10112 8116 10124
rect 8071 10084 8116 10112
rect 7745 10075 7803 10081
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 4724 10016 5365 10044
rect 4724 9920 4752 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5353 10007 5411 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 7760 10044 7788 10075
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8662 10112 8668 10124
rect 8527 10084 8668 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 8496 10044 8524 10075
rect 8662 10072 8668 10084
rect 8720 10112 8726 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8720 10084 9137 10112
rect 8720 10072 8726 10084
rect 9125 10081 9137 10084
rect 9171 10112 9183 10115
rect 9582 10112 9588 10124
rect 9171 10084 9588 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 7024 10016 7788 10044
rect 7852 10016 8524 10044
rect 8757 10047 8815 10053
rect 7024 9920 7052 10016
rect 7852 9920 7880 10016
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 8803 10016 9689 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9677 10013 9689 10016
rect 9723 10044 9735 10047
rect 11054 10044 11060 10056
rect 9723 10016 11060 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11974 10044 11980 10056
rect 11935 10016 11980 10044
rect 11517 10007 11575 10013
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 10597 9979 10655 9985
rect 10597 9976 10609 9979
rect 9824 9948 10609 9976
rect 9824 9936 9830 9948
rect 10597 9945 10609 9948
rect 10643 9976 10655 9979
rect 11146 9976 11152 9988
rect 10643 9948 11152 9976
rect 10643 9945 10655 9948
rect 10597 9939 10655 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11532 9976 11560 10007
rect 11974 10004 11980 10016
rect 12032 10044 12038 10056
rect 12618 10044 12624 10056
rect 12032 10016 12624 10044
rect 12032 10004 12038 10016
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 11882 9976 11888 9988
rect 11532 9948 11888 9976
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5350 9908 5356 9920
rect 5215 9880 5356 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 6457 9911 6515 9917
rect 6457 9877 6469 9911
rect 6503 9908 6515 9911
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6503 9880 6837 9908
rect 6503 9877 6515 9880
rect 6457 9871 6515 9877
rect 6825 9877 6837 9880
rect 6871 9908 6883 9911
rect 7006 9908 7012 9920
rect 6871 9880 7012 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 7156 9880 7205 9908
rect 7156 9868 7162 9880
rect 7193 9877 7205 9880
rect 7239 9908 7251 9911
rect 7834 9908 7840 9920
rect 7239 9880 7840 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 10962 9908 10968 9920
rect 10923 9880 10968 9908
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 12618 9704 12624 9716
rect 7524 9676 8248 9704
rect 7524 9664 7530 9676
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5810 9636 5816 9648
rect 5500 9608 5816 9636
rect 5500 9596 5506 9608
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 8220 9636 8248 9676
rect 12452 9676 12624 9704
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8220 9608 8585 9636
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8573 9599 8631 9605
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4223 9540 4721 9568
rect 4223 9509 4251 9540
rect 4709 9537 4721 9540
rect 4755 9568 4767 9571
rect 4798 9568 4804 9580
rect 4755 9540 4804 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 8202 9568 8208 9580
rect 6687 9540 8208 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 4208 9503 4266 9509
rect 4208 9469 4220 9503
rect 4254 9469 4266 9503
rect 4208 9463 4266 9469
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9500 6331 9503
rect 7098 9500 7104 9512
rect 6319 9472 7104 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7668 9509 7696 9540
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 8018 9500 8024 9512
rect 7699 9472 7733 9500
rect 7979 9472 8024 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 4065 9435 4123 9441
rect 4065 9401 4077 9435
rect 4111 9432 4123 9435
rect 4295 9435 4353 9441
rect 4295 9432 4307 9435
rect 4111 9404 4307 9432
rect 4111 9401 4123 9404
rect 4065 9395 4123 9401
rect 4295 9401 4307 9404
rect 4341 9432 4353 9435
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4341 9404 5273 9432
rect 4341 9401 4353 9404
rect 4295 9395 4353 9401
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5261 9395 5319 9401
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 5534 9432 5540 9444
rect 5408 9404 5540 9432
rect 5408 9392 5414 9404
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7576 9432 7604 9463
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8588 9500 8616 9599
rect 11054 9596 11060 9648
rect 11112 9636 11118 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 11112 9608 11253 9636
rect 11112 9596 11118 9608
rect 11241 9605 11253 9608
rect 11287 9605 11299 9639
rect 11241 9599 11299 9605
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 9364 9540 10885 9568
rect 9364 9528 9370 9540
rect 9122 9500 9128 9512
rect 8588 9472 9128 9500
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 9968 9509 9996 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 12452 9568 12480 9676
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 12452 9540 13308 9568
rect 10873 9531 10931 9537
rect 9585 9503 9643 9509
rect 9585 9500 9597 9503
rect 9548 9472 9597 9500
rect 9548 9460 9554 9472
rect 9585 9469 9597 9472
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 8386 9432 8392 9444
rect 7064 9404 8392 9432
rect 7064 9392 7070 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 10336 9432 10364 9463
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 12434 9500 12440 9512
rect 12492 9509 12498 9512
rect 12492 9503 12530 9509
rect 11480 9472 12440 9500
rect 11480 9460 11486 9472
rect 12434 9460 12440 9472
rect 12518 9500 12530 9503
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12518 9472 12909 9500
rect 12518 9469 12530 9472
rect 12492 9463 12530 9469
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 13280 9500 13308 9540
rect 13484 9503 13542 9509
rect 13484 9500 13496 9503
rect 13280 9472 13496 9500
rect 12897 9463 12955 9469
rect 13484 9469 13496 9472
rect 13530 9500 13542 9503
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13530 9472 13921 9500
rect 13530 9469 13542 9472
rect 13484 9463 13542 9469
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 12492 9460 12498 9463
rect 10686 9432 10692 9444
rect 9732 9404 10692 9432
rect 9732 9392 9738 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 12575 9435 12633 9441
rect 12575 9432 12587 9435
rect 11020 9404 12587 9432
rect 11020 9392 11026 9404
rect 12575 9401 12587 9404
rect 12621 9401 12633 9435
rect 12575 9395 12633 9401
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5994 9364 6000 9376
rect 5123 9336 6000 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 8904 9336 8953 9364
rect 8904 9324 8910 9336
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 9398 9364 9404 9376
rect 9359 9336 9404 9364
rect 8941 9327 8999 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11572 9336 11621 9364
rect 11572 9324 11578 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11974 9364 11980 9376
rect 11935 9336 11980 9364
rect 11609 9327 11667 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 13630 9373 13636 9376
rect 13587 9367 13636 9373
rect 13587 9333 13599 9367
rect 13633 9333 13636 9367
rect 13587 9327 13636 9333
rect 13630 9324 13636 9327
rect 13688 9324 13694 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 6638 9160 6644 9172
rect 6599 9132 6644 9160
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 4979 9095 5037 9101
rect 4979 9061 4991 9095
rect 5025 9092 5037 9095
rect 5074 9092 5080 9104
rect 5025 9064 5080 9092
rect 5025 9061 5037 9064
rect 4979 9055 5037 9061
rect 5074 9052 5080 9064
rect 5132 9052 5138 9104
rect 6273 9095 6331 9101
rect 6273 9061 6285 9095
rect 6319 9092 6331 9095
rect 6319 9064 7052 9092
rect 6319 9061 6331 9064
rect 6273 9055 6331 9061
rect 7024 9036 7052 9064
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 9548 9064 10180 9092
rect 9548 9052 9554 9064
rect 4614 9024 4620 9036
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 8993 6699 9027
rect 7006 9024 7012 9036
rect 6967 8996 7012 9024
rect 6641 8987 6699 8993
rect 6656 8956 6684 8987
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7190 9024 7196 9036
rect 7151 8996 7196 9024
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 9024 7803 9027
rect 8018 9024 8024 9036
rect 7791 8996 8024 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 7098 8956 7104 8968
rect 6656 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7650 8956 7656 8968
rect 7156 8928 7656 8956
rect 7156 8916 7162 8928
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 5905 8823 5963 8829
rect 5905 8789 5917 8823
rect 5951 8820 5963 8823
rect 5994 8820 6000 8832
rect 5951 8792 6000 8820
rect 5951 8789 5963 8792
rect 5905 8783 5963 8789
rect 5994 8780 6000 8792
rect 6052 8820 6058 8832
rect 7760 8820 7788 8987
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10042 9024 10048 9036
rect 9999 8996 10048 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10152 9033 10180 9064
rect 11146 9052 11152 9104
rect 11204 9092 11210 9104
rect 12158 9092 12164 9104
rect 11204 9064 12164 9092
rect 11204 9052 11210 9064
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 8993 10195 9027
rect 10137 8987 10195 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10520 8956 10548 8987
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10744 8996 10885 9024
rect 10744 8984 10750 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 13538 8984 13544 9036
rect 13596 9033 13602 9036
rect 13596 9027 13634 9033
rect 13622 8993 13634 9027
rect 13596 8987 13634 8993
rect 13596 8984 13602 8987
rect 12066 8956 12072 8968
rect 9732 8928 10548 8956
rect 12027 8928 12072 8956
rect 9732 8916 9738 8928
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 11974 8888 11980 8900
rect 11204 8860 11980 8888
rect 11204 8848 11210 8860
rect 11974 8848 11980 8860
rect 12032 8888 12038 8900
rect 12360 8888 12388 8919
rect 12032 8860 12388 8888
rect 12032 8848 12038 8860
rect 8110 8820 8116 8832
rect 6052 8792 7788 8820
rect 8071 8792 8116 8820
rect 6052 8780 6058 8792
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8757 8823 8815 8829
rect 8757 8820 8769 8823
rect 8444 8792 8769 8820
rect 8444 8780 8450 8792
rect 8757 8789 8769 8792
rect 8803 8820 8815 8823
rect 9490 8820 9496 8832
rect 8803 8792 9496 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 13679 8823 13737 8829
rect 13679 8820 13691 8823
rect 12400 8792 13691 8820
rect 12400 8780 12406 8792
rect 13679 8789 13691 8792
rect 13725 8789 13737 8823
rect 13679 8783 13737 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4295 8619 4353 8625
rect 4295 8585 4307 8619
rect 4341 8616 4353 8619
rect 4706 8616 4712 8628
rect 4341 8588 4712 8616
rect 4341 8585 4353 8588
rect 4295 8579 4353 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 7190 8616 7196 8628
rect 6503 8588 7196 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 8168 8588 9137 8616
rect 8168 8576 8174 8588
rect 9125 8585 9137 8588
rect 9171 8616 9183 8619
rect 9674 8616 9680 8628
rect 9171 8588 9680 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 10100 8588 11253 8616
rect 10100 8576 10106 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11241 8579 11299 8585
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12158 8616 12164 8628
rect 12115 8588 12164 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 6730 8548 6736 8560
rect 6236 8520 6736 8548
rect 6236 8508 6242 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 7285 8551 7343 8557
rect 7285 8517 7297 8551
rect 7331 8548 7343 8551
rect 7834 8548 7840 8560
rect 7331 8520 7840 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 7834 8508 7840 8520
rect 7892 8548 7898 8560
rect 8570 8548 8576 8560
rect 7892 8520 8576 8548
rect 7892 8508 7898 8520
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10686 8508 10692 8560
rect 10744 8548 10750 8560
rect 10873 8551 10931 8557
rect 10873 8548 10885 8551
rect 10744 8520 10885 8548
rect 10744 8508 10750 8520
rect 10873 8517 10885 8520
rect 10919 8517 10931 8551
rect 10873 8511 10931 8517
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 13538 8548 13544 8560
rect 11940 8520 13544 8548
rect 11940 8508 11946 8520
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5626 8480 5632 8492
rect 5307 8452 5632 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5902 8480 5908 8492
rect 5863 8452 5908 8480
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 8662 8480 8668 8492
rect 8312 8452 8668 8480
rect 4208 8415 4266 8421
rect 4208 8381 4220 8415
rect 4254 8412 4266 8415
rect 4254 8381 4267 8412
rect 4208 8375 4267 8381
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 4239 8276 4267 8375
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5920 8344 5948 8440
rect 7650 8412 7656 8424
rect 7611 8384 7656 8412
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 8312 8421 8340 8452
rect 8662 8440 8668 8452
rect 8720 8480 8726 8492
rect 9306 8480 9312 8492
rect 8720 8452 9312 8480
rect 8720 8440 8726 8452
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 8113 8375 8171 8381
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8381 8355 8415
rect 8570 8412 8576 8424
rect 8531 8384 8576 8412
rect 8297 8375 8355 8381
rect 5408 8316 5453 8344
rect 5552 8316 5948 8344
rect 8128 8344 8156 8375
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 8904 8384 9505 8412
rect 8904 8372 8910 8384
rect 9493 8381 9505 8384
rect 9539 8381 9551 8415
rect 9674 8412 9680 8424
rect 9635 8384 9680 8412
rect 9493 8375 9551 8381
rect 8386 8344 8392 8356
rect 8128 8316 8392 8344
rect 5408 8304 5414 8316
rect 4617 8279 4675 8285
rect 4617 8276 4629 8279
rect 1544 8248 4629 8276
rect 1544 8236 1550 8248
rect 4617 8245 4629 8248
rect 4663 8276 4675 8279
rect 4798 8276 4804 8288
rect 4663 8248 4804 8276
rect 4663 8245 4675 8248
rect 4617 8239 4675 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 5074 8276 5080 8288
rect 5035 8248 5080 8276
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5552 8276 5580 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 9508 8344 9536 8375
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 12434 8372 12440 8424
rect 12492 8421 12498 8424
rect 12492 8415 12530 8421
rect 12518 8412 12530 8415
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12518 8384 12909 8412
rect 12518 8381 12530 8384
rect 12492 8375 12530 8381
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12492 8372 12498 8375
rect 9998 8347 10056 8353
rect 9998 8344 10010 8347
rect 9508 8316 10010 8344
rect 9998 8313 10010 8316
rect 10044 8313 10056 8347
rect 9998 8307 10056 8313
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11609 8347 11667 8353
rect 11609 8344 11621 8347
rect 11112 8316 11621 8344
rect 11112 8304 11118 8316
rect 11609 8313 11621 8316
rect 11655 8344 11667 8347
rect 12066 8344 12072 8356
rect 11655 8316 12072 8344
rect 11655 8313 11667 8316
rect 11609 8307 11667 8313
rect 12066 8304 12072 8316
rect 12124 8304 12130 8356
rect 12618 8353 12624 8356
rect 12575 8347 12624 8353
rect 12575 8313 12587 8347
rect 12621 8313 12624 8347
rect 12575 8307 12624 8313
rect 12618 8304 12624 8307
rect 12676 8304 12682 8356
rect 8754 8276 8760 8288
rect 5500 8248 5580 8276
rect 8715 8248 8760 8276
rect 5500 8236 5506 8248
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 10594 8276 10600 8288
rect 10555 8248 10600 8276
rect 10594 8236 10600 8248
rect 10652 8236 10658 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 4614 8072 4620 8084
rect 4575 8044 4620 8072
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7524 8044 7665 8072
rect 7524 8032 7530 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8662 8072 8668 8084
rect 8067 8044 8668 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8812 8044 9045 8072
rect 8812 8032 8818 8044
rect 9033 8041 9045 8044
rect 9079 8072 9091 8075
rect 9674 8072 9680 8084
rect 9079 8044 9680 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 5718 8004 5724 8016
rect 5132 7976 5724 8004
rect 5132 7964 5138 7976
rect 5718 7964 5724 7976
rect 5776 8004 5782 8016
rect 6042 8007 6100 8013
rect 6042 8004 6054 8007
rect 5776 7976 6054 8004
rect 5776 7964 5782 7976
rect 6042 7973 6054 7976
rect 6088 7973 6100 8007
rect 8386 8004 8392 8016
rect 8299 7976 8392 8004
rect 6042 7967 6100 7973
rect 8386 7964 8392 7976
rect 8444 8004 8450 8016
rect 9401 8007 9459 8013
rect 9401 8004 9413 8007
rect 8444 7976 9413 8004
rect 8444 7964 8450 7976
rect 9401 7973 9413 7976
rect 9447 7973 9459 8007
rect 9858 8004 9864 8016
rect 9819 7976 9864 8004
rect 9401 7967 9459 7973
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 11425 8007 11483 8013
rect 11425 8004 11437 8007
rect 10652 7976 11437 8004
rect 10652 7964 10658 7976
rect 11425 7973 11437 7976
rect 11471 7973 11483 8007
rect 11425 7967 11483 7973
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5350 7936 5356 7948
rect 5307 7908 5356 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 5408 7908 6653 7936
rect 5408 7896 5414 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 6641 7899 6699 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 8352 7908 8493 7936
rect 8352 7896 8358 7908
rect 8481 7905 8493 7908
rect 8527 7905 8539 7939
rect 8481 7899 8539 7905
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7377 7871 7435 7877
rect 7377 7868 7389 7871
rect 7055 7840 7389 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7377 7837 7389 7840
rect 7423 7868 7435 7871
rect 7650 7868 7656 7880
rect 7423 7840 7656 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 5736 7800 5764 7831
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 9950 7868 9956 7880
rect 9815 7840 9956 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 10778 7868 10784 7880
rect 10459 7840 10784 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 10778 7828 10784 7840
rect 10836 7868 10842 7880
rect 11146 7868 11152 7880
rect 10836 7840 11152 7868
rect 10836 7828 10842 7840
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 12342 7868 12348 7880
rect 11379 7840 12348 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 6638 7800 6644 7812
rect 5736 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 10928 7772 11897 7800
rect 10928 7760 10934 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 5626 7732 5632 7744
rect 5539 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7732 5690 7744
rect 5902 7732 5908 7744
rect 5684 7704 5908 7732
rect 5684 7692 5690 7704
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6638 7528 6644 7540
rect 6227 7500 6644 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12342 7528 12348 7540
rect 11931 7500 12348 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 7650 7392 7656 7404
rect 7607 7364 7656 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 10502 7392 10508 7404
rect 10463 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 10778 7392 10784 7404
rect 10739 7364 10784 7392
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 8662 7324 8668 7336
rect 8623 7296 8668 7324
rect 6917 7287 6975 7293
rect 6932 7256 6960 7287
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 7466 7256 7472 7268
rect 6932 7228 7472 7256
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 5718 7188 5724 7200
rect 5408 7160 5724 7188
rect 5408 7148 5414 7160
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6638 7188 6644 7200
rect 6599 7160 6644 7188
rect 6638 7148 6644 7160
rect 6696 7188 6702 7200
rect 6932 7188 6960 7228
rect 7466 7216 7472 7228
rect 7524 7256 7530 7268
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7524 7228 7849 7256
rect 7524 7216 7530 7228
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 8986 7259 9044 7265
rect 8986 7256 8998 7259
rect 8904 7228 8998 7256
rect 8904 7216 8910 7228
rect 8986 7225 8998 7228
rect 9032 7225 9044 7259
rect 8986 7219 9044 7225
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 10652 7228 10697 7256
rect 10652 7216 10658 7228
rect 6696 7160 6960 7188
rect 6696 7148 6702 7160
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8352 7160 8493 7188
rect 8352 7148 8358 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 10612 7188 10640 7216
rect 11425 7191 11483 7197
rect 11425 7188 11437 7191
rect 10367 7160 11437 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 11425 7157 11437 7160
rect 11471 7157 11483 7191
rect 11425 7151 11483 7157
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 8720 6956 9137 6984
rect 8720 6944 8726 6956
rect 9125 6953 9137 6956
rect 9171 6984 9183 6987
rect 9582 6984 9588 6996
rect 9171 6956 9588 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10137 6987 10195 6993
rect 10137 6984 10149 6987
rect 10008 6956 10149 6984
rect 10008 6944 10014 6956
rect 10137 6953 10149 6956
rect 10183 6953 10195 6987
rect 10502 6984 10508 6996
rect 10463 6956 10508 6984
rect 10137 6947 10195 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4960 6851 5018 6857
rect 4960 6848 4972 6851
rect 4396 6820 4972 6848
rect 4396 6808 4402 6820
rect 4960 6817 4972 6820
rect 5006 6848 5018 6851
rect 5442 6848 5448 6860
rect 5006 6820 5448 6848
rect 5006 6817 5018 6820
rect 4960 6811 5018 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 7285 6851 7343 6857
rect 7285 6848 7297 6851
rect 7248 6820 7297 6848
rect 7248 6808 7254 6820
rect 7285 6817 7297 6820
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 9674 6808 9680 6860
rect 9732 6857 9738 6860
rect 9732 6851 9770 6857
rect 9758 6817 9770 6851
rect 9732 6811 9770 6817
rect 9815 6851 9873 6857
rect 9815 6817 9827 6851
rect 9861 6848 9873 6851
rect 10962 6848 10968 6860
rect 9861 6820 10968 6848
rect 9861 6817 9873 6820
rect 9815 6811 9873 6817
rect 9732 6808 9738 6811
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 5031 6715 5089 6721
rect 5031 6712 5043 6715
rect 3936 6684 5043 6712
rect 3936 6672 3942 6684
rect 5031 6681 5043 6684
rect 5077 6681 5089 6715
rect 5031 6675 5089 6681
rect 7469 6715 7527 6721
rect 7469 6681 7481 6715
rect 7515 6712 7527 6715
rect 8110 6712 8116 6724
rect 7515 6684 8116 6712
rect 7515 6681 7527 6684
rect 7469 6675 7527 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 8665 6647 8723 6653
rect 8665 6644 8677 6647
rect 8536 6616 8677 6644
rect 8536 6604 8542 6616
rect 8665 6613 8677 6616
rect 8711 6644 8723 6647
rect 8846 6644 8852 6656
rect 8711 6616 8852 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 4338 6440 4344 6452
rect 4299 6412 4344 6440
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 7190 6440 7196 6452
rect 7151 6412 7196 6440
rect 7190 6400 7196 6412
rect 7248 6440 7254 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7248 6412 7941 6440
rect 7248 6400 7254 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8665 6443 8723 6449
rect 8665 6440 8677 6443
rect 8628 6412 8677 6440
rect 8628 6400 8634 6412
rect 8665 6409 8677 6412
rect 8711 6409 8723 6443
rect 8665 6403 8723 6409
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6564 6208 7021 6236
rect 4706 6168 4712 6180
rect 4619 6140 4712 6168
rect 4706 6128 4712 6140
rect 4764 6168 4770 6180
rect 5261 6171 5319 6177
rect 5261 6168 5273 6171
rect 4764 6140 5273 6168
rect 4764 6128 4770 6140
rect 5261 6137 5273 6140
rect 5307 6137 5319 6171
rect 5261 6131 5319 6137
rect 5353 6171 5411 6177
rect 5353 6137 5365 6171
rect 5399 6168 5411 6171
rect 5442 6168 5448 6180
rect 5399 6140 5448 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5368 6100 5396 6131
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5902 6168 5908 6180
rect 5863 6140 5908 6168
rect 5902 6128 5908 6140
rect 5960 6128 5966 6180
rect 5123 6072 5396 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 6564 6109 6592 6208
rect 7009 6205 7021 6208
rect 7055 6236 7067 6239
rect 8294 6236 8300 6248
rect 7055 6208 8300 6236
rect 7055 6205 7067 6208
rect 7009 6199 7067 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8527 6208 9076 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 9048 6109 9076 6208
rect 9674 6168 9680 6180
rect 9635 6140 9680 6168
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 6549 6103 6607 6109
rect 6549 6100 6561 6103
rect 6236 6072 6561 6100
rect 6236 6060 6242 6072
rect 6549 6069 6561 6072
rect 6595 6069 6607 6103
rect 6549 6063 6607 6069
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9306 6100 9312 6112
rect 9079 6072 9312 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 4387 5899 4445 5905
rect 4387 5865 4399 5899
rect 4433 5896 4445 5899
rect 4706 5896 4712 5908
rect 4433 5868 4712 5896
rect 4433 5865 4445 5868
rect 4387 5859 4445 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7190 5896 7196 5908
rect 6963 5868 7196 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 7558 5896 7564 5908
rect 7331 5868 7564 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 5169 5831 5227 5837
rect 5169 5797 5181 5831
rect 5215 5828 5227 5831
rect 5442 5828 5448 5840
rect 5215 5800 5448 5828
rect 5215 5797 5227 5800
rect 5169 5791 5227 5797
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 7208 5828 7236 5856
rect 7650 5828 7656 5840
rect 7208 5800 7656 5828
rect 7650 5788 7656 5800
rect 7708 5828 7714 5840
rect 7708 5800 8248 5828
rect 7708 5788 7714 5800
rect 4246 5720 4252 5772
rect 4304 5769 4310 5772
rect 4304 5763 4342 5769
rect 4330 5729 4342 5763
rect 4304 5723 4342 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7282 5760 7288 5772
rect 6595 5732 7288 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 4304 5720 4310 5723
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7558 5760 7564 5772
rect 7519 5732 7564 5760
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7834 5760 7840 5772
rect 7795 5732 7840 5760
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8220 5769 8248 5800
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 4120 5664 5365 5692
rect 4120 5652 4126 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5810 5692 5816 5704
rect 5771 5664 5816 5692
rect 5353 5655 5411 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 3099 5355 3157 5361
rect 3099 5321 3111 5355
rect 3145 5352 3157 5355
rect 3881 5355 3939 5361
rect 3881 5352 3893 5355
rect 3145 5324 3893 5352
rect 3145 5321 3157 5324
rect 3099 5315 3157 5321
rect 3881 5321 3893 5324
rect 3927 5352 3939 5355
rect 4062 5352 4068 5364
rect 3927 5324 4068 5352
rect 3927 5321 3939 5324
rect 3881 5315 3939 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4304 5324 4445 5352
rect 4304 5312 4310 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5905 5355 5963 5361
rect 5905 5352 5917 5355
rect 5592 5324 5917 5352
rect 5592 5312 5598 5324
rect 5905 5321 5917 5324
rect 5951 5321 5963 5355
rect 5905 5315 5963 5321
rect 3510 5284 3516 5296
rect 3471 5256 3516 5284
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 9953 5287 10011 5293
rect 9953 5253 9965 5287
rect 9999 5284 10011 5287
rect 11330 5284 11336 5296
rect 9999 5256 11336 5284
rect 9999 5253 10011 5256
rect 9953 5247 10011 5253
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 3028 5151 3086 5157
rect 3028 5117 3040 5151
rect 3074 5148 3086 5151
rect 3528 5148 3556 5244
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 7668 5188 8585 5216
rect 7668 5160 7696 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 3074 5120 3556 5148
rect 4024 5151 4082 5157
rect 3074 5117 3086 5120
rect 3028 5111 3086 5117
rect 4024 5117 4036 5151
rect 4070 5148 4082 5151
rect 4070 5117 4108 5148
rect 4024 5111 4108 5117
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 4080 5080 4108 5111
rect 4798 5108 4804 5160
rect 4856 5148 4862 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4856 5120 4997 5148
rect 4856 5108 4862 5120
rect 4985 5117 4997 5120
rect 5031 5148 5043 5151
rect 6638 5148 6644 5160
rect 5031 5120 5488 5148
rect 6551 5120 6644 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5350 5089 5356 5092
rect 5347 5080 5356 5089
rect 3936 5052 4936 5080
rect 5311 5052 5356 5080
rect 3936 5040 3942 5052
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4908 5021 4936 5052
rect 5347 5043 5356 5052
rect 5350 5040 5356 5043
rect 5408 5040 5414 5092
rect 5460 5080 5488 5120
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 7006 5148 7012 5160
rect 6696 5120 7012 5148
rect 6696 5108 6702 5120
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7374 5148 7380 5160
rect 7335 5120 7380 5148
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7650 5148 7656 5160
rect 7611 5120 7656 5148
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8202 5148 8208 5160
rect 8163 5120 8208 5148
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 9766 5148 9772 5160
rect 9727 5120 9772 5148
rect 9766 5108 9772 5120
rect 9824 5148 9830 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 9824 5120 10333 5148
rect 9824 5108 9830 5120
rect 10321 5117 10333 5120
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 5460 5052 6960 5080
rect 4111 5015 4169 5021
rect 4111 5012 4123 5015
rect 4028 4984 4123 5012
rect 4028 4972 4034 4984
rect 4111 4981 4123 4984
rect 4157 4981 4169 5015
rect 4111 4975 4169 4981
rect 4893 5015 4951 5021
rect 4893 4981 4905 5015
rect 4939 5012 4951 5015
rect 4982 5012 4988 5024
rect 4939 4984 4988 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 6638 5012 6644 5024
rect 6319 4984 6644 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 6932 5021 6960 5052
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 4981 6975 5015
rect 6917 4975 6975 4981
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 7892 4984 8953 5012
rect 7892 4972 7898 4984
rect 8941 4981 8953 4984
rect 8987 5012 8999 5015
rect 9582 5012 9588 5024
rect 8987 4984 9588 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7800 4780 8217 4808
rect 7800 4768 7806 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 5626 4740 5632 4752
rect 5587 4712 5632 4740
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 4430 4632 4436 4684
rect 4488 4681 4494 4684
rect 4488 4675 4526 4681
rect 4514 4641 4526 4675
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 4488 4635 4526 4641
rect 4488 4632 4494 4635
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7834 4672 7840 4684
rect 7795 4644 7840 4672
rect 7653 4635 7711 4641
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5810 4604 5816 4616
rect 5771 4576 5816 4604
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7558 4604 7564 4616
rect 6696 4576 7564 4604
rect 6696 4564 6702 4576
rect 7558 4564 7564 4576
rect 7616 4604 7622 4616
rect 7668 4604 7696 4635
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8846 4604 8852 4616
rect 7616 4576 8852 4604
rect 7616 4564 7622 4576
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 5077 4539 5135 4545
rect 5077 4505 5089 4539
rect 5123 4536 5135 4539
rect 5350 4536 5356 4548
rect 5123 4508 5356 4536
rect 5123 4505 5135 4508
rect 5077 4499 5135 4505
rect 5350 4496 5356 4508
rect 5408 4536 5414 4548
rect 6178 4536 6184 4548
rect 5408 4508 6184 4536
rect 5408 4496 5414 4508
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4571 4471 4629 4477
rect 4571 4468 4583 4471
rect 4387 4440 4583 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4571 4437 4583 4440
rect 4617 4468 4629 4471
rect 4890 4468 4896 4480
rect 4617 4440 4896 4468
rect 4617 4437 4629 4440
rect 4571 4431 4629 4437
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 5994 4468 6000 4480
rect 5776 4440 6000 4468
rect 5776 4428 5782 4440
rect 5994 4428 6000 4440
rect 6052 4468 6058 4480
rect 6457 4471 6515 4477
rect 6457 4468 6469 4471
rect 6052 4440 6469 4468
rect 6052 4428 6058 4440
rect 6457 4437 6469 4440
rect 6503 4437 6515 4471
rect 6457 4431 6515 4437
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7374 4468 7380 4480
rect 6963 4440 7380 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7374 4428 7380 4440
rect 7432 4468 7438 4480
rect 7650 4468 7656 4480
rect 7432 4440 7656 4468
rect 7432 4428 7438 4440
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8720 4440 8769 4468
rect 8720 4428 8726 4440
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 3789 4267 3847 4273
rect 3789 4233 3801 4267
rect 3835 4264 3847 4267
rect 3970 4264 3976 4276
rect 3835 4236 3976 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 4430 4264 4436 4276
rect 4391 4236 4436 4264
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8159 4236 8984 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 4948 4100 5273 4128
rect 4948 4088 4954 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5902 4128 5908 4140
rect 5863 4100 5908 4128
rect 5261 4091 5319 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6273 4131 6331 4137
rect 6273 4128 6285 4131
rect 6052 4100 6285 4128
rect 6052 4088 6058 4100
rect 6273 4097 6285 4100
rect 6319 4128 6331 4131
rect 8128 4128 8156 4227
rect 8846 4196 8852 4208
rect 8807 4168 8852 4196
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 8956 4140 8984 4236
rect 9582 4156 9588 4208
rect 9640 4156 9646 4208
rect 8754 4137 8760 4140
rect 6319 4100 8156 4128
rect 8720 4131 8760 4137
rect 6319 4097 6331 4100
rect 6273 4091 6331 4097
rect 5074 4060 5080 4072
rect 5035 4032 5080 4060
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 7208 4069 7236 4100
rect 8720 4097 8732 4131
rect 8720 4091 8760 4097
rect 8754 4088 8760 4091
rect 8812 4088 8818 4140
rect 8938 4128 8944 4140
rect 8899 4100 8944 4128
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9306 4128 9312 4140
rect 9267 4100 9312 4128
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9600 4128 9628 4156
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 9600 4100 10609 4128
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7340 4032 7757 4060
rect 7340 4020 7346 4032
rect 7745 4029 7757 4032
rect 7791 4060 7803 4063
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 7791 4032 9689 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 9677 4023 9735 4029
rect 9784 4032 10333 4060
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 5350 3992 5356 4004
rect 4203 3964 5356 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 6270 3952 6276 4004
rect 6328 3952 6334 4004
rect 8573 3995 8631 4001
rect 8573 3992 8585 3995
rect 7852 3964 8585 3992
rect 6288 3924 6316 3952
rect 7852 3936 7880 3964
rect 8573 3961 8585 3964
rect 8619 3992 8631 3995
rect 8662 3992 8668 4004
rect 8619 3964 8668 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 6638 3924 6644 3936
rect 6288 3896 6644 3924
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7834 3884 7840 3936
rect 7892 3884 7898 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8754 3924 8760 3936
rect 8527 3896 8760 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8754 3884 8760 3896
rect 8812 3924 8818 3936
rect 9784 3924 9812 4032
rect 10321 4029 10333 4032
rect 10367 4060 10379 4063
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10367 4032 10977 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 13538 4060 13544 4072
rect 13495 4032 13544 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13538 4020 13544 4032
rect 13596 4060 13602 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13596 4032 14013 4060
rect 13596 4020 13602 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 10137 3995 10195 4001
rect 10137 3961 10149 3995
rect 10183 3961 10195 3995
rect 10137 3955 10195 3961
rect 9950 3924 9956 3936
rect 8812 3896 9812 3924
rect 9911 3896 9956 3924
rect 8812 3884 8818 3896
rect 9950 3884 9956 3896
rect 10008 3924 10014 3936
rect 10152 3924 10180 3955
rect 13630 3924 13636 3936
rect 10008 3896 10180 3924
rect 13591 3896 13636 3924
rect 10008 3884 10014 3896
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5350 3720 5356 3732
rect 4939 3692 5356 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5350 3680 5356 3692
rect 5408 3720 5414 3732
rect 5626 3720 5632 3732
rect 5408 3692 5632 3720
rect 5408 3680 5414 3692
rect 5626 3680 5632 3692
rect 5684 3720 5690 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 5684 3692 6745 3720
rect 5684 3680 5690 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 10318 3720 10324 3732
rect 10279 3692 10324 3720
rect 6733 3683 6791 3689
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 11425 3723 11483 3729
rect 11425 3689 11437 3723
rect 11471 3720 11483 3723
rect 12802 3720 12808 3732
rect 11471 3692 12808 3720
rect 11471 3689 11483 3692
rect 11425 3683 11483 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 6178 3661 6184 3664
rect 6175 3652 6184 3661
rect 6139 3624 6184 3652
rect 6175 3615 6184 3624
rect 6178 3612 6184 3615
rect 6236 3612 6242 3664
rect 7101 3655 7159 3661
rect 7101 3621 7113 3655
rect 7147 3652 7159 3655
rect 8110 3652 8116 3664
rect 7147 3624 8116 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 8720 3624 9076 3652
rect 8720 3612 8726 3624
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 7742 3584 7748 3596
rect 7607 3556 7748 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 7742 3544 7748 3556
rect 7800 3584 7806 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 7800 3556 8953 3584
rect 7800 3544 7806 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 9048 3584 9076 3624
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9048 3556 9689 3584
rect 8941 3547 8999 3553
rect 9677 3553 9689 3556
rect 9723 3584 9735 3587
rect 9950 3584 9956 3596
rect 9723 3556 9956 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 11238 3584 11244 3596
rect 11199 3556 11244 3584
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 13446 3584 13452 3596
rect 13407 3556 13452 3584
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 290 3476 296 3528
rect 348 3516 354 3528
rect 1302 3516 1308 3528
rect 348 3488 1308 3516
rect 348 3476 354 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 4525 3519 4583 3525
rect 4525 3485 4537 3519
rect 4571 3516 4583 3519
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 4571 3488 5825 3516
rect 4571 3485 4583 3488
rect 4525 3479 4583 3485
rect 5813 3485 5825 3488
rect 5859 3516 5871 3519
rect 6822 3516 6828 3528
rect 5859 3488 6828 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8754 3516 8760 3528
rect 7975 3488 8760 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 7377 3451 7435 3457
rect 7377 3448 7389 3451
rect 5276 3420 7389 3448
rect 5276 3392 5304 3420
rect 7377 3417 7389 3420
rect 7423 3417 7435 3451
rect 7377 3411 7435 3417
rect 7726 3451 7784 3457
rect 7726 3417 7738 3451
rect 7772 3448 7784 3451
rect 8570 3448 8576 3460
rect 7772 3420 8576 3448
rect 7772 3417 7784 3420
rect 7726 3411 7784 3417
rect 5258 3380 5264 3392
rect 5219 3352 5264 3380
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5534 3380 5540 3392
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 7392 3380 7420 3411
rect 8570 3408 8576 3420
rect 8628 3448 8634 3460
rect 8938 3448 8944 3460
rect 8628 3420 8944 3448
rect 8628 3408 8634 3420
rect 8938 3408 8944 3420
rect 8996 3448 9002 3460
rect 9582 3448 9588 3460
rect 8996 3420 9588 3448
rect 8996 3408 9002 3420
rect 9582 3408 9588 3420
rect 9640 3448 9646 3460
rect 10060 3448 10088 3479
rect 10410 3448 10416 3460
rect 9640 3420 10416 3448
rect 9640 3408 9646 3420
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 7834 3380 7840 3392
rect 7392 3352 7840 3380
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8665 3383 8723 3389
rect 8665 3380 8677 3383
rect 8168 3352 8677 3380
rect 8168 3340 8174 3352
rect 8665 3349 8677 3352
rect 8711 3380 8723 3383
rect 8846 3380 8852 3392
rect 8711 3352 8852 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 9398 3380 9404 3392
rect 9359 3352 9404 3380
rect 9398 3340 9404 3352
rect 9456 3380 9462 3392
rect 9815 3383 9873 3389
rect 9815 3380 9827 3383
rect 9456 3352 9827 3380
rect 9456 3340 9462 3352
rect 9815 3349 9827 3352
rect 9861 3349 9873 3383
rect 9950 3380 9956 3392
rect 9911 3352 9956 3380
rect 9815 3343 9873 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 13630 3380 13636 3392
rect 13591 3352 13636 3380
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 5334 3179 5392 3185
rect 5334 3145 5346 3179
rect 5380 3176 5392 3179
rect 5534 3176 5540 3188
rect 5380 3148 5540 3176
rect 5380 3145 5392 3148
rect 5334 3139 5392 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 6086 3176 6092 3188
rect 5859 3148 6092 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7742 3176 7748 3188
rect 7703 3148 7748 3176
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 8849 3179 8907 3185
rect 8849 3176 8861 3179
rect 8812 3148 8861 3176
rect 8812 3136 8818 3148
rect 8849 3145 8861 3148
rect 8895 3145 8907 3179
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 8849 3139 8907 3145
rect 4709 3111 4767 3117
rect 4709 3077 4721 3111
rect 4755 3108 4767 3111
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 4755 3080 5457 3108
rect 4755 3077 4767 3080
rect 4709 3071 4767 3077
rect 5445 3077 5457 3080
rect 5491 3108 5503 3111
rect 7760 3108 7788 3136
rect 5491 3080 7788 3108
rect 5491 3077 5503 3080
rect 5445 3071 5503 3077
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 5123 3012 5549 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 5537 3009 5549 3012
rect 5583 3040 5595 3043
rect 5994 3040 6000 3052
rect 5583 3012 6000 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 7377 3043 7435 3049
rect 6687 3012 7328 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 4120 2944 4169 2972
rect 4120 2932 4126 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 7300 2972 7328 3012
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7423 3012 8340 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 8312 2984 8340 3012
rect 8110 2972 8116 2984
rect 7300 2944 8116 2972
rect 4157 2935 4215 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8864 2972 8892 3139
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11514 3176 11520 3188
rect 11296 3148 11520 3176
rect 11296 3136 11302 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 12768 3148 13001 3176
rect 12768 3136 12774 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 12989 3139 13047 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 8938 3068 8944 3120
rect 8996 3108 9002 3120
rect 9950 3108 9956 3120
rect 8996 3080 9956 3108
rect 8996 3068 9002 3080
rect 9950 3068 9956 3080
rect 10008 3108 10014 3120
rect 10045 3111 10103 3117
rect 10045 3108 10057 3111
rect 10008 3080 10057 3108
rect 10008 3068 10014 3080
rect 10045 3077 10057 3080
rect 10091 3077 10103 3111
rect 10045 3071 10103 3077
rect 11149 3111 11207 3117
rect 11149 3077 11161 3111
rect 11195 3108 11207 3111
rect 12526 3108 12532 3120
rect 11195 3080 12532 3108
rect 11195 3077 11207 3080
rect 11149 3071 11207 3077
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3108 12679 3111
rect 13170 3108 13176 3120
rect 12667 3080 13176 3108
rect 12667 3077 12679 3080
rect 12621 3071 12679 3077
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3040 9094 3052
rect 9398 3040 9404 3052
rect 9088 3012 9404 3040
rect 9088 3000 9094 3012
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8352 2944 9137 2972
rect 8352 2932 8358 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10778 2932 10784 2984
rect 10836 2972 10842 2984
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 10836 2944 10977 2972
rect 10836 2932 10842 2944
rect 10965 2941 10977 2944
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12710 2972 12716 2984
rect 12483 2944 12716 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 5169 2907 5227 2913
rect 5169 2873 5181 2907
rect 5215 2904 5227 2907
rect 5258 2904 5264 2916
rect 5215 2876 5264 2904
rect 5215 2873 5227 2876
rect 5169 2867 5227 2873
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 5718 2836 5724 2848
rect 4387 2808 5724 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6273 2839 6331 2845
rect 6273 2836 6285 2839
rect 6236 2808 6285 2836
rect 6236 2796 6242 2808
rect 6273 2805 6285 2808
rect 6319 2836 6331 2839
rect 8478 2836 8484 2848
rect 6319 2808 8484 2836
rect 6319 2805 6331 2808
rect 6273 2799 6331 2805
rect 8478 2796 8484 2808
rect 8536 2836 8542 2848
rect 10134 2836 10140 2848
rect 8536 2808 10140 2836
rect 8536 2796 8542 2808
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 7009 2635 7067 2641
rect 7009 2632 7021 2635
rect 6880 2604 7021 2632
rect 6880 2592 6886 2604
rect 7009 2601 7021 2604
rect 7055 2601 7067 2635
rect 7009 2595 7067 2601
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 9493 2635 9551 2641
rect 9493 2632 9505 2635
rect 8720 2604 9505 2632
rect 8720 2592 8726 2604
rect 9493 2601 9505 2604
rect 9539 2601 9551 2635
rect 9493 2595 9551 2601
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13722 2632 13728 2644
rect 13311 2604 13728 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4816 2496 4844 2592
rect 5258 2564 5264 2576
rect 5219 2536 5264 2564
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 6696 2536 7788 2564
rect 6696 2524 6702 2536
rect 4203 2468 4844 2496
rect 5169 2499 5227 2505
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5810 2496 5816 2508
rect 5215 2468 5816 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 7006 2496 7012 2508
rect 6411 2468 7012 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 7650 2496 7656 2508
rect 7611 2468 7656 2496
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 7760 2505 7788 2536
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 8202 2456 8208 2508
rect 8260 2496 8266 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 8260 2468 8309 2496
rect 8260 2456 8266 2468
rect 8297 2465 8309 2468
rect 8343 2496 8355 2499
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8343 2468 9045 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9732 2468 9781 2496
rect 9732 2456 9738 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9815 2468 10333 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10321 2465 10333 2468
rect 10367 2465 10379 2499
rect 10870 2496 10876 2508
rect 10783 2468 10876 2496
rect 10321 2459 10379 2465
rect 10870 2456 10876 2468
rect 10928 2496 10934 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 10928 2468 11437 2496
rect 10928 2456 10934 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 13078 2496 13084 2508
rect 13039 2468 13084 2496
rect 11425 2459 11483 2465
rect 13078 2456 13084 2468
rect 13136 2496 13142 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13136 2468 13645 2496
rect 13136 2456 13142 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 7668 2428 7696 2456
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 7668 2400 8677 2428
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 4338 2360 4344 2372
rect 4299 2332 4344 2360
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2360 10011 2363
rect 10686 2360 10692 2372
rect 9999 2332 10692 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11974 2360 11980 2372
rect 11103 2332 11980 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 11974 2320 11980 2332
rect 12032 2320 12038 2372
rect 6638 2292 6644 2304
rect 6599 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 8484 35640 8536 35692
rect 9312 35640 9364 35692
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 8208 35232 8260 35284
rect 5540 35096 5592 35148
rect 5632 35096 5684 35148
rect 5816 35096 5868 35148
rect 7656 35139 7708 35148
rect 7656 35105 7665 35139
rect 7665 35105 7699 35139
rect 7699 35105 7708 35139
rect 7656 35096 7708 35105
rect 5632 35003 5684 35012
rect 5632 34969 5641 35003
rect 5641 34969 5675 35003
rect 5675 34969 5684 35003
rect 5632 34960 5684 34969
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 4804 34688 4856 34740
rect 10968 34688 11020 34740
rect 13636 34731 13688 34740
rect 13636 34697 13645 34731
rect 13645 34697 13679 34731
rect 13679 34697 13688 34731
rect 13636 34688 13688 34697
rect 10140 34620 10192 34672
rect 5540 34484 5592 34536
rect 7656 34484 7708 34536
rect 8208 34484 8260 34536
rect 9312 34484 9364 34536
rect 9496 34527 9548 34536
rect 9496 34493 9505 34527
rect 9505 34493 9539 34527
rect 9539 34493 9548 34527
rect 9496 34484 9548 34493
rect 12532 34484 12584 34536
rect 5356 34391 5408 34400
rect 5356 34357 5365 34391
rect 5365 34357 5399 34391
rect 5399 34357 5408 34391
rect 5356 34348 5408 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 2136 31696 2188 31748
rect 3976 31696 4028 31748
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 5724 29044 5776 29096
rect 5816 29044 5868 29096
rect 3148 28976 3200 29028
rect 3516 28976 3568 29028
rect 12716 28976 12768 29028
rect 12808 28976 12860 29028
rect 3976 28908 4028 28960
rect 4344 28908 4396 28960
rect 8668 28908 8720 28960
rect 9312 28908 9364 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 5264 27548 5316 27600
rect 5724 27548 5776 27600
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 112 26868 164 26920
rect 1308 26868 1360 26920
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 7104 22423 7156 22432
rect 7104 22389 7113 22423
rect 7113 22389 7147 22423
rect 7147 22389 7156 22423
rect 7104 22380 7156 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 20 22108 72 22160
rect 388 22108 440 22160
rect 6644 22083 6696 22092
rect 6644 22049 6688 22083
rect 6688 22049 6696 22083
rect 8024 22083 8076 22092
rect 6644 22040 6696 22049
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 6552 21972 6604 22024
rect 7656 22015 7708 22024
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 10508 21675 10560 21684
rect 10508 21641 10517 21675
rect 10517 21641 10551 21675
rect 10551 21641 10560 21675
rect 10508 21632 10560 21641
rect 6644 21607 6696 21616
rect 6644 21573 6653 21607
rect 6653 21573 6687 21607
rect 6687 21573 6696 21607
rect 6644 21564 6696 21573
rect 8116 21564 8168 21616
rect 7104 21496 7156 21548
rect 8116 21403 8168 21412
rect 7196 21335 7248 21344
rect 7196 21301 7205 21335
rect 7205 21301 7239 21335
rect 7239 21301 7248 21335
rect 8116 21369 8125 21403
rect 8125 21369 8159 21403
rect 8159 21369 8168 21403
rect 8116 21360 8168 21369
rect 7196 21292 7248 21301
rect 8024 21292 8076 21344
rect 8576 21292 8628 21344
rect 10784 21292 10836 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 7104 21088 7156 21140
rect 7196 21020 7248 21072
rect 7932 21063 7984 21072
rect 7932 21029 7941 21063
rect 7941 21029 7975 21063
rect 7975 21029 7984 21063
rect 7932 21020 7984 21029
rect 8116 21020 8168 21072
rect 9772 20995 9824 21004
rect 9772 20961 9790 20995
rect 9790 20961 9824 20995
rect 9772 20952 9824 20961
rect 8300 20884 8352 20936
rect 9680 20748 9732 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 7656 20587 7708 20596
rect 7656 20553 7665 20587
rect 7665 20553 7699 20587
rect 7699 20553 7708 20587
rect 7656 20544 7708 20553
rect 8300 20476 8352 20528
rect 9588 20544 9640 20596
rect 7288 20247 7340 20256
rect 7288 20213 7297 20247
rect 7297 20213 7331 20247
rect 7331 20213 7340 20247
rect 7288 20204 7340 20213
rect 7656 20204 7708 20256
rect 8300 20272 8352 20324
rect 9772 20247 9824 20256
rect 9772 20213 9781 20247
rect 9781 20213 9815 20247
rect 9815 20213 9824 20247
rect 9772 20204 9824 20213
rect 10968 20204 11020 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 8116 20000 8168 20052
rect 8576 20000 8628 20052
rect 8024 19975 8076 19984
rect 8024 19941 8033 19975
rect 8033 19941 8067 19975
rect 8067 19941 8076 19975
rect 8024 19932 8076 19941
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 8116 19456 8168 19508
rect 4068 19320 4120 19372
rect 4344 19320 4396 19372
rect 8668 19320 8720 19372
rect 8760 19320 8812 19372
rect 12624 19320 12676 19372
rect 12900 19320 12952 19372
rect 6920 19295 6972 19304
rect 6920 19261 6929 19295
rect 6929 19261 6963 19295
rect 6963 19261 6972 19295
rect 6920 19252 6972 19261
rect 12348 19252 12400 19304
rect 12532 19252 12584 19304
rect 6828 19227 6880 19236
rect 6828 19193 6837 19227
rect 6837 19193 6871 19227
rect 6871 19193 6880 19227
rect 6828 19184 6880 19193
rect 8024 19116 8076 19168
rect 8392 19116 8444 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 5632 18819 5684 18828
rect 5632 18785 5650 18819
rect 5650 18785 5684 18819
rect 9496 18912 9548 18964
rect 11336 18912 11388 18964
rect 6828 18844 6880 18896
rect 5632 18776 5684 18785
rect 11060 18776 11112 18828
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 7196 18683 7248 18692
rect 7196 18649 7205 18683
rect 7205 18649 7239 18683
rect 7239 18649 7248 18683
rect 7196 18640 7248 18649
rect 8300 18572 8352 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 4160 18368 4212 18420
rect 5632 18411 5684 18420
rect 5632 18377 5641 18411
rect 5641 18377 5675 18411
rect 5675 18377 5684 18411
rect 5632 18368 5684 18377
rect 6828 18368 6880 18420
rect 6920 18368 6972 18420
rect 3056 18300 3108 18352
rect 5816 18300 5868 18352
rect 7196 18300 7248 18352
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 7288 18232 7340 18241
rect 8300 18232 8352 18284
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 6644 18096 6696 18148
rect 6920 18139 6972 18148
rect 6920 18105 6929 18139
rect 6929 18105 6963 18139
rect 6963 18105 6972 18139
rect 6920 18096 6972 18105
rect 7104 18096 7156 18148
rect 8116 18139 8168 18148
rect 8116 18105 8125 18139
rect 8125 18105 8159 18139
rect 8159 18105 8168 18139
rect 8116 18096 8168 18105
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 11060 18028 11112 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 5448 17824 5500 17833
rect 6644 17824 6696 17876
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 6828 17756 6880 17808
rect 7288 17799 7340 17808
rect 7288 17765 7297 17799
rect 7297 17765 7331 17799
rect 7331 17765 7340 17799
rect 7288 17756 7340 17765
rect 10232 17756 10284 17808
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 7104 17620 7156 17672
rect 9864 17620 9916 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 11060 17620 11112 17672
rect 6920 17484 6972 17536
rect 10140 17484 10192 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 6828 17280 6880 17332
rect 9864 17323 9916 17332
rect 6644 17212 6696 17264
rect 6920 17144 6972 17196
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 10232 17280 10284 17332
rect 10600 17255 10652 17264
rect 10600 17221 10609 17255
rect 10609 17221 10643 17255
rect 10643 17221 10652 17255
rect 10600 17212 10652 17221
rect 6644 17076 6696 17128
rect 6184 16940 6236 16992
rect 8300 17051 8352 17060
rect 8300 17017 8309 17051
rect 8309 17017 8343 17051
rect 8343 17017 8352 17051
rect 8300 17008 8352 17017
rect 10048 17051 10100 17060
rect 10048 17017 10057 17051
rect 10057 17017 10091 17051
rect 10091 17017 10100 17051
rect 10048 17008 10100 17017
rect 10140 17051 10192 17060
rect 10140 17017 10149 17051
rect 10149 17017 10183 17051
rect 10183 17017 10192 17051
rect 10140 17008 10192 17017
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 8116 16779 8168 16788
rect 8116 16745 8125 16779
rect 8125 16745 8159 16779
rect 8159 16745 8168 16779
rect 8116 16736 8168 16745
rect 10140 16736 10192 16788
rect 7840 16668 7892 16720
rect 9772 16668 9824 16720
rect 11704 16668 11756 16720
rect 6092 16600 6144 16652
rect 6828 16600 6880 16652
rect 7288 16532 7340 16584
rect 7748 16532 7800 16584
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 11060 16532 11112 16584
rect 10048 16464 10100 16516
rect 6644 16396 6696 16448
rect 9404 16439 9456 16448
rect 9404 16405 9413 16439
rect 9413 16405 9447 16439
rect 9447 16405 9456 16439
rect 9404 16396 9456 16405
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 8392 16192 8444 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 6184 15988 6236 16040
rect 7748 15988 7800 16040
rect 8760 15988 8812 16040
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 11152 16031 11204 16040
rect 11152 15997 11196 16031
rect 11196 15997 11204 16031
rect 11152 15988 11204 15997
rect 7840 15920 7892 15972
rect 6092 15852 6144 15904
rect 9588 15920 9640 15972
rect 9772 15963 9824 15972
rect 9772 15929 9775 15963
rect 9775 15929 9809 15963
rect 9809 15929 9824 15963
rect 9772 15920 9824 15929
rect 10416 15920 10468 15972
rect 9404 15852 9456 15904
rect 9496 15852 9548 15904
rect 11704 15920 11756 15972
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 8852 15648 8904 15700
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 9772 15648 9824 15700
rect 6644 15623 6696 15632
rect 6644 15589 6653 15623
rect 6653 15589 6687 15623
rect 6687 15589 6696 15623
rect 6644 15580 6696 15589
rect 7840 15623 7892 15632
rect 7840 15589 7843 15623
rect 7843 15589 7877 15623
rect 7877 15589 7892 15623
rect 7840 15580 7892 15589
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 10048 15580 10100 15632
rect 6000 15555 6052 15564
rect 6000 15521 6009 15555
rect 6009 15521 6043 15555
rect 6043 15521 6052 15555
rect 6000 15512 6052 15521
rect 6920 15512 6972 15564
rect 7564 15444 7616 15496
rect 10416 15444 10468 15496
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 6000 15147 6052 15156
rect 6000 15113 6009 15147
rect 6009 15113 6043 15147
rect 6043 15113 6052 15147
rect 6000 15104 6052 15113
rect 7840 15104 7892 15156
rect 10416 15104 10468 15156
rect 8116 14968 8168 15020
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 9496 14900 9548 14952
rect 6920 14764 6972 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 9680 14560 9732 14612
rect 6184 14535 6236 14544
rect 6184 14501 6187 14535
rect 6187 14501 6221 14535
rect 6221 14501 6236 14535
rect 6184 14492 6236 14501
rect 8760 14535 8812 14544
rect 8760 14501 8769 14535
rect 8769 14501 8803 14535
rect 8803 14501 8812 14535
rect 8760 14492 8812 14501
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8392 14424 8444 14476
rect 9680 14467 9732 14476
rect 6644 14356 6696 14408
rect 6736 14356 6788 14408
rect 6920 14356 6972 14408
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 10324 14424 10376 14476
rect 5356 14220 5408 14272
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 8392 14016 8444 14068
rect 9680 14016 9732 14068
rect 7840 13948 7892 14000
rect 8576 13948 8628 14000
rect 5448 13880 5500 13932
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 8668 13855 8720 13864
rect 6644 13812 6696 13821
rect 5356 13787 5408 13796
rect 5356 13753 5365 13787
rect 5365 13753 5399 13787
rect 5399 13753 5408 13787
rect 5908 13787 5960 13796
rect 5356 13744 5408 13753
rect 5908 13753 5917 13787
rect 5917 13753 5951 13787
rect 5951 13753 5960 13787
rect 5908 13744 5960 13753
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 6920 13744 6972 13796
rect 7840 13744 7892 13796
rect 8576 13744 8628 13796
rect 5172 13676 5224 13728
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 6000 13472 6052 13524
rect 6920 13515 6972 13524
rect 5172 13404 5224 13456
rect 5816 13404 5868 13456
rect 6092 13404 6144 13456
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 8024 13404 8076 13456
rect 7840 13379 7892 13388
rect 4620 13268 4672 13320
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 7656 13268 7708 13320
rect 9772 13268 9824 13320
rect 5356 13132 5408 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 8760 13132 8812 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 6828 12724 6880 12776
rect 7380 12792 7432 12844
rect 5080 12656 5132 12708
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 7840 12724 7892 12776
rect 9312 12792 9364 12844
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 5356 12656 5408 12665
rect 8116 12656 8168 12708
rect 8760 12656 8812 12708
rect 5172 12588 5224 12640
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 7656 12588 7708 12640
rect 9404 12631 9456 12640
rect 9404 12597 9413 12631
rect 9413 12597 9447 12631
rect 9447 12597 9456 12631
rect 9404 12588 9456 12597
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 5356 12384 5408 12436
rect 5448 12384 5500 12436
rect 8668 12427 8720 12436
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 9588 12384 9640 12436
rect 7656 12316 7708 12368
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8668 12291 8720 12300
rect 8668 12257 8677 12291
rect 8677 12257 8711 12291
rect 8711 12257 8720 12291
rect 8668 12248 8720 12257
rect 9588 12248 9640 12300
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 10876 12180 10928 12232
rect 5080 12044 5132 12096
rect 5448 12044 5500 12096
rect 6000 12044 6052 12096
rect 7840 12044 7892 12096
rect 10600 12044 10652 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 7380 11840 7432 11892
rect 8576 11883 8628 11892
rect 8576 11849 8585 11883
rect 8585 11849 8619 11883
rect 8619 11849 8628 11883
rect 8576 11840 8628 11849
rect 9772 11840 9824 11892
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 9036 11704 9088 11756
rect 9404 11704 9456 11756
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11980 11704 12032 11756
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 8576 11568 8628 11620
rect 10600 11611 10652 11620
rect 10600 11577 10609 11611
rect 10609 11577 10643 11611
rect 10643 11577 10652 11611
rect 10600 11568 10652 11577
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 7656 11296 7708 11348
rect 9036 11339 9088 11348
rect 9036 11305 9045 11339
rect 9045 11305 9079 11339
rect 9079 11305 9088 11339
rect 9036 11296 9088 11305
rect 9496 11339 9548 11348
rect 9496 11305 9505 11339
rect 9505 11305 9539 11339
rect 9539 11305 9548 11339
rect 9496 11296 9548 11305
rect 9772 11228 9824 11280
rect 8116 11203 8168 11212
rect 8116 11169 8160 11203
rect 8160 11169 8168 11203
rect 8116 11160 8168 11169
rect 10600 11160 10652 11212
rect 10876 11160 10928 11212
rect 11060 11160 11112 11212
rect 10968 11092 11020 11144
rect 10416 11024 10468 11076
rect 7104 10956 7156 11008
rect 8024 10956 8076 11008
rect 8208 10956 8260 11008
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 11060 10752 11112 10804
rect 12716 10752 12768 10804
rect 8116 10727 8168 10736
rect 8116 10693 8125 10727
rect 8125 10693 8159 10727
rect 8159 10693 8168 10727
rect 8116 10684 8168 10693
rect 10416 10616 10468 10668
rect 8576 10548 8628 10600
rect 9404 10548 9456 10600
rect 8852 10480 8904 10532
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 10876 10523 10928 10532
rect 9772 10412 9824 10464
rect 9864 10412 9916 10464
rect 10876 10489 10885 10523
rect 10885 10489 10919 10523
rect 10919 10489 10928 10523
rect 10876 10480 10928 10489
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 5356 10140 5408 10192
rect 8852 10140 8904 10192
rect 11520 10140 11572 10192
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 8116 10115 8168 10124
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8668 10072 8720 10124
rect 9588 10072 9640 10124
rect 11060 10004 11112 10056
rect 11980 10047 12032 10056
rect 9772 9936 9824 9988
rect 11152 9936 11204 9988
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 12624 10004 12676 10056
rect 11888 9936 11940 9988
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5356 9868 5408 9920
rect 7012 9868 7064 9920
rect 7104 9868 7156 9920
rect 7840 9868 7892 9920
rect 10968 9911 11020 9920
rect 10968 9877 10977 9911
rect 10977 9877 11011 9911
rect 11011 9877 11020 9911
rect 10968 9868 11020 9877
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 7472 9664 7524 9716
rect 5448 9596 5500 9648
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 4804 9528 4856 9580
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 8208 9528 8260 9580
rect 8024 9503 8076 9512
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 5540 9392 5592 9444
rect 7012 9392 7064 9444
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 11060 9596 11112 9648
rect 9312 9528 9364 9580
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9496 9460 9548 9512
rect 12624 9664 12676 9716
rect 8392 9392 8444 9444
rect 9680 9392 9732 9444
rect 11428 9460 11480 9512
rect 12440 9503 12492 9512
rect 12440 9469 12484 9503
rect 12484 9469 12492 9503
rect 12440 9460 12492 9469
rect 10692 9392 10744 9444
rect 10968 9392 11020 9444
rect 6000 9324 6052 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 8852 9324 8904 9376
rect 9404 9367 9456 9376
rect 9404 9333 9413 9367
rect 9413 9333 9447 9367
rect 9447 9333 9456 9367
rect 9404 9324 9456 9333
rect 11520 9324 11572 9376
rect 11980 9367 12032 9376
rect 11980 9333 11989 9367
rect 11989 9333 12023 9367
rect 12023 9333 12032 9367
rect 11980 9324 12032 9333
rect 13636 9324 13688 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 6644 9163 6696 9172
rect 6644 9129 6653 9163
rect 6653 9129 6687 9163
rect 6687 9129 6696 9163
rect 6644 9120 6696 9129
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 5080 9052 5132 9104
rect 9496 9052 9548 9104
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 7012 9027 7064 9036
rect 7012 8993 7021 9027
rect 7021 8993 7055 9027
rect 7055 8993 7064 9027
rect 7012 8984 7064 8993
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7104 8916 7156 8968
rect 7656 8916 7708 8968
rect 6000 8780 6052 8832
rect 8024 8984 8076 9036
rect 10048 8984 10100 9036
rect 11152 9052 11204 9104
rect 12164 9095 12216 9104
rect 12164 9061 12173 9095
rect 12173 9061 12207 9095
rect 12207 9061 12216 9095
rect 12164 9052 12216 9061
rect 9680 8916 9732 8968
rect 10692 8984 10744 9036
rect 13544 9027 13596 9036
rect 13544 8993 13588 9027
rect 13588 8993 13596 9027
rect 13544 8984 13596 8993
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 11152 8848 11204 8900
rect 11980 8848 12032 8900
rect 8116 8823 8168 8832
rect 8116 8789 8125 8823
rect 8125 8789 8159 8823
rect 8159 8789 8168 8823
rect 8116 8780 8168 8789
rect 8392 8780 8444 8832
rect 9496 8780 9548 8832
rect 12348 8780 12400 8832
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4712 8576 4764 8628
rect 7196 8576 7248 8628
rect 8116 8576 8168 8628
rect 9680 8576 9732 8628
rect 10048 8576 10100 8628
rect 12164 8576 12216 8628
rect 6184 8508 6236 8560
rect 6736 8508 6788 8560
rect 7840 8508 7892 8560
rect 8576 8508 8628 8560
rect 10692 8508 10744 8560
rect 11888 8508 11940 8560
rect 13544 8551 13596 8560
rect 13544 8517 13553 8551
rect 13553 8517 13587 8551
rect 13587 8517 13596 8551
rect 13544 8508 13596 8517
rect 5632 8440 5684 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 1492 8236 1544 8288
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 7656 8372 7708 8381
rect 8668 8440 8720 8492
rect 9312 8440 9364 8492
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 8852 8372 8904 8424
rect 9680 8415 9732 8424
rect 5356 8304 5408 8313
rect 4804 8236 4856 8288
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 5448 8236 5500 8288
rect 8392 8304 8444 8356
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 12440 8415 12492 8424
rect 12440 8381 12484 8415
rect 12484 8381 12492 8415
rect 12440 8372 12492 8381
rect 11060 8304 11112 8356
rect 12072 8304 12124 8356
rect 12624 8304 12676 8356
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 10600 8279 10652 8288
rect 10600 8245 10609 8279
rect 10609 8245 10643 8279
rect 10643 8245 10652 8279
rect 10600 8236 10652 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 7472 8032 7524 8084
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 8760 8032 8812 8084
rect 9680 8032 9732 8084
rect 5080 7964 5132 8016
rect 5724 7964 5776 8016
rect 8392 8007 8444 8016
rect 8392 7973 8401 8007
rect 8401 7973 8435 8007
rect 8435 7973 8444 8007
rect 8392 7964 8444 7973
rect 9864 8007 9916 8016
rect 9864 7973 9873 8007
rect 9873 7973 9907 8007
rect 9907 7973 9916 8007
rect 9864 7964 9916 7973
rect 10600 7964 10652 8016
rect 5356 7896 5408 7948
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 8300 7896 8352 7948
rect 7656 7828 7708 7880
rect 9956 7828 10008 7880
rect 10784 7828 10836 7880
rect 11152 7828 11204 7880
rect 12348 7828 12400 7880
rect 6644 7760 6696 7812
rect 10876 7760 10928 7812
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 5908 7692 5960 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 6644 7488 6696 7540
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 12348 7488 12400 7540
rect 7656 7352 7708 7404
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 5356 7148 5408 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 7472 7216 7524 7268
rect 8852 7216 8904 7268
rect 10600 7259 10652 7268
rect 10600 7225 10609 7259
rect 10609 7225 10643 7259
rect 10643 7225 10652 7259
rect 10600 7216 10652 7225
rect 6644 7148 6696 7157
rect 8300 7148 8352 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 8668 6944 8720 6996
rect 9588 6944 9640 6996
rect 9956 6944 10008 6996
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 4344 6808 4396 6860
rect 5448 6808 5500 6860
rect 7196 6808 7248 6860
rect 9680 6851 9732 6860
rect 9680 6817 9724 6851
rect 9724 6817 9732 6851
rect 9680 6808 9732 6817
rect 10968 6808 11020 6860
rect 3884 6672 3936 6724
rect 8116 6672 8168 6724
rect 8484 6604 8536 6656
rect 8852 6604 8904 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 4344 6443 4396 6452
rect 4344 6409 4353 6443
rect 4353 6409 4387 6443
rect 4387 6409 4396 6443
rect 4344 6400 4396 6409
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 8576 6400 8628 6452
rect 4712 6171 4764 6180
rect 4712 6137 4721 6171
rect 4721 6137 4755 6171
rect 4755 6137 4764 6171
rect 4712 6128 4764 6137
rect 5448 6128 5500 6180
rect 5908 6171 5960 6180
rect 5908 6137 5917 6171
rect 5917 6137 5951 6171
rect 5951 6137 5960 6171
rect 5908 6128 5960 6137
rect 6184 6060 6236 6112
rect 8300 6196 8352 6248
rect 9680 6171 9732 6180
rect 9680 6137 9689 6171
rect 9689 6137 9723 6171
rect 9723 6137 9732 6171
rect 9680 6128 9732 6137
rect 9312 6060 9364 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 4712 5856 4764 5908
rect 7196 5856 7248 5908
rect 7564 5856 7616 5908
rect 5448 5831 5500 5840
rect 5448 5797 5457 5831
rect 5457 5797 5491 5831
rect 5491 5797 5500 5831
rect 5448 5788 5500 5797
rect 7656 5788 7708 5840
rect 4252 5763 4304 5772
rect 4252 5729 4296 5763
rect 4296 5729 4304 5763
rect 4252 5720 4304 5729
rect 7288 5763 7340 5772
rect 7288 5729 7297 5763
rect 7297 5729 7331 5763
rect 7331 5729 7340 5763
rect 7288 5720 7340 5729
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 4068 5652 4120 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4068 5312 4120 5364
rect 4252 5312 4304 5364
rect 5540 5312 5592 5364
rect 3516 5287 3568 5296
rect 3516 5253 3525 5287
rect 3525 5253 3559 5287
rect 3559 5253 3568 5287
rect 3516 5244 3568 5253
rect 11336 5244 11388 5296
rect 3884 5040 3936 5092
rect 4804 5108 4856 5160
rect 6644 5151 6696 5160
rect 5356 5083 5408 5092
rect 3976 4972 4028 5024
rect 5356 5049 5359 5083
rect 5359 5049 5393 5083
rect 5393 5049 5408 5083
rect 5356 5040 5408 5049
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 7012 5151 7064 5160
rect 6644 5108 6696 5117
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 4988 4972 5040 5024
rect 6644 4972 6696 5024
rect 7840 4972 7892 5024
rect 9588 4972 9640 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 7748 4768 7800 4820
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 4436 4675 4488 4684
rect 4436 4641 4480 4675
rect 4480 4641 4488 4675
rect 7288 4675 7340 4684
rect 4436 4632 4488 4641
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 7840 4675 7892 4684
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 6644 4564 6696 4616
rect 7564 4564 7616 4616
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8852 4564 8904 4616
rect 5356 4496 5408 4548
rect 6184 4496 6236 4548
rect 4896 4428 4948 4480
rect 5724 4428 5776 4480
rect 6000 4428 6052 4480
rect 7380 4428 7432 4480
rect 7656 4428 7708 4480
rect 8668 4428 8720 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 3976 4224 4028 4276
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 4896 4088 4948 4140
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 6000 4088 6052 4140
rect 8852 4199 8904 4208
rect 8852 4165 8861 4199
rect 8861 4165 8895 4199
rect 8895 4165 8904 4199
rect 8852 4156 8904 4165
rect 9588 4156 9640 4208
rect 8760 4131 8812 4140
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 8760 4097 8766 4131
rect 8766 4097 8812 4131
rect 8760 4088 8812 4097
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 7288 4020 7340 4072
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5356 3952 5408 3961
rect 6276 3952 6328 4004
rect 8668 3952 8720 4004
rect 6644 3927 6696 3936
rect 6644 3893 6653 3927
rect 6653 3893 6687 3927
rect 6687 3893 6696 3927
rect 6644 3884 6696 3893
rect 7840 3884 7892 3936
rect 8760 3884 8812 3936
rect 13544 4020 13596 4072
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 13636 3927 13688 3936
rect 9956 3884 10008 3893
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 5356 3680 5408 3732
rect 5632 3680 5684 3732
rect 10324 3723 10376 3732
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 12808 3680 12860 3732
rect 6184 3655 6236 3664
rect 6184 3621 6187 3655
rect 6187 3621 6221 3655
rect 6221 3621 6236 3655
rect 6184 3612 6236 3621
rect 8116 3612 8168 3664
rect 8668 3612 8720 3664
rect 7748 3544 7800 3596
rect 9956 3544 10008 3596
rect 11244 3587 11296 3596
rect 11244 3553 11253 3587
rect 11253 3553 11287 3587
rect 11287 3553 11296 3587
rect 11244 3544 11296 3553
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 296 3476 348 3528
rect 1308 3476 1360 3528
rect 6828 3476 6880 3528
rect 8760 3476 8812 3528
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 8576 3408 8628 3460
rect 8944 3408 8996 3460
rect 9588 3408 9640 3460
rect 10416 3408 10468 3460
rect 7840 3383 7892 3392
rect 7840 3349 7849 3383
rect 7849 3349 7883 3383
rect 7883 3349 7892 3383
rect 7840 3340 7892 3349
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 8116 3340 8168 3392
rect 8852 3340 8904 3392
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9404 3340 9456 3349
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 5540 3136 5592 3188
rect 6092 3136 6144 3188
rect 7748 3179 7800 3188
rect 7748 3145 7757 3179
rect 7757 3145 7791 3179
rect 7791 3145 7800 3179
rect 7748 3136 7800 3145
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 8760 3136 8812 3188
rect 10416 3179 10468 3188
rect 6000 3000 6052 3052
rect 4068 2932 4120 2984
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 8300 2932 8352 2984
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11244 3136 11296 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 12716 3136 12768 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 8944 3068 8996 3120
rect 9956 3068 10008 3120
rect 12532 3068 12584 3120
rect 13176 3068 13228 3120
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9404 3000 9456 3052
rect 10784 2932 10836 2984
rect 12716 2932 12768 2984
rect 5264 2864 5316 2916
rect 5724 2796 5776 2848
rect 6184 2796 6236 2848
rect 8484 2796 8536 2848
rect 10140 2796 10192 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 6828 2592 6880 2644
rect 8668 2592 8720 2644
rect 13728 2592 13780 2644
rect 5264 2567 5316 2576
rect 5264 2533 5273 2567
rect 5273 2533 5307 2567
rect 5307 2533 5316 2567
rect 5264 2524 5316 2533
rect 6644 2524 6696 2576
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 8208 2456 8260 2508
rect 9680 2456 9732 2508
rect 10876 2499 10928 2508
rect 10876 2465 10885 2499
rect 10885 2465 10919 2499
rect 10919 2465 10928 2499
rect 10876 2456 10928 2465
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 4344 2363 4396 2372
rect 4344 2329 4353 2363
rect 4353 2329 4387 2363
rect 4387 2329 4396 2363
rect 4344 2320 4396 2329
rect 10692 2320 10744 2372
rect 11980 2320 12032 2372
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
<< metal2 >>
rect 386 39520 442 40000
rect 1214 39522 1270 40000
rect 1214 39520 1348 39522
rect 2134 39520 2190 40000
rect 3054 39520 3110 40000
rect 3882 39520 3938 40000
rect 4802 39520 4858 40000
rect 5722 39522 5778 40000
rect 5644 39520 5778 39522
rect 6550 39520 6606 40000
rect 7470 39522 7526 40000
rect 6932 39520 7526 39522
rect 8390 39520 8446 40000
rect 9218 39520 9274 40000
rect 10138 39520 10194 40000
rect 11058 39520 11114 40000
rect 11886 39520 11942 40000
rect 12806 39520 12862 40000
rect 13726 39520 13782 40000
rect 14554 39520 14610 40000
rect 15474 39520 15530 40000
rect 112 26920 164 26926
rect 112 26862 164 26868
rect 20 22160 72 22166
rect 20 22102 72 22108
rect 32 6225 60 22102
rect 124 16153 152 26862
rect 400 22166 428 39520
rect 1228 39494 1348 39520
rect 1320 26926 1348 39494
rect 2148 31754 2176 39520
rect 2136 31748 2188 31754
rect 2136 31690 2188 31696
rect 1308 26920 1360 26926
rect 1308 26862 1360 26868
rect 388 22160 440 22166
rect 388 22102 440 22108
rect 3068 18358 3096 39520
rect 3896 37210 3924 39520
rect 3528 37182 3924 37210
rect 3422 33416 3478 33425
rect 3422 33351 3478 33360
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 21049 3188 28970
rect 3436 22001 3464 33351
rect 3528 29034 3556 37182
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 4816 34746 4844 39520
rect 5644 39494 5764 39520
rect 5644 35154 5672 39494
rect 6564 37754 6592 39520
rect 6932 39494 7512 39520
rect 6564 37726 6776 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5632 35148 5684 35154
rect 5632 35090 5684 35096
rect 5816 35148 5868 35154
rect 5816 35090 5868 35096
rect 4804 34740 4856 34746
rect 4804 34682 4856 34688
rect 5552 34542 5580 35090
rect 5630 35048 5686 35057
rect 5630 34983 5632 34992
rect 5684 34983 5686 34992
rect 5632 34954 5684 34960
rect 5540 34536 5592 34542
rect 5460 34484 5540 34490
rect 5460 34478 5592 34484
rect 5460 34462 5580 34478
rect 5356 34400 5408 34406
rect 5356 34342 5408 34348
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3976 31748 4028 31754
rect 3976 31690 4028 31696
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3516 29028 3568 29034
rect 3516 28970 3568 28976
rect 3988 28966 4016 31690
rect 3976 28960 4028 28966
rect 3976 28902 4028 28908
rect 4344 28960 4396 28966
rect 4344 28902 4396 28908
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3422 21992 3478 22001
rect 3422 21927 3478 21936
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3146 21040 3202 21049
rect 3146 20975 3202 20984
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 4158 20088 4214 20097
rect 4158 20023 4214 20032
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 19258 4108 19314
rect 3988 19230 4108 19258
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 110 16144 166 16153
rect 110 16079 166 16088
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 1306 10704 1362 10713
rect 1306 10639 1362 10648
rect 18 6216 74 6225
rect 18 6151 74 6160
rect 846 3904 902 3913
rect 846 3839 902 3848
rect 296 3528 348 3534
rect 296 3470 348 3476
rect 308 480 336 3470
rect 860 480 888 3839
rect 1320 3534 1348 10639
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 2778 8392 2834 8401
rect 2700 8350 2778 8378
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 2134 8256 2190 8265
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1504 480 1532 8230
rect 2134 8191 2190 8200
rect 2148 480 2176 8191
rect 2700 480 2728 8350
rect 2778 8327 2834 8336
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3882 6760 3938 6769
rect 3882 6695 3884 6704
rect 3936 6695 3938 6704
rect 3884 6666 3936 6672
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3988 5352 4016 19230
rect 4172 18426 4200 20023
rect 4356 19378 4384 28902
rect 5264 27600 5316 27606
rect 5264 27542 5316 27548
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 5276 18057 5304 27542
rect 5368 22681 5396 34342
rect 5354 22672 5410 22681
rect 5354 22607 5410 22616
rect 5460 22522 5488 34462
rect 5828 29102 5856 35090
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 5724 29096 5776 29102
rect 5724 29038 5776 29044
rect 5816 29096 5868 29102
rect 5816 29038 5868 29044
rect 5736 27606 5764 29038
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 5368 22494 5488 22522
rect 5262 18048 5318 18057
rect 5262 17983 5318 17992
rect 5368 17218 5396 22494
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6552 22024 6604 22030
rect 6550 21992 6552 22001
rect 6604 21992 6606 22001
rect 6550 21927 6606 21936
rect 6656 21622 6684 22034
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5644 18426 5672 18770
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5446 18184 5502 18193
rect 5446 18119 5502 18128
rect 5460 17882 5488 18119
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5276 17190 5396 17218
rect 4250 16144 4306 16153
rect 4250 16079 4306 16088
rect 4264 5778 4292 16079
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6458 4384 6802
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5370 4108 5646
rect 4264 5370 4292 5714
rect 3896 5324 4016 5352
rect 4068 5364 4120 5370
rect 3516 5296 3568 5302
rect 3514 5264 3516 5273
rect 3568 5264 3570 5273
rect 3514 5199 3570 5208
rect 3896 5098 3924 5324
rect 4068 5306 4120 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4593 4016 4966
rect 3974 4584 4030 4593
rect 3974 4519 4030 4528
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3988 4282 4016 4519
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4080 4162 4108 5199
rect 4264 5137 4292 5306
rect 4250 5128 4306 5137
rect 4250 5063 4306 5072
rect 4448 4690 4476 15807
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13462 5212 13670
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 12782 4660 13262
rect 4620 12776 4672 12782
rect 4618 12744 4620 12753
rect 4672 12744 4674 12753
rect 4618 12679 4674 12688
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 5092 12102 5120 12650
rect 5184 12646 5212 13398
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4618 9072 4674 9081
rect 4618 9007 4620 9016
rect 4672 9007 4674 9016
rect 4620 8978 4672 8984
rect 4632 8090 4660 8978
rect 4724 8634 4752 9862
rect 4802 9616 4858 9625
rect 4858 9560 4936 9568
rect 4802 9551 4804 9560
rect 4856 9540 4936 9560
rect 4804 9522 4856 9528
rect 4802 8664 4858 8673
rect 4712 8628 4764 8634
rect 4802 8599 4858 8608
rect 4712 8570 4764 8576
rect 4816 8294 4844 8599
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5914 4752 6122
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5166 4844 5510
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4908 5012 4936 9540
rect 5080 9104 5132 9110
rect 5184 9092 5212 12582
rect 5132 9064 5212 9092
rect 5080 9046 5132 9052
rect 5092 8294 5120 9046
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8022 5120 8230
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 5170 7304 5226 7313
rect 5170 7239 5226 7248
rect 4816 4984 4936 5012
rect 4988 5024 5040 5030
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4448 4282 4476 4626
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 3988 4134 4108 4162
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3330 1456 3386 1465
rect 3330 1391 3386 1400
rect 3344 480 3372 1391
rect 3988 480 4016 4134
rect 4448 3913 4476 4218
rect 4434 3904 4490 3913
rect 4434 3839 4490 3848
rect 4066 3224 4122 3233
rect 4066 3159 4068 3168
rect 4120 3159 4122 3168
rect 4068 3130 4120 3136
rect 4080 2990 4108 3130
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4816 2650 4844 4984
rect 4988 4966 5040 4972
rect 5000 4729 5028 4966
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4146 4936 4422
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5080 4072 5132 4078
rect 5078 4040 5080 4049
rect 5132 4040 5134 4049
rect 5078 3975 5134 3984
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4526 2544 4582 2553
rect 4526 2479 4582 2488
rect 4342 2408 4398 2417
rect 4342 2343 4344 2352
rect 4396 2343 4398 2352
rect 4344 2314 4396 2320
rect 4540 480 4568 2479
rect 5184 480 5212 7239
rect 5276 5273 5304 17190
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13802 5396 14214
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12714 5396 13126
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12442 5396 12650
rect 5460 12442 5488 13874
rect 5644 12458 5672 18362
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5722 18048 5778 18057
rect 5722 17983 5778 17992
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5619 12430 5672 12458
rect 5736 12458 5764 17983
rect 5828 13462 5856 18294
rect 6656 18154 6684 18702
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6656 17882 6684 18090
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 17270 6684 17614
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6644 17128 6696 17134
rect 6090 17096 6146 17105
rect 6644 17070 6696 17076
rect 6090 17031 6146 17040
rect 6104 16658 6132 17031
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6104 15910 6132 16594
rect 6196 16046 6224 16934
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6656 16454 6684 17070
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 15904 6144 15910
rect 6090 15872 6092 15881
rect 6144 15872 6146 15881
rect 6090 15807 6146 15816
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6012 15162 6040 15506
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5920 12850 5948 13738
rect 6012 13530 6040 15098
rect 6196 14550 6224 15982
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6656 15638 6684 16390
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6748 14498 6776 37726
rect 6932 19394 6960 39494
rect 8404 35306 8432 39520
rect 9232 37210 9260 39520
rect 9232 37182 9352 37210
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9324 35698 9352 37182
rect 8484 35692 8536 35698
rect 8484 35634 8536 35640
rect 9312 35692 9364 35698
rect 9312 35634 9364 35640
rect 8220 35290 8432 35306
rect 8208 35284 8432 35290
rect 8260 35278 8432 35284
rect 8208 35226 8260 35232
rect 7656 35148 7708 35154
rect 7656 35090 7708 35096
rect 7668 34542 7696 35090
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7116 21554 7144 22374
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7116 21146 7144 21490
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7208 21078 7236 21286
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7668 20602 7696 21966
rect 8036 21350 8064 22034
rect 8116 21616 8168 21622
rect 8116 21558 8168 21564
rect 8128 21418 8156 21558
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7668 20262 7696 20538
rect 7288 20256 7340 20262
rect 7286 20224 7288 20233
rect 7656 20256 7708 20262
rect 7340 20224 7342 20233
rect 7944 20233 7972 21014
rect 7656 20198 7708 20204
rect 7930 20224 7986 20233
rect 7286 20159 7342 20168
rect 7930 20159 7986 20168
rect 8036 19990 8064 21286
rect 8128 21078 8156 21354
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 6932 19366 7052 19394
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18902 6868 19178
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 18426 6868 18838
rect 6932 18426 6960 19246
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6840 17338 6868 17750
rect 6932 17542 6960 18090
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6932 17202 6960 17478
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6826 16688 6882 16697
rect 6826 16623 6828 16632
rect 6880 16623 6882 16632
rect 6828 16594 6880 16600
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6932 14822 6960 15506
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6196 13734 6224 14486
rect 6748 14470 6868 14498
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6656 13870 6684 14350
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6184 13728 6236 13734
rect 6748 13716 6776 14350
rect 6184 13670 6236 13676
rect 6656 13688 6776 13716
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5736 12430 5799 12458
rect 5619 12356 5647 12430
rect 5771 12424 5799 12430
rect 5771 12396 5856 12424
rect 5619 12328 5764 12356
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10198 5396 10406
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5368 9926 5396 10134
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9450 5396 9862
rect 5460 9654 5488 12038
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 9178 5580 9386
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5644 8498 5672 9998
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7954 5396 8298
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5262 5264 5318 5273
rect 5262 5199 5318 5208
rect 5368 5098 5396 7142
rect 5460 6866 5488 8230
rect 5644 7750 5672 8434
rect 5736 8265 5764 12328
rect 5828 9761 5856 12396
rect 5814 9752 5870 9761
rect 5814 9687 5870 9696
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5722 8256 5778 8265
rect 5722 8191 5778 8200
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5736 7206 5764 7958
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5846 5488 6122
rect 5448 5840 5500 5846
rect 5500 5788 5580 5794
rect 5448 5782 5580 5788
rect 5460 5766 5580 5782
rect 5552 5370 5580 5766
rect 5828 5710 5856 9590
rect 5920 8498 5948 12786
rect 6104 12458 6132 13398
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6656 12458 6684 13688
rect 6840 13546 6868 14470
rect 6932 14414 6960 14758
rect 7024 14498 7052 19366
rect 8036 19174 8064 19926
rect 8128 19514 8156 19994
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7208 18358 7236 18634
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7102 18184 7158 18193
rect 7102 18119 7104 18128
rect 7156 18119 7158 18128
rect 7104 18090 7156 18096
rect 7208 18034 7236 18294
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7116 18006 7236 18034
rect 7116 17678 7144 18006
rect 7300 17814 7328 18226
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 7288 17808 7340 17814
rect 7288 17750 7340 17756
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 8128 16794 8156 18090
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7300 15366 7328 16526
rect 7760 16046 7788 16526
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14822 7328 15302
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7024 14470 7328 14498
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6748 13518 6868 13546
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6748 12628 6776 13518
rect 6920 13466 6972 13472
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 12782 6868 13330
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 6932 12646 6960 12679
rect 6920 12640 6972 12646
rect 6748 12600 6868 12628
rect 6104 12430 6177 12458
rect 6656 12430 6776 12458
rect 6149 12424 6177 12430
rect 6149 12396 6224 12424
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 9382 6040 12038
rect 6090 9480 6146 9489
rect 6090 9415 6146 9424
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 8838 6040 9318
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 6186 5948 7686
rect 5908 6180 5960 6186
rect 5908 6122 5960 6128
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5368 4554 5396 5034
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4616 5592 4622
rect 5538 4584 5540 4593
rect 5592 4584 5594 4593
rect 5356 4548 5408 4554
rect 5538 4519 5594 4528
rect 5356 4490 5408 4496
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5368 3738 5396 3946
rect 5644 3738 5672 4694
rect 5828 4622 5856 5646
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5276 2922 5304 3334
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5552 3097 5580 3130
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 5736 2961 5764 4422
rect 5920 4146 5948 6122
rect 6012 4486 6040 8774
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6012 3058 6040 4082
rect 6104 3194 6132 9415
rect 6196 8566 6224 12396
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6748 9489 6776 12430
rect 6734 9480 6790 9489
rect 6734 9415 6790 9424
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 7818 6684 9114
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7546 6684 7754
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 4706 6224 6054
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6656 5166 6684 7142
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6196 4678 6316 4706
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 3670 6224 4490
rect 6288 4010 6316 4678
rect 6656 4622 6684 4966
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5722 2952 5778 2961
rect 5264 2916 5316 2922
rect 5722 2887 5778 2896
rect 5264 2858 5316 2864
rect 5276 2582 5304 2858
rect 5736 2854 5764 2887
rect 6196 2854 6224 3606
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6656 2582 6684 3878
rect 6748 3505 6776 8502
rect 6840 5114 6868 12600
rect 6920 12582 6972 12588
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 9926 7052 10406
rect 7116 9926 7144 10950
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7024 9450 7052 9862
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9081 6960 9318
rect 6918 9072 6974 9081
rect 7024 9042 7052 9386
rect 6918 9007 6974 9016
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7116 8974 7144 9454
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7208 8634 7236 8978
rect 7300 8945 7328 14470
rect 7576 14278 7604 15438
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7392 12306 7420 12786
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 11898 7420 12242
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7392 11778 7420 11834
rect 7392 11750 7512 11778
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7392 10470 7420 11630
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7286 8936 7342 8945
rect 7286 8871 7342 8880
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7208 6866 7236 8570
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7208 6458 7236 6802
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 5914 7236 6394
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7012 5160 7064 5166
rect 6840 5086 6960 5114
rect 7012 5102 7064 5108
rect 6932 3913 6960 5086
rect 6918 3904 6974 3913
rect 6918 3839 6974 3848
rect 6828 3528 6880 3534
rect 6734 3496 6790 3505
rect 6828 3470 6880 3476
rect 6734 3431 6790 3440
rect 6840 2650 6868 3470
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5828 480 5856 2450
rect 6656 2310 6684 2518
rect 7024 2514 7052 5102
rect 7300 4690 7328 5714
rect 7392 5166 7420 10406
rect 7484 10130 7512 11750
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7484 9722 7512 10066
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7484 8090 7512 9658
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7484 7274 7512 7890
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7576 5914 7604 14214
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12646 7696 13262
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12374 7696 12582
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7668 11762 7696 12310
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11354 7696 11698
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 8537 7696 8910
rect 7654 8528 7710 8537
rect 7654 8463 7710 8472
rect 7668 8430 7696 8463
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 7886 7696 8366
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7668 7410 7696 7822
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7656 5840 7708 5846
rect 7656 5782 7708 5788
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4078 7328 4626
rect 7392 4486 7420 5102
rect 7576 4622 7604 5714
rect 7668 5166 7696 5782
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7760 4826 7788 15982
rect 7852 15978 7880 16662
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7852 15638 7880 15914
rect 7840 15632 7892 15638
rect 7840 15574 7892 15580
rect 7852 15162 7880 15574
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7852 14006 7880 15098
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14482 8156 14962
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8022 14376 8078 14385
rect 8022 14311 8078 14320
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7852 13394 7880 13738
rect 8036 13462 8064 14311
rect 8128 13734 8156 14418
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 12782 7880 13330
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7852 12102 7880 12718
rect 8036 12594 8064 13398
rect 8128 12714 8156 13670
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 8036 12566 8156 12594
rect 8128 12306 8156 12566
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 8128 11370 8156 12242
rect 8036 11342 8156 11370
rect 8036 11014 8064 11342
rect 8220 11234 8248 34478
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8312 20534 8340 20878
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8312 20330 8340 20470
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8312 19854 8340 20266
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8312 18290 8340 18566
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17105 8340 17682
rect 8298 17096 8354 17105
rect 8298 17031 8300 17040
rect 8352 17031 8354 17040
rect 8300 17002 8352 17008
rect 8404 16250 8432 19110
rect 8496 17882 8524 35634
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 10152 34678 10180 39520
rect 10506 35728 10562 35737
rect 10506 35663 10562 35672
rect 10140 34672 10192 34678
rect 10140 34614 10192 34620
rect 9312 34536 9364 34542
rect 9312 34478 9364 34484
rect 9496 34536 9548 34542
rect 9496 34478 9548 34484
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9324 28966 9352 34478
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8588 20058 8616 21286
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8680 19378 8708 28902
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8850 20224 8906 20233
rect 8850 20159 8906 20168
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8772 17218 8800 19314
rect 8496 17190 8800 17218
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8404 14074 8432 14418
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8128 11218 8248 11234
rect 8116 11212 8248 11218
rect 8168 11206 8248 11212
rect 8116 11154 8168 11160
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10554 8064 10950
rect 8128 10742 8156 11154
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8116 10736 8168 10742
rect 8114 10704 8116 10713
rect 8168 10704 8170 10713
rect 8114 10639 8170 10648
rect 8036 10526 8156 10554
rect 8128 10130 8156 10526
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 8566 7880 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 9042 8064 9454
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8128 8838 8156 10066
rect 8220 10033 8248 10950
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8634 8156 8774
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 8128 6730 8156 8570
rect 8220 8242 8248 9522
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8838 8432 9386
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8362 8432 8774
rect 8496 8673 8524 17190
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 14550 8800 15982
rect 8864 15706 8892 20159
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9508 18970 9536 34478
rect 10520 21690 10548 35663
rect 11072 34762 11100 39520
rect 11900 37754 11928 39520
rect 11900 37726 12020 37754
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11992 35737 12020 37726
rect 11978 35728 12034 35737
rect 11978 35663 12034 35672
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 10980 34746 11100 34762
rect 10968 34740 11100 34746
rect 11020 34734 11100 34740
rect 10968 34682 11020 34688
rect 12532 34536 12584 34542
rect 12532 34478 12584 34484
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11334 30152 11390 30161
rect 11334 30087 11390 30096
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 9770 21040 9826 21049
rect 9770 20975 9772 20984
rect 9824 20975 9826 20984
rect 9772 20946 9824 20952
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20618 9720 20742
rect 9600 20602 9720 20618
rect 9588 20596 9720 20602
rect 9640 20590 9720 20596
rect 9588 20538 9640 20544
rect 9784 20262 9812 20946
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9876 17338 9904 17614
rect 10152 17542 10180 18158
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10244 17814 10272 18022
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 10152 17066 10180 17478
rect 10244 17338 10272 17750
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10612 17270 10640 17614
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9416 16046 9444 16390
rect 9404 16040 9456 16046
rect 9692 15994 9720 16594
rect 9404 15982 9456 15988
rect 9600 15978 9720 15994
rect 9784 15978 9812 16662
rect 10060 16522 10088 17002
rect 10152 16794 10180 17002
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9588 15972 9720 15978
rect 9640 15966 9720 15972
rect 9588 15914 9640 15920
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9416 15706 9444 15846
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9508 14958 9536 15846
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9692 14618 9720 15966
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15706 9812 15914
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 10060 15638 10088 16458
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9876 15026 9904 15574
rect 10428 15502 10456 15914
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15162 10456 15438
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9692 14385 9720 14418
rect 9678 14376 9734 14385
rect 9678 14311 9734 14320
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9692 14074 9720 14311
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8588 13802 8616 13942
rect 10336 13870 10364 14418
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 11898 8616 13738
rect 8680 13190 8708 13806
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8680 12442 8708 13126
rect 8772 12714 8800 13126
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8772 12322 8800 12650
rect 8680 12306 8800 12322
rect 8668 12300 8800 12306
rect 8720 12294 8800 12300
rect 8668 12242 8720 12248
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8588 11626 8616 11834
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10606 8616 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8680 10130 8708 12242
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11354 9076 11698
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 10198 8892 10474
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8864 9382 8892 10134
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9324 9586 9352 12786
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 11762 9444 12582
rect 9600 12442 9628 13670
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9588 12436 9640 12442
rect 9508 12396 9588 12424
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9508 11354 9536 12396
rect 9588 12378 9640 12384
rect 9692 12322 9720 12718
rect 9600 12306 9720 12322
rect 9588 12300 9720 12306
rect 9640 12294 9720 12300
rect 9588 12242 9640 12248
rect 9784 12238 9812 13262
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11898 9812 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8588 8430 8616 8502
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8220 8214 8340 8242
rect 8312 7954 8340 8214
rect 8404 8022 8432 8298
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7206 8340 7890
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8312 6254 8340 7142
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5030 7880 5714
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7852 4690 7880 4966
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7668 2514 7696 4422
rect 7852 4049 7880 4626
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 3194 7788 3538
rect 7852 3398 7880 3878
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8128 3398 8156 3606
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8036 3233 8064 3334
rect 8022 3224 8078 3233
rect 7748 3188 7800 3194
rect 8022 3159 8078 3168
rect 7748 3130 7800 3136
rect 8128 2990 8156 3334
rect 8116 2984 8168 2990
rect 8220 2961 8248 5102
rect 8312 4690 8340 6190
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8300 2984 8352 2990
rect 8116 2926 8168 2932
rect 8206 2952 8262 2961
rect 8300 2926 8352 2932
rect 8206 2887 8262 2896
rect 8220 2514 8248 2887
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 1850 6684 2246
rect 6380 1822 6684 1850
rect 6380 480 6408 1822
rect 7024 480 7052 2450
rect 7668 480 7696 2450
rect 8312 480 8340 2926
rect 8496 2854 8524 6598
rect 8588 6458 8616 8366
rect 8680 8090 8708 8434
rect 8864 8430 8892 9318
rect 9140 9178 9168 9454
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9324 8498 9352 9522
rect 9416 9382 9444 10542
rect 9784 10470 9812 11222
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9600 9466 9628 10066
rect 9784 9994 9812 10406
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9508 9110 9536 9454
rect 9600 9450 9720 9466
rect 9600 9444 9732 9450
rect 9600 9438 9680 9444
rect 9680 9386 9732 9392
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9586 9072 9642 9081
rect 9508 8838 9536 9046
rect 9586 9007 9642 9016
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 8090 8800 8230
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 7002 8708 7278
rect 8864 7274 8892 8366
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9600 7546 9628 9007
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8634 9720 8910
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8090 9720 8366
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8864 6662 8892 7210
rect 9784 7018 9812 9114
rect 9876 8022 9904 10406
rect 9954 10024 10010 10033
rect 9954 9959 10010 9968
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9876 7546 9904 7958
rect 9968 7886 9996 9959
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8634 10088 8978
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10060 8537 10088 8570
rect 10046 8528 10102 8537
rect 10046 8463 10102 8472
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9600 7002 9812 7018
rect 9968 7002 9996 7822
rect 9588 6996 9812 7002
rect 9640 6990 9812 6996
rect 9956 6996 10008 7002
rect 9588 6938 9640 6944
rect 9956 6938 10008 6944
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 9692 6225 9720 6802
rect 9678 6216 9734 6225
rect 9678 6151 9680 6160
rect 9732 6151 9734 6160
rect 9680 6122 9732 6128
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4010 8708 4422
rect 8864 4214 8892 4558
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8680 3670 8708 3946
rect 8772 3942 8800 4082
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8588 3194 8616 3402
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8680 2650 8708 3606
rect 8772 3534 8800 3878
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 3194 8800 3470
rect 8864 3398 8892 4150
rect 9324 4146 9352 6054
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4214 9628 4966
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8956 3466 8984 4082
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8864 3108 8892 3334
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8944 3120 8996 3126
rect 8864 3080 8944 3108
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8864 480 8892 3080
rect 8944 3062 8996 3068
rect 9034 3088 9090 3097
rect 9416 3058 9444 3334
rect 9034 3023 9036 3032
rect 9088 3023 9090 3032
rect 9404 3052 9456 3058
rect 9036 2994 9088 3000
rect 9404 2994 9456 3000
rect 9600 2530 9628 3402
rect 9508 2502 9628 2530
rect 9692 2514 9720 6122
rect 9772 5160 9824 5166
rect 9770 5128 9772 5137
rect 9824 5128 9826 5137
rect 9770 5063 9826 5072
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3602 9996 3878
rect 10336 3738 10364 13806
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11626 10640 12038
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10612 11218 10640 11562
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 10674 10456 11018
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9042 10732 9386
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10704 8566 10732 8978
rect 10692 8560 10744 8566
rect 10796 8537 10824 21286
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10980 16130 11008 20198
rect 11348 18970 11376 30087
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 12544 19310 12572 34478
rect 12820 31770 12848 39520
rect 13634 35184 13690 35193
rect 13634 35119 13690 35128
rect 13648 34746 13676 35119
rect 13740 35057 13768 39520
rect 14568 37210 14596 39520
rect 13832 37182 14596 37210
rect 13726 35048 13782 35057
rect 13726 34983 13782 34992
rect 13636 34740 13688 34746
rect 13636 34682 13688 34688
rect 12728 31742 12848 31770
rect 12728 29034 12756 31742
rect 12716 29028 12768 29034
rect 12716 28970 12768 28976
rect 12808 29028 12860 29034
rect 12808 28970 12860 28976
rect 12820 28914 12848 28970
rect 12820 28886 12940 28914
rect 12912 19378 12940 28886
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12636 19258 12664 19314
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18086 11100 18770
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17678 11100 18022
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11704 16720 11756 16726
rect 11058 16688 11114 16697
rect 11704 16662 11756 16668
rect 11058 16623 11114 16632
rect 11072 16590 11100 16623
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16250 11100 16526
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11150 16144 11206 16153
rect 10980 16102 11100 16130
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11762 10916 12174
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 11072 11218 11100 16102
rect 11150 16079 11206 16088
rect 11164 16046 11192 16079
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11716 15978 11744 16662
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10888 10538 10916 11154
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10692 8502 10744 8508
rect 10782 8528 10838 8537
rect 10782 8463 10838 8472
rect 10506 8392 10562 8401
rect 10506 8327 10562 8336
rect 10520 7410 10548 8327
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 8022 10640 8230
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 7002 10548 7346
rect 10612 7274 10640 7958
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7410 10824 7822
rect 10888 7818 10916 10474
rect 10980 9926 11008 11086
rect 11072 10810 11100 11154
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9450 11008 9862
rect 11072 9654 11100 9998
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 11164 9110 11192 9930
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11060 8356 11112 8362
rect 10980 8316 11060 8344
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10980 6866 11008 8316
rect 11060 8298 11112 8304
rect 11164 7886 11192 8842
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11440 7313 11468 9454
rect 11532 9382 11560 10134
rect 11992 10062 12020 11698
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11520 9376 11572 9382
rect 11900 9364 11928 9930
rect 12360 9636 12388 19246
rect 12636 19230 12756 19258
rect 12728 12322 12756 19230
rect 12728 12294 12848 12322
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12360 9608 12480 9636
rect 12452 9518 12480 9608
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 11980 9376 12032 9382
rect 11900 9336 11980 9364
rect 11520 9318 11572 9324
rect 11980 9318 12032 9324
rect 11532 9081 11560 9318
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11518 9072 11574 9081
rect 11518 9007 11574 9016
rect 11886 8936 11942 8945
rect 11992 8906 12020 9318
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11886 8871 11942 8880
rect 11980 8900 12032 8906
rect 11900 8566 11928 8871
rect 11980 8842 12032 8848
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 12084 8362 12112 8910
rect 12176 8634 12204 9046
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8356 12124 8362
rect 12072 8298 12124 8304
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 12360 7886 12388 8774
rect 12438 8528 12494 8537
rect 12438 8463 12494 8472
rect 12452 8430 12480 8463
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12622 8392 12678 8401
rect 12622 8327 12624 8336
rect 12676 8327 12678 8336
rect 12624 8298 12676 8304
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12360 7546 12388 7822
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 11426 7304 11482 7313
rect 11426 7239 11482 7248
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 10874 4720 10930 4729
rect 10874 4655 10930 4664
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10782 3496 10838 3505
rect 10416 3460 10468 3466
rect 10782 3431 10838 3440
rect 10416 3402 10468 3408
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3126 9996 3334
rect 10428 3194 10456 3402
rect 10796 3194 10824 3431
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10796 2990 10824 3130
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9680 2508 9732 2514
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 9508 480 9536 2502
rect 9680 2450 9732 2456
rect 10152 480 10180 2790
rect 10888 2514 10916 4655
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11256 3194 11284 3538
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10704 480 10732 2314
rect 11348 480 11376 5238
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 12728 3194 12756 10746
rect 12820 3738 12848 12294
rect 13634 10024 13690 10033
rect 13634 9959 13690 9968
rect 13648 9382 13676 9959
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8566 13584 8978
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13556 4078 13584 8502
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13450 3632 13506 3641
rect 13450 3567 13452 3576
rect 13504 3567 13506 3576
rect 13452 3538 13504 3544
rect 13464 3194 13492 3538
rect 13648 3505 13676 3878
rect 13634 3496 13690 3505
rect 13634 3431 13690 3440
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 11532 1465 11560 3130
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11518 1456 11574 1465
rect 11518 1391 11574 1400
rect 11992 480 12020 2314
rect 12544 480 12572 3062
rect 12728 2990 12756 3130
rect 13176 3120 13228 3126
rect 13648 3097 13676 3334
rect 13176 3062 13228 3068
rect 13634 3088 13690 3097
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 13082 2544 13138 2553
rect 13082 2479 13084 2488
rect 13136 2479 13138 2488
rect 13084 2450 13136 2456
rect 13188 480 13216 3062
rect 13634 3023 13690 3032
rect 13728 2644 13780 2650
rect 13832 2632 13860 37182
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 15488 35193 15516 39520
rect 15474 35184 15530 35193
rect 15474 35119 15530 35128
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13910 22672 13966 22681
rect 13910 22607 13966 22616
rect 13780 2604 13860 2632
rect 13728 2586 13780 2592
rect 13924 2428 13952 22607
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 15658 3496 15714 3505
rect 15658 3431 15714 3440
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 15014 3088 15070 3097
rect 15014 3023 15070 3032
rect 13832 2400 13952 2428
rect 14186 2408 14242 2417
rect 13832 480 13860 2400
rect 14186 2343 14242 2352
rect 14200 1986 14228 2343
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14200 1958 14412 1986
rect 14384 480 14412 1958
rect 15028 480 15056 3023
rect 15672 480 15700 3431
rect 294 0 350 480
rect 846 0 902 480
rect 1490 0 1546 480
rect 2134 0 2190 480
rect 2686 0 2742 480
rect 3330 0 3386 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5170 0 5226 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 7010 0 7066 480
rect 7654 0 7710 480
rect 8298 0 8354 480
rect 8850 0 8906 480
rect 9494 0 9550 480
rect 10138 0 10194 480
rect 10690 0 10746 480
rect 11334 0 11390 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13818 0 13874 480
rect 14370 0 14426 480
rect 15014 0 15070 480
rect 15658 0 15714 480
<< via2 >>
rect 3422 33360 3478 33416
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 5630 35012 5686 35048
rect 5630 34992 5632 35012
rect 5632 34992 5684 35012
rect 5684 34992 5686 35012
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3422 21936 3478 21992
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3146 20984 3202 21040
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 4158 20032 4214 20088
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 110 16088 166 16144
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 1306 10648 1362 10704
rect 18 6160 74 6216
rect 846 3848 902 3904
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 2134 8200 2190 8256
rect 2778 8336 2834 8392
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3882 6724 3938 6760
rect 3882 6704 3884 6724
rect 3884 6704 3936 6724
rect 3936 6704 3938 6724
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 5354 22616 5410 22672
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 5262 17992 5318 18048
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6550 21972 6552 21992
rect 6552 21972 6604 21992
rect 6604 21972 6606 21992
rect 6550 21936 6606 21972
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 5446 18128 5502 18184
rect 4250 16088 4306 16144
rect 4434 15816 4490 15872
rect 3514 5244 3516 5264
rect 3516 5244 3568 5264
rect 3568 5244 3570 5264
rect 3514 5208 3570 5244
rect 4066 5208 4122 5264
rect 3974 4528 4030 4584
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4250 5072 4306 5128
rect 4618 12724 4620 12744
rect 4620 12724 4672 12744
rect 4672 12724 4674 12744
rect 4618 12688 4674 12724
rect 4618 9036 4674 9072
rect 4618 9016 4620 9036
rect 4620 9016 4672 9036
rect 4672 9016 4674 9036
rect 4802 9580 4858 9616
rect 4802 9560 4804 9580
rect 4804 9560 4856 9580
rect 4856 9560 4858 9580
rect 4802 8608 4858 8664
rect 5170 7248 5226 7304
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3330 1400 3386 1456
rect 4434 3848 4490 3904
rect 4066 3188 4122 3224
rect 4066 3168 4068 3188
rect 4068 3168 4120 3188
rect 4120 3168 4122 3188
rect 4986 4664 5042 4720
rect 5078 4020 5080 4040
rect 5080 4020 5132 4040
rect 5132 4020 5134 4040
rect 5078 3984 5134 4020
rect 4526 2488 4582 2544
rect 4342 2372 4398 2408
rect 4342 2352 4344 2372
rect 4344 2352 4396 2372
rect 4396 2352 4398 2372
rect 5722 17992 5778 18048
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6090 17040 6146 17096
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6090 15852 6092 15872
rect 6092 15852 6144 15872
rect 6144 15852 6146 15872
rect 6090 15816 6146 15852
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 7286 20204 7288 20224
rect 7288 20204 7340 20224
rect 7340 20204 7342 20224
rect 7286 20168 7342 20204
rect 7930 20168 7986 20224
rect 6826 16652 6882 16688
rect 6826 16632 6828 16652
rect 6828 16632 6880 16652
rect 6880 16632 6882 16652
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 5262 5208 5318 5264
rect 5814 9696 5870 9752
rect 5722 8200 5778 8256
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 7102 18148 7158 18184
rect 7102 18128 7104 18148
rect 7104 18128 7156 18148
rect 7156 18128 7158 18148
rect 6918 12688 6974 12744
rect 6090 9424 6146 9480
rect 5538 4564 5540 4584
rect 5540 4564 5592 4584
rect 5592 4564 5594 4584
rect 5538 4528 5594 4564
rect 5538 3032 5594 3088
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6734 9424 6790 9480
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 5722 2896 5778 2952
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 6918 9016 6974 9072
rect 7286 8880 7342 8936
rect 6918 3848 6974 3904
rect 6734 3440 6790 3496
rect 7654 8472 7710 8528
rect 8022 14320 8078 14376
rect 8298 17060 8354 17096
rect 8298 17040 8300 17060
rect 8300 17040 8352 17060
rect 8352 17040 8354 17060
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 10506 35672 10562 35728
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8850 20168 8906 20224
rect 8114 10684 8116 10704
rect 8116 10684 8168 10704
rect 8168 10684 8170 10704
rect 8114 10648 8170 10684
rect 8206 9968 8262 10024
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11978 35672 12034 35728
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11334 30096 11390 30152
rect 9770 21004 9826 21040
rect 9770 20984 9772 21004
rect 9772 20984 9824 21004
rect 9824 20984 9826 21004
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 9678 14320 9734 14376
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8482 8608 8538 8664
rect 7838 3984 7894 4040
rect 8022 3168 8078 3224
rect 8206 2896 8262 2952
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 9586 9016 9642 9072
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 9954 9968 10010 10024
rect 10046 8472 10102 8528
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9678 6180 9734 6216
rect 9678 6160 9680 6180
rect 9680 6160 9732 6180
rect 9732 6160 9734 6180
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9034 3052 9090 3088
rect 9034 3032 9036 3052
rect 9036 3032 9088 3052
rect 9088 3032 9090 3052
rect 9770 5108 9772 5128
rect 9772 5108 9824 5128
rect 9824 5108 9826 5128
rect 9770 5072 9826 5108
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 13634 35128 13690 35184
rect 13726 34992 13782 35048
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11058 16632 11114 16688
rect 11150 16088 11206 16144
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 10782 8472 10838 8528
rect 10506 8336 10562 8392
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11518 9016 11574 9072
rect 11886 8880 11942 8936
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 12438 8472 12494 8528
rect 12622 8356 12678 8392
rect 12622 8336 12624 8356
rect 12624 8336 12676 8356
rect 12676 8336 12678 8356
rect 11426 7248 11482 7304
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 10874 4664 10930 4720
rect 10782 3440 10838 3496
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 13634 9968 13690 10024
rect 13450 3596 13506 3632
rect 13450 3576 13452 3596
rect 13452 3576 13504 3596
rect 13504 3576 13506 3596
rect 13634 3440 13690 3496
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 11518 1400 11574 1456
rect 13082 2508 13138 2544
rect 13082 2488 13084 2508
rect 13084 2488 13136 2508
rect 13136 2488 13138 2508
rect 13634 3032 13690 3088
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 15474 35128 15530 35184
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 13910 22616 13966 22672
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 15658 3440 15714 3496
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 15014 3032 15070 3088
rect 14186 2352 14242 2408
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 10501 35730 10567 35733
rect 11973 35730 12039 35733
rect 10501 35728 12039 35730
rect 10501 35672 10506 35728
rect 10562 35672 11978 35728
rect 12034 35672 12039 35728
rect 10501 35670 12039 35672
rect 10501 35667 10567 35670
rect 11973 35667 12039 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 13629 35186 13695 35189
rect 15469 35186 15535 35189
rect 13629 35184 15535 35186
rect 13629 35128 13634 35184
rect 13690 35128 15474 35184
rect 15530 35128 15535 35184
rect 13629 35126 15535 35128
rect 13629 35123 13695 35126
rect 15469 35123 15535 35126
rect 5625 35050 5691 35053
rect 13721 35050 13787 35053
rect 5625 35048 13787 35050
rect 5625 34992 5630 35048
rect 5686 34992 13726 35048
rect 13782 34992 13787 35048
rect 5625 34990 13787 34992
rect 5625 34987 5691 34990
rect 13721 34987 13787 34990
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 0 33418 480 33448
rect 3417 33418 3483 33421
rect 0 33416 3483 33418
rect 0 33360 3422 33416
rect 3478 33360 3483 33416
rect 0 33358 3483 33360
rect 0 33328 480 33358
rect 3417 33355 3483 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 11329 30154 11395 30157
rect 11329 30152 15532 30154
rect 11329 30096 11334 30152
rect 11390 30096 15532 30152
rect 11329 30094 15532 30096
rect 11329 30091 11395 30094
rect 15472 30048 15532 30094
rect 15472 29958 16000 30048
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 5349 22674 5415 22677
rect 13905 22674 13971 22677
rect 5349 22672 13971 22674
rect 5349 22616 5354 22672
rect 5410 22616 13910 22672
rect 13966 22616 13971 22672
rect 5349 22614 13971 22616
rect 5349 22611 5415 22614
rect 13905 22611 13971 22614
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 3417 21994 3483 21997
rect 6545 21994 6611 21997
rect 3417 21992 6611 21994
rect 3417 21936 3422 21992
rect 3478 21936 6550 21992
rect 6606 21936 6611 21992
rect 3417 21934 6611 21936
rect 3417 21931 3483 21934
rect 6545 21931 6611 21934
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3141 21042 3207 21045
rect 9765 21042 9831 21045
rect 3141 21040 9831 21042
rect 3141 20984 3146 21040
rect 3202 20984 9770 21040
rect 9826 20984 9831 21040
rect 3141 20982 9831 20984
rect 3141 20979 3207 20982
rect 9765 20979 9831 20982
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 7281 20226 7347 20229
rect 7925 20226 7991 20229
rect 8845 20226 8911 20229
rect 7281 20224 8911 20226
rect 7281 20168 7286 20224
rect 7342 20168 7930 20224
rect 7986 20168 8850 20224
rect 8906 20168 8911 20224
rect 7281 20166 8911 20168
rect 7281 20163 7347 20166
rect 7925 20163 7991 20166
rect 8845 20163 8911 20166
rect 6277 20160 6597 20161
rect 0 20090 480 20120
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 4153 20090 4219 20093
rect 0 20088 4219 20090
rect 0 20032 4158 20088
rect 4214 20032 4219 20088
rect 0 20030 4219 20032
rect 0 20000 480 20030
rect 4153 20027 4219 20030
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 5441 18186 5507 18189
rect 7097 18186 7163 18189
rect 5441 18184 7163 18186
rect 5441 18128 5446 18184
rect 5502 18128 7102 18184
rect 7158 18128 7163 18184
rect 5441 18126 7163 18128
rect 5441 18123 5507 18126
rect 7097 18123 7163 18126
rect 5257 18050 5323 18053
rect 5717 18050 5783 18053
rect 5257 18048 5783 18050
rect 5257 17992 5262 18048
rect 5318 17992 5722 18048
rect 5778 17992 5783 18048
rect 5257 17990 5783 17992
rect 5257 17987 5323 17990
rect 5717 17987 5783 17990
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 6085 17098 6151 17101
rect 8293 17098 8359 17101
rect 6085 17096 8359 17098
rect 6085 17040 6090 17096
rect 6146 17040 8298 17096
rect 8354 17040 8359 17096
rect 6085 17038 8359 17040
rect 6085 17035 6151 17038
rect 8293 17035 8359 17038
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 6821 16690 6887 16693
rect 11053 16690 11119 16693
rect 6821 16688 11119 16690
rect 6821 16632 6826 16688
rect 6882 16632 11058 16688
rect 11114 16632 11119 16688
rect 6821 16630 11119 16632
rect 6821 16627 6887 16630
rect 11053 16627 11119 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 105 16146 171 16149
rect 4245 16146 4311 16149
rect 11145 16146 11211 16149
rect 105 16144 11211 16146
rect 105 16088 110 16144
rect 166 16088 4250 16144
rect 4306 16088 11150 16144
rect 11206 16088 11211 16144
rect 105 16086 11211 16088
rect 105 16083 171 16086
rect 4245 16083 4311 16086
rect 11145 16083 11211 16086
rect 4429 15874 4495 15877
rect 6085 15874 6151 15877
rect 4429 15872 6151 15874
rect 4429 15816 4434 15872
rect 4490 15816 6090 15872
rect 6146 15816 6151 15872
rect 4429 15814 6151 15816
rect 4429 15811 4495 15814
rect 6085 15811 6151 15814
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 8017 14378 8083 14381
rect 9673 14378 9739 14381
rect 8017 14376 9739 14378
rect 8017 14320 8022 14376
rect 8078 14320 9678 14376
rect 9734 14320 9739 14376
rect 8017 14318 9739 14320
rect 8017 14315 8083 14318
rect 9673 14315 9739 14318
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 4613 12746 4679 12749
rect 6913 12746 6979 12749
rect 4613 12744 6979 12746
rect 4613 12688 4618 12744
rect 4674 12688 6918 12744
rect 6974 12688 6979 12744
rect 4613 12686 6979 12688
rect 4613 12683 4679 12686
rect 6913 12683 6979 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 1301 10706 1367 10709
rect 8109 10706 8175 10709
rect 1301 10704 8175 10706
rect 1301 10648 1306 10704
rect 1362 10648 8114 10704
rect 8170 10648 8175 10704
rect 1301 10646 8175 10648
rect 1301 10643 1367 10646
rect 8109 10643 8175 10646
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 8201 10026 8267 10029
rect 9949 10026 10015 10029
rect 8201 10024 10015 10026
rect 8201 9968 8206 10024
rect 8262 9968 9954 10024
rect 10010 9968 10015 10024
rect 8201 9966 10015 9968
rect 8201 9963 8267 9966
rect 9949 9963 10015 9966
rect 13629 10026 13695 10029
rect 15520 10026 16000 10056
rect 13629 10024 16000 10026
rect 13629 9968 13634 10024
rect 13690 9968 16000 10024
rect 13629 9966 16000 9968
rect 13629 9963 13695 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 5809 9754 5875 9757
rect 5766 9752 5875 9754
rect 5766 9696 5814 9752
rect 5870 9696 5875 9752
rect 5766 9691 5875 9696
rect 4797 9618 4863 9621
rect 5766 9618 5826 9691
rect 4797 9616 5826 9618
rect 4797 9560 4802 9616
rect 4858 9560 5826 9616
rect 4797 9558 5826 9560
rect 4797 9555 4863 9558
rect 6085 9482 6151 9485
rect 6729 9482 6795 9485
rect 6085 9480 6795 9482
rect 6085 9424 6090 9480
rect 6146 9424 6734 9480
rect 6790 9424 6795 9480
rect 6085 9422 6795 9424
rect 6085 9419 6151 9422
rect 6729 9419 6795 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 4613 9074 4679 9077
rect 6913 9074 6979 9077
rect 4613 9072 6979 9074
rect 4613 9016 4618 9072
rect 4674 9016 6918 9072
rect 6974 9016 6979 9072
rect 4613 9014 6979 9016
rect 4613 9011 4679 9014
rect 6913 9011 6979 9014
rect 9581 9074 9647 9077
rect 11513 9074 11579 9077
rect 9581 9072 11579 9074
rect 9581 9016 9586 9072
rect 9642 9016 11518 9072
rect 11574 9016 11579 9072
rect 9581 9014 11579 9016
rect 9581 9011 9647 9014
rect 11513 9011 11579 9014
rect 7281 8938 7347 8941
rect 11881 8938 11947 8941
rect 7281 8936 11947 8938
rect 7281 8880 7286 8936
rect 7342 8880 11886 8936
rect 11942 8880 11947 8936
rect 7281 8878 11947 8880
rect 7281 8875 7347 8878
rect 11881 8875 11947 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 4797 8666 4863 8669
rect 8477 8666 8543 8669
rect 4797 8664 8543 8666
rect 4797 8608 4802 8664
rect 4858 8608 8482 8664
rect 8538 8608 8543 8664
rect 4797 8606 8543 8608
rect 4797 8603 4863 8606
rect 8477 8603 8543 8606
rect 7649 8530 7715 8533
rect 10041 8530 10107 8533
rect 10777 8530 10843 8533
rect 12433 8530 12499 8533
rect 7649 8528 10107 8530
rect 7649 8472 7654 8528
rect 7710 8472 10046 8528
rect 10102 8472 10107 8528
rect 7649 8470 10107 8472
rect 7649 8467 7715 8470
rect 10041 8467 10107 8470
rect 10182 8528 12499 8530
rect 10182 8472 10782 8528
rect 10838 8472 12438 8528
rect 12494 8472 12499 8528
rect 10182 8470 12499 8472
rect 2773 8394 2839 8397
rect 10182 8394 10242 8470
rect 10777 8467 10843 8470
rect 12433 8467 12499 8470
rect 2773 8392 10242 8394
rect 2773 8336 2778 8392
rect 2834 8336 10242 8392
rect 2773 8334 10242 8336
rect 10501 8394 10567 8397
rect 12617 8394 12683 8397
rect 10501 8392 12683 8394
rect 10501 8336 10506 8392
rect 10562 8336 12622 8392
rect 12678 8336 12683 8392
rect 10501 8334 12683 8336
rect 2773 8331 2839 8334
rect 10501 8331 10567 8334
rect 12617 8331 12683 8334
rect 2129 8258 2195 8261
rect 5717 8258 5783 8261
rect 2129 8256 5783 8258
rect 2129 8200 2134 8256
rect 2190 8200 5722 8256
rect 5778 8200 5783 8256
rect 2129 8198 5783 8200
rect 2129 8195 2195 8198
rect 5717 8195 5783 8198
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 5165 7306 5231 7309
rect 11421 7306 11487 7309
rect 5165 7304 11487 7306
rect 5165 7248 5170 7304
rect 5226 7248 11426 7304
rect 11482 7248 11487 7304
rect 5165 7246 11487 7248
rect 5165 7243 5231 7246
rect 11421 7243 11487 7246
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 0 6762 480 6792
rect 3877 6762 3943 6765
rect 0 6760 3943 6762
rect 0 6704 3882 6760
rect 3938 6704 3943 6760
rect 0 6702 3943 6704
rect 0 6672 480 6702
rect 3877 6699 3943 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 13 6218 79 6221
rect 9673 6218 9739 6221
rect 13 6216 9739 6218
rect 13 6160 18 6216
rect 74 6160 9678 6216
rect 9734 6160 9739 6216
rect 13 6158 9739 6160
rect 13 6155 79 6158
rect 9673 6155 9739 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 3509 5266 3575 5269
rect 4061 5266 4127 5269
rect 5257 5266 5323 5269
rect 3509 5264 5323 5266
rect 3509 5208 3514 5264
rect 3570 5208 4066 5264
rect 4122 5208 5262 5264
rect 5318 5208 5323 5264
rect 3509 5206 5323 5208
rect 3509 5203 3575 5206
rect 4061 5203 4127 5206
rect 5257 5203 5323 5206
rect 4245 5130 4311 5133
rect 9765 5130 9831 5133
rect 4245 5128 9831 5130
rect 4245 5072 4250 5128
rect 4306 5072 9770 5128
rect 9826 5072 9831 5128
rect 4245 5070 9831 5072
rect 4245 5067 4311 5070
rect 9765 5067 9831 5070
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 4981 4722 5047 4725
rect 10869 4722 10935 4725
rect 4981 4720 10935 4722
rect 4981 4664 4986 4720
rect 5042 4664 10874 4720
rect 10930 4664 10935 4720
rect 4981 4662 10935 4664
rect 4981 4659 5047 4662
rect 10869 4659 10935 4662
rect 3969 4586 4035 4589
rect 5533 4586 5599 4589
rect 3969 4584 5599 4586
rect 3969 4528 3974 4584
rect 4030 4528 5538 4584
rect 5594 4528 5599 4584
rect 3969 4526 5599 4528
rect 3969 4523 4035 4526
rect 5533 4523 5599 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 5073 4042 5139 4045
rect 7833 4042 7899 4045
rect 5073 4040 7899 4042
rect 5073 3984 5078 4040
rect 5134 3984 7838 4040
rect 7894 3984 7899 4040
rect 5073 3982 7899 3984
rect 5073 3979 5139 3982
rect 7833 3979 7899 3982
rect 841 3906 907 3909
rect 4429 3906 4495 3909
rect 841 3904 4495 3906
rect 841 3848 846 3904
rect 902 3848 4434 3904
rect 4490 3848 4495 3904
rect 841 3846 4495 3848
rect 841 3843 907 3846
rect 4429 3843 4495 3846
rect 6913 3904 6979 3909
rect 6913 3848 6918 3904
rect 6974 3848 6979 3904
rect 6913 3843 6979 3848
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 6916 3634 6976 3843
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 13445 3634 13511 3637
rect 6916 3632 13511 3634
rect 6916 3576 13450 3632
rect 13506 3576 13511 3632
rect 6916 3574 13511 3576
rect 13445 3571 13511 3574
rect 6729 3498 6795 3501
rect 10777 3498 10843 3501
rect 6729 3496 10843 3498
rect 6729 3440 6734 3496
rect 6790 3440 10782 3496
rect 10838 3440 10843 3496
rect 6729 3438 10843 3440
rect 6729 3435 6795 3438
rect 10777 3435 10843 3438
rect 13629 3498 13695 3501
rect 15653 3498 15719 3501
rect 13629 3496 15719 3498
rect 13629 3440 13634 3496
rect 13690 3440 15658 3496
rect 15714 3440 15719 3496
rect 13629 3438 15719 3440
rect 13629 3435 13695 3438
rect 15653 3435 15719 3438
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 4061 3226 4127 3229
rect 8017 3226 8083 3229
rect 4061 3224 8083 3226
rect 4061 3168 4066 3224
rect 4122 3168 8022 3224
rect 8078 3168 8083 3224
rect 4061 3166 8083 3168
rect 4061 3163 4127 3166
rect 8017 3163 8083 3166
rect 5533 3090 5599 3093
rect 9029 3090 9095 3093
rect 5533 3088 9095 3090
rect 5533 3032 5538 3088
rect 5594 3032 9034 3088
rect 9090 3032 9095 3088
rect 5533 3030 9095 3032
rect 5533 3027 5599 3030
rect 9029 3027 9095 3030
rect 13629 3090 13695 3093
rect 15009 3090 15075 3093
rect 13629 3088 15075 3090
rect 13629 3032 13634 3088
rect 13690 3032 15014 3088
rect 15070 3032 15075 3088
rect 13629 3030 15075 3032
rect 13629 3027 13695 3030
rect 15009 3027 15075 3030
rect 5717 2954 5783 2957
rect 8201 2954 8267 2957
rect 5717 2952 8267 2954
rect 5717 2896 5722 2952
rect 5778 2896 8206 2952
rect 8262 2896 8267 2952
rect 5717 2894 8267 2896
rect 5717 2891 5783 2894
rect 8201 2891 8267 2894
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 4521 2546 4587 2549
rect 13077 2546 13143 2549
rect 4521 2544 13143 2546
rect 4521 2488 4526 2544
rect 4582 2488 13082 2544
rect 13138 2488 13143 2544
rect 4521 2486 13143 2488
rect 4521 2483 4587 2486
rect 13077 2483 13143 2486
rect 4337 2410 4403 2413
rect 14181 2410 14247 2413
rect 4337 2408 14247 2410
rect 4337 2352 4342 2408
rect 4398 2352 14186 2408
rect 14242 2352 14247 2408
rect 4337 2350 14247 2352
rect 4337 2347 4403 2350
rect 14181 2347 14247 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 3325 1458 3391 1461
rect 11513 1458 11579 1461
rect 3325 1456 11579 1458
rect 3325 1400 3330 1456
rect 3386 1400 11518 1456
rect 11574 1400 11579 1456
rect 3325 1398 11579 1400
rect 3325 1395 3391 1398
rect 11513 1395 11579 1398
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_1  _47_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _78_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_40 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__B
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__33__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _58_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _33_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__53__C
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_nor4_4  _53_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1602 592
use scs8hd_inv_8  _45_
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__C
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_82
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__D
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__B
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _54_
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__B
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_103
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _82_
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_115 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_114 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__88__A
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__58__D
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__C
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_42
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_50
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use scs8hd_or4_4  _46_
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__64__B
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__B
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_66
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__B
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__D
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use scs8hd_or4_4  _55_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__C
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _88_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_30
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__C
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _61_
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__64__D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _34_
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__34__C
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _62_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__B
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 774 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_39
timestamp 1586364061
transform 1 0 4692 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _64_
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__52__B
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__D
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__D
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _52_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__D
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__C
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_83
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 590 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_37
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _31_
timestamp 1586364061
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use scs8hd_nor4_4  _63_
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__C
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _35_
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_1  _32_
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_100
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_47
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _39_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_93
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _29_
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _37_
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__42__C
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__B
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__B
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _42_
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__C
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__D
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__41__C
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__D
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_104
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_137
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_145
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__50__D
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _50_
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__50__B
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__C
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__B
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_nor4_4  _41_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_38
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__D
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__B
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__B
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__D
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _51_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_nor4_4  _43_
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 1602 592
use scs8hd_nor4_4  _44_
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__D
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_89
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__C
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_137
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_133
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use scs8hd_buf_1  _40_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__36__B
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__C
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__D
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_inv_8  _30_
timestamp 1586364061
transform 1 0 6900 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_76
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_80
timestamp 1586364061
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_119
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _73_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_42
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use scs8hd_nor4_4  _36_
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__49__B
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__B
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__D
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__38__B
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_118
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_40
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_20_52
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 590 592
use scs8hd_nor4_4  _48_
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _49_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__C
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__C
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__D
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _38_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 1602 592
use scs8hd_conb_1  _71_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__C
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_96
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_120
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_120
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__D
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__B
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_70
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__B
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_113
timestamp 1586364061
transform 1 0 11500 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_121
timestamp 1586364061
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__B
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _57_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  FILLER_22_72
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _56_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _60_
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__B
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _66_
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_75
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _59_
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_114
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_138
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _74_
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_77
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__92__A
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_89
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_81
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 774 592
use scs8hd_conb_1  _72_
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_121
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _67_
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _92_
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_82
timestamp 1586364061
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_119
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_42
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_75
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use scs8hd_inv_8  _65_
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_111
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_51
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_112
timestamp 1586364061
transform 1 0 11408 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_124
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_136
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_inv_8  _68_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_91
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_103
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_82
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_90
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_52
timestamp 1586364061
transform 1 0 5888 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_70
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _69_
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_85
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_89
timestamp 1586364061
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_108
timestamp 1586364061
transform 1 0 11040 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_132
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_144
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8924 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_81
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use scs8hd_buf_2  _89_
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__89__A
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_104
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_108
timestamp 1586364061
transform 1 0 11040 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_120
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _70_
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_36_63
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_conb_1  _75_
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_68
timestamp 1586364061
transform 1 0 7360 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_104
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_141
timestamp 1586364061
transform 1 0 14076 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_141
timestamp 1586364061
transform 1 0 14076 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 5152 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _87_
timestamp 1586364061
transform 1 0 5428 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 5704 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_48
timestamp 1586364061
transform 1 0 5520 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_59_52
timestamp 1586364061
transform 1 0 5888 0 1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_51
timestamp 1586364061
transform 1 0 5796 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _93_
timestamp 1586364061
transform 1 0 7636 0 -1 35360
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__93__A
timestamp 1586364061
transform 1 0 7636 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_60
timestamp 1586364061
transform 1 0 6624 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_59_70
timestamp 1586364061
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_60_63
timestamp 1586364061
transform 1 0 6900 0 -1 35360
box -38 -48 774 592
use scs8hd_buf_2  _91_
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__91__A
timestamp 1586364061
transform 1 0 8924 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_73
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 590 592
use scs8hd_fill_2  FILLER_59_83
timestamp 1586364061
transform 1 0 8740 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_87
timestamp 1586364061
transform 1 0 9108 0 1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_75
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_87
timestamp 1586364061
transform 1 0 9108 0 -1 35360
box -38 -48 406 592
use scs8hd_buf_2  _90_
timestamp 1586364061
transform 1 0 9476 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__90__A
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_99
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_60_91
timestamp 1586364061
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_111
timestamp 1586364061
transform 1 0 11316 0 1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_59_119
timestamp 1586364061
transform 1 0 12052 0 1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 13432 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_131
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_138
timestamp 1586364061
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_142
timestamp 1586364061
transform 1 0 14168 0 1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 6366 0 6422 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 7010 0 7066 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 7654 0 7710 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 8298 0 8354 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 8850 0 8906 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 9494 0 9550 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 294 0 350 480 6 chany_bottom_in[0]
port 6 nsew default input
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[1]
port 7 nsew default input
rlabel metal2 s 1490 0 1546 480 6 chany_bottom_in[2]
port 8 nsew default input
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_in[3]
port 9 nsew default input
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_in[4]
port 10 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_in[5]
port 11 nsew default input
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_in[6]
port 12 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[7]
port 13 nsew default input
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_in[8]
port 14 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_out[0]
port 15 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_out[1]
port 16 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_out[2]
port 17 nsew default tristate
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_out[3]
port 18 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[4]
port 19 nsew default tristate
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_out[5]
port 20 nsew default tristate
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_out[6]
port 21 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[7]
port 22 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_out[8]
port 23 nsew default tristate
rlabel metal2 s 386 39520 442 40000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 1214 39520 1270 40000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 3054 39520 3110 40000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 3882 39520 3938 40000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 4802 39520 4858 40000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 7470 39520 7526 40000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 8390 39520 8446 40000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 9218 39520 9274 40000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 11058 39520 11114 40000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 11886 39520 11942 40000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 12806 39520 12862 40000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 15474 39520 15530 40000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 10138 0 10194 480 6 data_in
port 42 nsew default input
rlabel metal2 s 5814 0 5870 480 6 enable
port 43 nsew default input
rlabel metal3 s 0 6672 480 6792 6 left_grid_pin_1_
port 44 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 left_grid_pin_5_
port 45 nsew default tristate
rlabel metal3 s 0 33328 480 33448 6 left_grid_pin_9_
port 46 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 right_grid_pin_3_
port 47 nsew default tristate
rlabel metal3 s 15520 29928 16000 30048 6 right_grid_pin_7_
port 48 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 49 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 50 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
