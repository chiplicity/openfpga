magic
tech EFS8A
magscale 1 2
timestamp 1602532119
<< locali >>
rect 11287 22049 11322 22083
rect 12725 19295 12759 19397
rect 1443 18785 1478 18819
rect 12667 18785 12702 18819
rect 2547 17697 2582 17731
rect 10425 17187 10459 17289
rect 10051 16745 10057 16779
rect 10051 16677 10085 16745
rect 15485 16031 15519 16201
rect 4807 15895 4841 15963
rect 4807 15861 4813 15895
rect 8493 15419 8527 15521
rect 20027 13821 20062 13855
rect 3617 13379 3651 13481
rect 19199 13413 19244 13447
rect 9999 13345 10034 13379
rect 3341 12631 3375 12801
rect 19251 12393 19257 12427
rect 19251 12325 19285 12393
rect 20855 12257 20982 12291
rect 5733 11203 5767 11305
rect 13863 11169 13898 11203
rect 15703 11169 15830 11203
rect 5641 11067 5675 11169
rect 6561 9979 6595 10217
rect 23615 10081 23650 10115
rect 4629 9027 4663 9129
rect 4721 8959 4755 9129
rect 15669 8381 15795 8415
rect 4261 8279 4295 8381
rect 19349 7327 19383 7497
rect 24627 6817 24662 6851
rect 7113 6647 7147 6749
rect 4629 6239 4663 6273
rect 4629 6205 4790 6239
rect 5365 6103 5399 6409
rect 1547 5865 1685 5899
rect 13863 5729 13898 5763
rect 4721 5083 4755 5253
rect 8539 5185 8677 5219
rect 12265 5015 12299 5117
rect 12627 4777 12633 4811
rect 12627 4709 12661 4777
rect 14047 4641 14082 4675
rect 11483 3961 11621 3995
rect 5399 3553 5434 3587
rect 18463 3553 18498 3587
rect 3617 2941 3778 2975
rect 3617 2839 3651 2941
rect 4583 2533 4721 2567
<< viali >>
rect 1476 24225 1510 24259
rect 8344 24225 8378 24259
rect 1547 24021 1581 24055
rect 8447 24021 8481 24055
rect 1869 23817 1903 23851
rect 8769 23817 8803 23851
rect 9505 23817 9539 23851
rect 14749 23817 14783 23851
rect 19901 23817 19935 23851
rect 21649 23817 21683 23851
rect 25145 23817 25179 23851
rect 9137 23681 9171 23715
rect 1444 23613 1478 23647
rect 2237 23613 2271 23647
rect 6904 23613 6938 23647
rect 7297 23613 7331 23647
rect 8344 23613 8378 23647
rect 9321 23613 9355 23647
rect 9873 23613 9907 23647
rect 14565 23613 14599 23647
rect 16932 23613 16966 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 21465 23613 21499 23647
rect 22017 23613 22051 23647
rect 24660 23613 24694 23647
rect 1547 23477 1581 23511
rect 6975 23477 7009 23511
rect 8447 23477 8481 23511
rect 15209 23477 15243 23511
rect 17003 23477 17037 23511
rect 17417 23477 17451 23511
rect 24731 23477 24765 23511
rect 10103 23273 10137 23307
rect 1476 23137 1510 23171
rect 10032 23137 10066 23171
rect 1547 22933 1581 22967
rect 1593 22729 1627 22763
rect 9045 22729 9079 22763
rect 10149 22729 10183 22763
rect 24777 22729 24811 22763
rect 8861 22525 8895 22559
rect 9965 22525 9999 22559
rect 24593 22525 24627 22559
rect 25145 22525 25179 22559
rect 9505 22389 9539 22423
rect 9781 22389 9815 22423
rect 10517 22389 10551 22423
rect 11391 22185 11425 22219
rect 8284 22049 8318 22083
rect 9873 22049 9907 22083
rect 11253 22049 11287 22083
rect 8355 21845 8389 21879
rect 9965 21845 9999 21879
rect 10793 21845 10827 21879
rect 9367 21641 9401 21675
rect 8769 21505 8803 21539
rect 10517 21505 10551 21539
rect 10885 21505 10919 21539
rect 7573 21437 7607 21471
rect 8309 21437 8343 21471
rect 9264 21437 9298 21471
rect 10241 21369 10275 21403
rect 10609 21369 10643 21403
rect 8125 21301 8159 21335
rect 9045 21301 9079 21335
rect 9781 21301 9815 21335
rect 11437 21301 11471 21335
rect 1593 21097 1627 21131
rect 10057 21097 10091 21131
rect 7665 21029 7699 21063
rect 7849 21029 7883 21063
rect 7941 21029 7975 21063
rect 10333 21029 10367 21063
rect 10885 21029 10919 21063
rect 1409 20961 1443 20995
rect 6377 20961 6411 20995
rect 11805 20961 11839 20995
rect 22820 20961 22854 20995
rect 8125 20893 8159 20927
rect 10241 20893 10275 20927
rect 11713 20893 11747 20927
rect 6561 20757 6595 20791
rect 8769 20757 8803 20791
rect 22891 20757 22925 20791
rect 9873 20553 9907 20587
rect 11069 20553 11103 20587
rect 11713 20553 11747 20587
rect 14013 20553 14047 20587
rect 22845 20553 22879 20587
rect 9505 20485 9539 20519
rect 7021 20417 7055 20451
rect 8125 20417 8159 20451
rect 10057 20417 10091 20451
rect 12449 20417 12483 20451
rect 4721 20349 4755 20383
rect 5800 20349 5834 20383
rect 13528 20349 13562 20383
rect 8217 20281 8251 20315
rect 8769 20281 8803 20315
rect 10149 20281 10183 20315
rect 10701 20281 10735 20315
rect 1685 20213 1719 20247
rect 4905 20213 4939 20247
rect 5273 20213 5307 20247
rect 5871 20213 5905 20247
rect 6285 20213 6319 20247
rect 6653 20213 6687 20247
rect 7757 20213 7791 20247
rect 9045 20213 9079 20247
rect 13599 20213 13633 20247
rect 7205 19941 7239 19975
rect 8125 19941 8159 19975
rect 8217 19941 8251 19975
rect 8769 19941 8803 19975
rect 10057 19941 10091 19975
rect 10609 19941 10643 19975
rect 11621 19941 11655 19975
rect 13093 19941 13127 19975
rect 13185 19941 13219 19975
rect 4997 19873 5031 19907
rect 6561 19873 6595 19907
rect 4353 19805 4387 19839
rect 9965 19805 9999 19839
rect 11529 19805 11563 19839
rect 11805 19805 11839 19839
rect 13369 19805 13403 19839
rect 7665 19669 7699 19703
rect 14013 19669 14047 19703
rect 1593 19465 1627 19499
rect 3893 19465 3927 19499
rect 4997 19465 5031 19499
rect 6561 19465 6595 19499
rect 7389 19465 7423 19499
rect 10149 19465 10183 19499
rect 13277 19465 13311 19499
rect 5733 19397 5767 19431
rect 12725 19397 12759 19431
rect 12909 19397 12943 19431
rect 4353 19329 4387 19363
rect 8125 19329 8159 19363
rect 9045 19329 9079 19363
rect 10977 19329 11011 19363
rect 1409 19261 1443 19295
rect 1961 19261 1995 19295
rect 2580 19261 2614 19295
rect 5549 19261 5583 19295
rect 9137 19261 9171 19295
rect 9597 19261 9631 19295
rect 12516 19261 12550 19295
rect 12725 19261 12759 19295
rect 4077 19193 4111 19227
rect 4169 19193 4203 19227
rect 7665 19193 7699 19227
rect 7757 19193 7791 19227
rect 10333 19193 10367 19227
rect 10425 19193 10459 19227
rect 11805 19193 11839 19227
rect 13737 19193 13771 19227
rect 13829 19193 13863 19227
rect 14381 19193 14415 19227
rect 2651 19125 2685 19159
rect 3065 19125 3099 19159
rect 3433 19125 3467 19159
rect 6101 19125 6135 19159
rect 8585 19125 8619 19159
rect 9321 19125 9355 19159
rect 11437 19125 11471 19159
rect 12587 19125 12621 19159
rect 14657 19125 14691 19159
rect 1547 18921 1581 18955
rect 7665 18921 7699 18955
rect 8309 18921 8343 18955
rect 13093 18921 13127 18955
rect 5089 18853 5123 18887
rect 7107 18853 7141 18887
rect 10885 18853 10919 18887
rect 13829 18853 13863 18887
rect 14381 18853 14415 18887
rect 16497 18853 16531 18887
rect 16589 18853 16623 18887
rect 1409 18785 1443 18819
rect 8493 18785 8527 18819
rect 9724 18785 9758 18819
rect 12633 18785 12667 18819
rect 15368 18785 15402 18819
rect 2973 18717 3007 18751
rect 4997 18717 5031 18751
rect 6745 18717 6779 18751
rect 9827 18717 9861 18751
rect 10793 18717 10827 18751
rect 11253 18717 11287 18751
rect 13737 18717 13771 18751
rect 15945 18717 15979 18751
rect 16773 18717 16807 18751
rect 5549 18649 5583 18683
rect 10517 18649 10551 18683
rect 12771 18649 12805 18683
rect 7941 18581 7975 18615
rect 8677 18581 8711 18615
rect 10149 18581 10183 18615
rect 13461 18581 13495 18615
rect 15439 18581 15473 18615
rect 2329 18377 2363 18411
rect 4905 18377 4939 18411
rect 6009 18377 6043 18411
rect 6975 18377 7009 18411
rect 8769 18377 8803 18411
rect 11713 18377 11747 18411
rect 12265 18377 12299 18411
rect 15485 18377 15519 18411
rect 25145 18377 25179 18411
rect 2053 18309 2087 18343
rect 9045 18309 9079 18343
rect 13461 18309 13495 18343
rect 3525 18241 3559 18275
rect 4169 18241 4203 18275
rect 5089 18241 5123 18275
rect 5549 18241 5583 18275
rect 9689 18241 9723 18275
rect 12909 18241 12943 18275
rect 14749 18241 14783 18275
rect 16037 18241 16071 18275
rect 16313 18241 16347 18275
rect 1409 18173 1443 18207
rect 6904 18173 6938 18207
rect 7849 18173 7883 18207
rect 9505 18173 9539 18207
rect 11228 18173 11262 18207
rect 24660 18173 24694 18207
rect 3341 18105 3375 18139
rect 3617 18105 3651 18139
rect 5181 18105 5215 18139
rect 8170 18105 8204 18139
rect 9781 18105 9815 18139
rect 10333 18105 10367 18139
rect 13001 18105 13035 18139
rect 14289 18105 14323 18139
rect 14473 18105 14507 18139
rect 14565 18105 14599 18139
rect 16129 18105 16163 18139
rect 1593 18037 1627 18071
rect 4537 18037 4571 18071
rect 6653 18037 6687 18071
rect 7297 18037 7331 18071
rect 7757 18037 7791 18071
rect 10609 18037 10643 18071
rect 10977 18037 11011 18071
rect 11299 18037 11333 18071
rect 12633 18037 12667 18071
rect 13921 18037 13955 18071
rect 15761 18037 15795 18071
rect 16957 18037 16991 18071
rect 24731 18037 24765 18071
rect 1593 17833 1627 17867
rect 2053 17833 2087 17867
rect 3525 17833 3559 17867
rect 4353 17833 4387 17867
rect 7849 17833 7883 17867
rect 9413 17833 9447 17867
rect 10885 17833 10919 17867
rect 11161 17833 11195 17867
rect 12909 17833 12943 17867
rect 13553 17833 13587 17867
rect 16497 17833 16531 17867
rect 4629 17765 4663 17799
rect 4721 17765 4755 17799
rect 7291 17765 7325 17799
rect 9873 17765 9907 17799
rect 11529 17765 11563 17799
rect 13737 17765 13771 17799
rect 13829 17765 13863 17799
rect 16865 17765 16899 17799
rect 1409 17697 1443 17731
rect 2513 17697 2547 17731
rect 5641 17697 5675 17731
rect 15393 17697 15427 17731
rect 15761 17697 15795 17731
rect 2651 17629 2685 17663
rect 4905 17629 4939 17663
rect 6929 17629 6963 17663
rect 9781 17629 9815 17663
rect 10425 17629 10459 17663
rect 11437 17629 11471 17663
rect 14013 17629 14047 17663
rect 15853 17629 15887 17663
rect 11989 17561 12023 17595
rect 2329 17493 2363 17527
rect 2973 17493 3007 17527
rect 6837 17493 6871 17527
rect 4629 17289 4663 17323
rect 8769 17289 8803 17323
rect 9597 17289 9631 17323
rect 10241 17289 10275 17323
rect 10425 17289 10459 17323
rect 13001 17289 13035 17323
rect 14473 17289 14507 17323
rect 7389 17221 7423 17255
rect 14749 17221 14783 17255
rect 24777 17221 24811 17255
rect 3985 17153 4019 17187
rect 4905 17153 4939 17187
rect 5181 17153 5215 17187
rect 7849 17153 7883 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 10885 17153 10919 17187
rect 11529 17153 11563 17187
rect 16313 17153 16347 17187
rect 17233 17153 17267 17187
rect 1409 17085 1443 17119
rect 3157 17085 3191 17119
rect 3341 17085 3375 17119
rect 6904 17085 6938 17119
rect 12587 17085 12621 17119
rect 13553 17085 13587 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 4997 17017 5031 17051
rect 5825 17017 5859 17051
rect 6653 17017 6687 17051
rect 7757 17017 7791 17051
rect 8211 17017 8245 17051
rect 10977 17017 11011 17051
rect 12265 17017 12299 17051
rect 13915 17017 13949 17051
rect 16405 17017 16439 17051
rect 16957 17017 16991 17051
rect 1593 16949 1627 16983
rect 1961 16949 1995 16983
rect 2513 16949 2547 16983
rect 6193 16949 6227 16983
rect 6975 16949 7009 16983
rect 9781 16949 9815 16983
rect 11805 16949 11839 16983
rect 12679 16949 12713 16983
rect 13369 16949 13403 16983
rect 15393 16949 15427 16983
rect 15669 16949 15703 16983
rect 16129 16949 16163 16983
rect 1547 16745 1581 16779
rect 5365 16745 5399 16779
rect 5641 16745 5675 16779
rect 10057 16745 10091 16779
rect 10609 16745 10643 16779
rect 14657 16745 14691 16779
rect 4807 16677 4841 16711
rect 7205 16677 7239 16711
rect 12265 16677 12299 16711
rect 13737 16677 13771 16711
rect 13829 16677 13863 16711
rect 14381 16677 14415 16711
rect 16174 16677 16208 16711
rect 17785 16677 17819 16711
rect 1476 16609 1510 16643
rect 2513 16609 2547 16643
rect 2973 16609 3007 16643
rect 6469 16609 6503 16643
rect 6929 16609 6963 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 9689 16609 9723 16643
rect 15853 16609 15887 16643
rect 24593 16609 24627 16643
rect 3157 16541 3191 16575
rect 4445 16541 4479 16575
rect 7481 16541 7515 16575
rect 8769 16541 8803 16575
rect 12173 16541 12207 16575
rect 17049 16541 17083 16575
rect 17693 16541 17727 16575
rect 12725 16473 12759 16507
rect 18245 16473 18279 16507
rect 1869 16405 1903 16439
rect 2329 16405 2363 16439
rect 3433 16405 3467 16439
rect 3801 16405 3835 16439
rect 4353 16405 4387 16439
rect 7941 16405 7975 16439
rect 10885 16405 10919 16439
rect 13185 16405 13219 16439
rect 13461 16405 13495 16439
rect 16773 16405 16807 16439
rect 24777 16405 24811 16439
rect 2881 16201 2915 16235
rect 3893 16201 3927 16235
rect 5365 16201 5399 16235
rect 6101 16201 6135 16235
rect 9689 16201 9723 16235
rect 10609 16201 10643 16235
rect 11805 16201 11839 16235
rect 12587 16201 12621 16235
rect 15025 16201 15059 16235
rect 15485 16201 15519 16235
rect 15761 16201 15795 16235
rect 17693 16201 17727 16235
rect 24593 16201 24627 16235
rect 3617 16133 3651 16167
rect 13277 16133 13311 16167
rect 8769 16065 8803 16099
rect 11437 16065 11471 16099
rect 12173 16065 12207 16099
rect 13461 16065 13495 16099
rect 15347 16065 15381 16099
rect 16957 16065 16991 16099
rect 2053 15997 2087 16031
rect 3433 15997 3467 16031
rect 4445 15997 4479 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 7665 15997 7699 16031
rect 12484 15997 12518 16031
rect 14381 15997 14415 16031
rect 15260 15997 15294 16031
rect 15485 15997 15519 16031
rect 18112 15997 18146 16031
rect 18521 15997 18555 16031
rect 6469 15929 6503 15963
rect 7941 15929 7975 15963
rect 9131 15929 9165 15963
rect 10793 15929 10827 15963
rect 10885 15929 10919 15963
rect 12909 15929 12943 15963
rect 13782 15929 13816 15963
rect 14657 15929 14691 15963
rect 16313 15929 16347 15963
rect 16405 15929 16439 15963
rect 18199 15929 18233 15963
rect 1685 15861 1719 15895
rect 2513 15861 2547 15895
rect 3249 15861 3283 15895
rect 4353 15861 4387 15895
rect 4813 15861 4847 15895
rect 5641 15861 5675 15895
rect 8309 15861 8343 15895
rect 8677 15861 8711 15895
rect 9965 15861 9999 15895
rect 16037 15861 16071 15895
rect 17233 15861 17267 15895
rect 4721 15657 4755 15691
rect 6837 15657 6871 15691
rect 8125 15657 8159 15691
rect 9045 15657 9079 15691
rect 9413 15657 9447 15691
rect 13369 15657 13403 15691
rect 15853 15657 15887 15691
rect 17141 15657 17175 15691
rect 18061 15657 18095 15691
rect 1685 15589 1719 15623
rect 2237 15589 2271 15623
rect 4537 15589 4571 15623
rect 8677 15589 8711 15623
rect 10286 15589 10320 15623
rect 11897 15589 11931 15623
rect 16542 15589 16576 15623
rect 17693 15589 17727 15623
rect 4629 15521 4663 15555
rect 5273 15521 5307 15555
rect 5457 15521 5491 15555
rect 6009 15521 6043 15555
rect 6929 15521 6963 15555
rect 7389 15521 7423 15555
rect 7757 15521 7791 15555
rect 8309 15521 8343 15555
rect 8493 15521 8527 15555
rect 9965 15521 9999 15555
rect 13277 15521 13311 15555
rect 13829 15521 13863 15555
rect 14289 15521 14323 15555
rect 17969 15521 18003 15555
rect 18429 15521 18463 15555
rect 1593 15453 1627 15487
rect 11805 15453 11839 15487
rect 12081 15453 12115 15487
rect 16221 15453 16255 15487
rect 3893 15385 3927 15419
rect 6469 15385 6503 15419
rect 8493 15385 8527 15419
rect 11161 15385 11195 15419
rect 2605 15317 2639 15351
rect 2881 15317 2915 15351
rect 3433 15317 3467 15351
rect 10885 15317 10919 15351
rect 12725 15317 12759 15351
rect 1593 15113 1627 15147
rect 1961 15113 1995 15147
rect 4353 15113 4387 15147
rect 9551 15113 9585 15147
rect 11805 15113 11839 15147
rect 13461 15113 13495 15147
rect 15485 15113 15519 15147
rect 16589 15113 16623 15147
rect 17509 15113 17543 15147
rect 20177 15113 20211 15147
rect 3157 15045 3191 15079
rect 5825 15045 5859 15079
rect 8217 15045 8251 15079
rect 9321 15045 9355 15079
rect 2605 14977 2639 15011
rect 8585 14977 8619 15011
rect 12541 14977 12575 15011
rect 12817 14977 12851 15011
rect 17785 14977 17819 15011
rect 21557 14977 21591 15011
rect 1409 14909 1443 14943
rect 4629 14909 4663 14943
rect 5181 14909 5215 14943
rect 5273 14909 5307 14943
rect 5825 14909 5859 14943
rect 6837 14909 6871 14943
rect 7389 14909 7423 14943
rect 7665 14909 7699 14943
rect 8217 14909 8251 14943
rect 9448 14909 9482 14943
rect 9873 14909 9907 14943
rect 10425 14909 10459 14943
rect 14013 14909 14047 14943
rect 14105 14909 14139 14943
rect 14565 14909 14599 14943
rect 15669 14909 15703 14943
rect 18061 14909 18095 14943
rect 18521 14909 18555 14943
rect 19993 14909 20027 14943
rect 21164 14909 21198 14943
rect 2697 14841 2731 14875
rect 3985 14841 4019 14875
rect 10746 14841 10780 14875
rect 12265 14841 12299 14875
rect 12633 14841 12667 14875
rect 14841 14841 14875 14875
rect 15117 14841 15151 14875
rect 15990 14841 16024 14875
rect 16865 14841 16899 14875
rect 19073 14841 19107 14875
rect 2329 14773 2363 14807
rect 3617 14773 3651 14807
rect 6193 14773 6227 14807
rect 6561 14773 6595 14807
rect 10241 14773 10275 14807
rect 11345 14773 11379 14807
rect 18153 14773 18187 14807
rect 20637 14773 20671 14807
rect 21235 14773 21269 14807
rect 4353 14569 4387 14603
rect 4629 14569 4663 14603
rect 7205 14569 7239 14603
rect 9873 14569 9907 14603
rect 15577 14569 15611 14603
rect 17509 14569 17543 14603
rect 19073 14569 19107 14603
rect 2605 14501 2639 14535
rect 3157 14501 3191 14535
rect 7481 14501 7515 14535
rect 8769 14501 8803 14535
rect 10378 14501 10412 14535
rect 11621 14501 11655 14535
rect 11989 14501 12023 14535
rect 13461 14501 13495 14535
rect 13553 14501 13587 14535
rect 15990 14501 16024 14535
rect 16865 14501 16899 14535
rect 5089 14433 5123 14467
rect 6837 14433 6871 14467
rect 7021 14433 7055 14467
rect 8309 14433 8343 14467
rect 8493 14433 8527 14467
rect 15669 14433 15703 14467
rect 16589 14433 16623 14467
rect 17417 14433 17451 14467
rect 17877 14433 17911 14467
rect 18981 14433 19015 14467
rect 19441 14433 19475 14467
rect 21097 14433 21131 14467
rect 1409 14365 1443 14399
rect 2237 14365 2271 14399
rect 2513 14365 2547 14399
rect 5733 14365 5767 14399
rect 10057 14365 10091 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 13737 14365 13771 14399
rect 21741 14365 21775 14399
rect 3893 14297 3927 14331
rect 6193 14297 6227 14331
rect 1961 14229 1995 14263
rect 3525 14229 3559 14263
rect 6561 14229 6595 14263
rect 10977 14229 11011 14263
rect 13185 14229 13219 14263
rect 18429 14229 18463 14263
rect 20085 14229 20119 14263
rect 6285 14025 6319 14059
rect 9413 14025 9447 14059
rect 11529 14025 11563 14059
rect 11897 14025 11931 14059
rect 13921 14025 13955 14059
rect 17417 14025 17451 14059
rect 19809 14025 19843 14059
rect 20131 14025 20165 14059
rect 20637 14025 20671 14059
rect 21005 14025 21039 14059
rect 25145 14025 25179 14059
rect 3249 13957 3283 13991
rect 6653 13957 6687 13991
rect 14749 13957 14783 13991
rect 15669 13957 15703 13991
rect 17049 13957 17083 13991
rect 1501 13889 1535 13923
rect 8677 13889 8711 13923
rect 9045 13889 9079 13923
rect 10609 13889 10643 13923
rect 12173 13889 12207 13923
rect 16773 13889 16807 13923
rect 18889 13889 18923 13923
rect 21189 13889 21223 13923
rect 3893 13821 3927 13855
rect 4261 13821 4295 13855
rect 4537 13821 4571 13855
rect 5089 13821 5123 13855
rect 6837 13821 6871 13855
rect 7297 13821 7331 13855
rect 7757 13821 7791 13855
rect 8217 13821 8251 13855
rect 9321 13821 9355 13855
rect 14565 13821 14599 13855
rect 16037 13821 16071 13855
rect 16497 13821 16531 13855
rect 17785 13821 17819 13855
rect 19993 13821 20027 13855
rect 24660 13821 24694 13855
rect 1863 13753 1897 13787
rect 5549 13753 5583 13787
rect 9134 13753 9168 13787
rect 10971 13753 11005 13787
rect 13001 13753 13035 13787
rect 13093 13753 13127 13787
rect 13645 13753 13679 13787
rect 14289 13753 14323 13787
rect 18521 13753 18555 13787
rect 18613 13753 18647 13787
rect 21281 13753 21315 13787
rect 21833 13753 21867 13787
rect 2421 13685 2455 13719
rect 2789 13685 2823 13719
rect 3525 13685 3559 13719
rect 3801 13685 3835 13719
rect 5825 13685 5859 13719
rect 6929 13685 6963 13719
rect 10149 13685 10183 13719
rect 10425 13685 10459 13719
rect 12725 13685 12759 13719
rect 18245 13685 18279 13719
rect 19533 13685 19567 13719
rect 24731 13685 24765 13719
rect 3157 13481 3191 13515
rect 3617 13481 3651 13515
rect 3801 13481 3835 13515
rect 5917 13481 5951 13515
rect 6193 13481 6227 13515
rect 8217 13481 8251 13515
rect 9137 13481 9171 13515
rect 10701 13481 10735 13515
rect 12817 13481 12851 13515
rect 14013 13481 14047 13515
rect 16589 13481 16623 13515
rect 18061 13481 18095 13515
rect 18521 13481 18555 13515
rect 19809 13481 19843 13515
rect 21189 13481 21223 13515
rect 2558 13413 2592 13447
rect 4077 13413 4111 13447
rect 8723 13413 8757 13447
rect 11161 13413 11195 13447
rect 13185 13413 13219 13447
rect 13737 13413 13771 13447
rect 17462 13413 17496 13447
rect 19165 13413 19199 13447
rect 21833 13413 21867 13447
rect 3617 13345 3651 13379
rect 4169 13345 4203 13379
rect 6101 13345 6135 13379
rect 6561 13345 6595 13379
rect 7113 13345 7147 13379
rect 7389 13345 7423 13379
rect 8636 13345 8670 13379
rect 9965 13345 9999 13379
rect 15577 13345 15611 13379
rect 16037 13345 16071 13379
rect 23616 13345 23650 13379
rect 2237 13277 2271 13311
rect 11069 13277 11103 13311
rect 13093 13277 13127 13311
rect 16313 13277 16347 13311
rect 17141 13277 17175 13311
rect 18889 13277 18923 13311
rect 21741 13277 21775 13311
rect 22017 13277 22051 13311
rect 1685 13209 1719 13243
rect 11621 13209 11655 13243
rect 2053 13141 2087 13175
rect 5181 13141 5215 13175
rect 5457 13141 5491 13175
rect 7849 13141 7883 13175
rect 10103 13141 10137 13175
rect 20085 13141 20119 13175
rect 23719 13141 23753 13175
rect 3157 12937 3191 12971
rect 5457 12937 5491 12971
rect 11529 12937 11563 12971
rect 11805 12937 11839 12971
rect 12633 12937 12667 12971
rect 13093 12937 13127 12971
rect 15577 12937 15611 12971
rect 17877 12937 17911 12971
rect 22293 12937 22327 12971
rect 23397 12937 23431 12971
rect 7297 12869 7331 12903
rect 8861 12869 8895 12903
rect 9689 12869 9723 12903
rect 16037 12869 16071 12903
rect 17141 12869 17175 12903
rect 23811 12869 23845 12903
rect 1685 12801 1719 12835
rect 2329 12801 2363 12835
rect 3341 12801 3375 12835
rect 9321 12801 9355 12835
rect 10609 12801 10643 12835
rect 13645 12801 13679 12835
rect 14565 12801 14599 12835
rect 16221 12801 16255 12835
rect 18889 12801 18923 12835
rect 20085 12801 20119 12835
rect 20821 12801 20855 12835
rect 21373 12801 21407 12835
rect 21649 12801 21683 12835
rect 1777 12665 1811 12699
rect 3617 12733 3651 12767
rect 4261 12733 4295 12767
rect 4445 12733 4479 12767
rect 4997 12733 5031 12767
rect 7481 12733 7515 12767
rect 8125 12733 8159 12767
rect 8309 12733 8343 12767
rect 8861 12733 8895 12767
rect 12449 12733 12483 12767
rect 15025 12733 15059 12767
rect 23740 12733 23774 12767
rect 24133 12733 24167 12767
rect 6193 12665 6227 12699
rect 10930 12665 10964 12699
rect 13461 12665 13495 12699
rect 13737 12665 13771 12699
rect 14289 12665 14323 12699
rect 15117 12665 15151 12699
rect 16542 12665 16576 12699
rect 17417 12665 17451 12699
rect 18245 12665 18279 12699
rect 18337 12665 18371 12699
rect 19809 12665 19843 12699
rect 19901 12665 19935 12699
rect 21189 12665 21223 12699
rect 21465 12665 21499 12699
rect 2605 12597 2639 12631
rect 3341 12597 3375 12631
rect 3433 12597 3467 12631
rect 3709 12597 3743 12631
rect 5733 12597 5767 12631
rect 6561 12597 6595 12631
rect 10057 12597 10091 12631
rect 10517 12597 10551 12631
rect 12173 12597 12207 12631
rect 19165 12597 19199 12631
rect 19533 12597 19567 12631
rect 1593 12393 1627 12427
rect 2421 12393 2455 12427
rect 3341 12393 3375 12427
rect 9505 12393 9539 12427
rect 11529 12393 11563 12427
rect 13093 12393 13127 12427
rect 15439 12393 15473 12427
rect 16221 12393 16255 12427
rect 17693 12393 17727 12427
rect 18245 12393 18279 12427
rect 19257 12393 19291 12427
rect 20085 12393 20119 12427
rect 21741 12393 21775 12427
rect 3709 12325 3743 12359
rect 6469 12325 6503 12359
rect 10654 12325 10688 12359
rect 12817 12325 12851 12359
rect 13829 12325 13863 12359
rect 17094 12325 17128 12359
rect 22109 12325 22143 12359
rect 1409 12257 1443 12291
rect 4997 12257 5031 12291
rect 5457 12257 5491 12291
rect 5825 12257 5859 12291
rect 6285 12257 6319 12291
rect 7297 12257 7331 12291
rect 8033 12257 8067 12291
rect 8309 12257 8343 12291
rect 8677 12257 8711 12291
rect 11253 12257 11287 12291
rect 12725 12257 12759 12291
rect 15336 12257 15370 12291
rect 16773 12257 16807 12291
rect 18521 12257 18555 12291
rect 20821 12257 20855 12291
rect 24568 12257 24602 12291
rect 2053 12189 2087 12223
rect 2513 12189 2547 12223
rect 7205 12189 7239 12223
rect 8769 12189 8803 12223
rect 10333 12189 10367 12223
rect 13737 12189 13771 12223
rect 18889 12189 18923 12223
rect 22017 12189 22051 12223
rect 22661 12189 22695 12223
rect 23489 12189 23523 12223
rect 14289 12121 14323 12155
rect 4537 12053 4571 12087
rect 4905 12053 4939 12087
rect 6745 12053 6779 12087
rect 9045 12053 9079 12087
rect 9873 12053 9907 12087
rect 13553 12053 13587 12087
rect 15853 12053 15887 12087
rect 19809 12053 19843 12087
rect 21051 12053 21085 12087
rect 24639 12053 24673 12087
rect 6285 11849 6319 11883
rect 6653 11849 6687 11883
rect 7849 11849 7883 11883
rect 10885 11849 10919 11883
rect 12265 11849 12299 11883
rect 13829 11849 13863 11883
rect 14289 11849 14323 11883
rect 15301 11849 15335 11883
rect 16773 11849 16807 11883
rect 17141 11849 17175 11883
rect 21465 11849 21499 11883
rect 23029 11849 23063 11883
rect 24685 11849 24719 11883
rect 11897 11781 11931 11815
rect 17785 11781 17819 11815
rect 19625 11781 19659 11815
rect 20913 11781 20947 11815
rect 1501 11713 1535 11747
rect 3617 11713 3651 11747
rect 4353 11713 4387 11747
rect 5917 11713 5951 11747
rect 8677 11713 8711 11747
rect 10057 11713 10091 11747
rect 12909 11713 12943 11747
rect 19901 11713 19935 11747
rect 22109 11713 22143 11747
rect 3249 11645 3283 11679
rect 4445 11645 4479 11679
rect 5181 11645 5215 11679
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 8125 11645 8159 11679
rect 8401 11645 8435 11679
rect 8953 11645 8987 11679
rect 11412 11645 11446 11679
rect 14473 11645 14507 11679
rect 14933 11645 14967 11679
rect 15761 11645 15795 11679
rect 15945 11645 15979 11679
rect 18061 11645 18095 11679
rect 24200 11645 24234 11679
rect 1593 11577 1627 11611
rect 2145 11577 2179 11611
rect 2973 11577 3007 11611
rect 3065 11577 3099 11611
rect 3985 11577 4019 11611
rect 9597 11577 9631 11611
rect 9689 11577 9723 11611
rect 13001 11577 13035 11611
rect 13553 11577 13587 11611
rect 16221 11577 16255 11611
rect 18382 11577 18416 11611
rect 19257 11577 19291 11611
rect 19993 11577 20027 11611
rect 20545 11577 20579 11611
rect 22201 11577 22235 11611
rect 22753 11577 22787 11611
rect 2421 11509 2455 11543
rect 6929 11509 6963 11543
rect 7389 11509 7423 11543
rect 9321 11509 9355 11543
rect 10517 11509 10551 11543
rect 11483 11509 11517 11543
rect 12633 11509 12667 11543
rect 14657 11509 14691 11543
rect 18981 11509 19015 11543
rect 21925 11509 21959 11543
rect 24271 11509 24305 11543
rect 24961 11509 24995 11543
rect 3157 11305 3191 11339
rect 3433 11305 3467 11339
rect 3893 11305 3927 11339
rect 4353 11305 4387 11339
rect 5733 11305 5767 11339
rect 5917 11305 5951 11339
rect 6469 11305 6503 11339
rect 8493 11305 8527 11339
rect 12081 11305 12115 11339
rect 15577 11305 15611 11339
rect 20361 11305 20395 11339
rect 22109 11305 22143 11339
rect 1771 11237 1805 11271
rect 9781 11237 9815 11271
rect 9873 11237 9907 11271
rect 12357 11237 12391 11271
rect 12449 11237 12483 11271
rect 17094 11237 17128 11271
rect 19073 11237 19107 11271
rect 21097 11237 21131 11271
rect 22477 11237 22511 11271
rect 1409 11169 1443 11203
rect 2789 11169 2823 11203
rect 4169 11169 4203 11203
rect 4537 11169 4571 11203
rect 4905 11169 4939 11203
rect 5457 11169 5491 11203
rect 5641 11169 5675 11203
rect 5733 11169 5767 11203
rect 6377 11169 6411 11203
rect 6837 11169 6871 11203
rect 7205 11169 7239 11203
rect 7573 11169 7607 11203
rect 11320 11169 11354 11203
rect 13829 11169 13863 11203
rect 15669 11169 15703 11203
rect 22569 11169 22603 11203
rect 24593 11169 24627 11203
rect 9229 11101 9263 11135
rect 10057 11101 10091 11135
rect 11805 11101 11839 11135
rect 13967 11101 14001 11135
rect 16773 11101 16807 11135
rect 18981 11101 19015 11135
rect 19349 11101 19383 11135
rect 21005 11101 21039 11135
rect 5641 11033 5675 11067
rect 6285 11033 6319 11067
rect 8861 11033 8895 11067
rect 12909 11033 12943 11067
rect 21557 11033 21591 11067
rect 24777 11033 24811 11067
rect 2329 10965 2363 10999
rect 8217 10965 8251 10999
rect 10793 10965 10827 10999
rect 11391 10965 11425 10999
rect 13277 10965 13311 10999
rect 14289 10965 14323 10999
rect 15899 10965 15933 10999
rect 17693 10965 17727 10999
rect 18061 10965 18095 10999
rect 19901 10965 19935 10999
rect 3341 10761 3375 10795
rect 4169 10761 4203 10795
rect 6285 10761 6319 10795
rect 10609 10761 10643 10795
rect 20361 10761 20395 10795
rect 21557 10761 21591 10795
rect 22569 10761 22603 10795
rect 24685 10761 24719 10795
rect 17049 10693 17083 10727
rect 19625 10693 19659 10727
rect 20085 10693 20119 10727
rect 22017 10693 22051 10727
rect 1501 10625 1535 10659
rect 2145 10625 2179 10659
rect 12541 10625 12575 10659
rect 16497 10625 16531 10659
rect 17785 10625 17819 10659
rect 18889 10625 18923 10659
rect 22109 10625 22143 10659
rect 3249 10557 3283 10591
rect 4445 10557 4479 10591
rect 4997 10557 5031 10591
rect 5273 10557 5307 10591
rect 5825 10557 5859 10591
rect 6561 10557 6595 10591
rect 7113 10557 7147 10591
rect 7573 10557 7607 10591
rect 7941 10557 7975 10591
rect 8493 10557 8527 10591
rect 8585 10557 8619 10591
rect 9413 10557 9447 10591
rect 11228 10557 11262 10591
rect 11621 10557 11655 10591
rect 14013 10557 14047 10591
rect 21281 10557 21315 10591
rect 23740 10557 23774 10591
rect 24133 10557 24167 10591
rect 1593 10489 1627 10523
rect 3065 10489 3099 10523
rect 9321 10489 9355 10523
rect 9734 10489 9768 10523
rect 12633 10489 12667 10523
rect 13185 10489 13219 10523
rect 14334 10489 14368 10523
rect 15761 10489 15795 10523
rect 16313 10489 16347 10523
rect 16589 10489 16623 10523
rect 19073 10489 19107 10523
rect 19165 10489 19199 10523
rect 20637 10489 20671 10523
rect 20729 10489 20763 10523
rect 2421 10421 2455 10455
rect 2973 10421 3007 10455
rect 5641 10421 5675 10455
rect 8861 10421 8895 10455
rect 10333 10421 10367 10455
rect 11299 10421 11333 10455
rect 11989 10421 12023 10455
rect 13461 10421 13495 10455
rect 13829 10421 13863 10455
rect 14933 10421 14967 10455
rect 17417 10421 17451 10455
rect 18521 10421 18555 10455
rect 23811 10421 23845 10455
rect 1869 10217 1903 10251
rect 3157 10217 3191 10251
rect 3525 10217 3559 10251
rect 4261 10217 4295 10251
rect 6561 10217 6595 10251
rect 8033 10217 8067 10251
rect 9045 10217 9079 10251
rect 9413 10217 9447 10251
rect 9873 10217 9907 10251
rect 16497 10217 16531 10251
rect 21005 10217 21039 10251
rect 23719 10217 23753 10251
rect 2881 10149 2915 10183
rect 5825 10149 5859 10183
rect 2053 10081 2087 10115
rect 2973 10081 3007 10115
rect 4077 10081 4111 10115
rect 4537 10081 4571 10115
rect 5273 10081 5307 10115
rect 8769 10149 8803 10183
rect 11206 10149 11240 10183
rect 12817 10149 12851 10183
rect 13369 10149 13403 10183
rect 15485 10149 15519 10183
rect 17186 10149 17220 10183
rect 18981 10149 19015 10183
rect 6653 10081 6687 10115
rect 6929 10081 6963 10115
rect 8217 10081 8251 10115
rect 8401 10081 8435 10115
rect 9689 10081 9723 10115
rect 11805 10081 11839 10115
rect 12081 10081 12115 10115
rect 14197 10081 14231 10115
rect 16865 10081 16899 10115
rect 20913 10081 20947 10115
rect 21373 10081 21407 10115
rect 23581 10081 23615 10115
rect 24593 10081 24627 10115
rect 7389 10013 7423 10047
rect 10885 10013 10919 10047
rect 12725 10013 12759 10047
rect 15393 10013 15427 10047
rect 16037 10013 16071 10047
rect 18705 10013 18739 10047
rect 18889 10013 18923 10047
rect 19349 10013 19383 10047
rect 6377 9945 6411 9979
rect 6561 9945 6595 9979
rect 6745 9945 6779 9979
rect 7665 9945 7699 9979
rect 14381 9945 14415 9979
rect 2421 9877 2455 9911
rect 3893 9877 3927 9911
rect 4905 9877 4939 9911
rect 12449 9877 12483 9911
rect 14013 9877 14047 9911
rect 17785 9877 17819 9911
rect 18153 9877 18187 9911
rect 19901 9877 19935 9911
rect 20637 9877 20671 9911
rect 24777 9877 24811 9911
rect 5365 9673 5399 9707
rect 5917 9673 5951 9707
rect 6653 9673 6687 9707
rect 8953 9673 8987 9707
rect 15117 9673 15151 9707
rect 15485 9673 15519 9707
rect 15761 9673 15795 9707
rect 16957 9673 16991 9707
rect 17325 9673 17359 9707
rect 17785 9673 17819 9707
rect 19165 9673 19199 9707
rect 21327 9673 21361 9707
rect 24685 9673 24719 9707
rect 2053 9605 2087 9639
rect 6285 9605 6319 9639
rect 8585 9605 8619 9639
rect 16589 9605 16623 9639
rect 23857 9605 23891 9639
rect 9689 9537 9723 9571
rect 11161 9537 11195 9571
rect 11621 9537 11655 9571
rect 18797 9537 18831 9571
rect 3525 9469 3559 9503
rect 3985 9469 4019 9503
rect 4353 9469 4387 9503
rect 4905 9469 4939 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 7849 9469 7883 9503
rect 8217 9469 8251 9503
rect 9321 9469 9355 9503
rect 9965 9469 9999 9503
rect 10885 9469 10919 9503
rect 11069 9469 11103 9503
rect 12725 9469 12759 9503
rect 13001 9469 13035 9503
rect 14197 9469 14231 9503
rect 19533 9469 19567 9503
rect 19625 9469 19659 9503
rect 20085 9469 20119 9503
rect 21256 9469 21290 9503
rect 1501 9401 1535 9435
rect 1593 9401 1627 9435
rect 9137 9401 9171 9435
rect 10517 9401 10551 9435
rect 12265 9401 12299 9435
rect 14013 9401 14047 9435
rect 14518 9401 14552 9435
rect 16037 9401 16071 9435
rect 16129 9401 16163 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 20913 9401 20947 9435
rect 2421 9333 2455 9367
rect 3065 9333 3099 9367
rect 3433 9333 3467 9367
rect 3617 9333 3651 9367
rect 7113 9333 7147 9367
rect 12541 9333 12575 9367
rect 13461 9333 13495 9367
rect 19717 9333 19751 9367
rect 21649 9333 21683 9367
rect 2697 9129 2731 9163
rect 4629 9129 4663 9163
rect 1771 9061 1805 9095
rect 1409 8993 1443 9027
rect 4353 8993 4387 9027
rect 4629 8993 4663 9027
rect 4721 9129 4755 9163
rect 6469 9129 6503 9163
rect 7297 9129 7331 9163
rect 9137 9129 9171 9163
rect 9873 9129 9907 9163
rect 11069 9129 11103 9163
rect 16313 9129 16347 9163
rect 21051 9129 21085 9163
rect 21373 9129 21407 9163
rect 7665 9061 7699 9095
rect 11523 9061 11557 9095
rect 13093 9061 13127 9095
rect 15025 9061 15059 9095
rect 15485 9061 15519 9095
rect 17601 9061 17635 9095
rect 5181 8993 5215 9027
rect 5365 8993 5399 9027
rect 5641 8993 5675 9027
rect 8217 8993 8251 9027
rect 9689 8993 9723 9027
rect 11161 8993 11195 9027
rect 12081 8993 12115 9027
rect 14197 8993 14231 9027
rect 16037 8993 16071 9027
rect 17141 8993 17175 9027
rect 17325 8993 17359 9027
rect 18613 8993 18647 9027
rect 18889 8993 18923 9027
rect 20948 8993 20982 9027
rect 4721 8925 4755 8959
rect 5825 8925 5859 8959
rect 8585 8925 8619 8959
rect 10701 8925 10735 8959
rect 13001 8925 13035 8959
rect 13277 8925 13311 8959
rect 15393 8925 15427 8959
rect 18981 8925 19015 8959
rect 5457 8857 5491 8891
rect 2329 8789 2363 8823
rect 2973 8789 3007 8823
rect 3617 8789 3651 8823
rect 4537 8789 4571 8823
rect 4813 8789 4847 8823
rect 6837 8789 6871 8823
rect 10149 8789 10183 8823
rect 12541 8789 12575 8823
rect 14657 8789 14691 8823
rect 18153 8789 18187 8823
rect 19625 8789 19659 8823
rect 2789 8585 2823 8619
rect 4353 8585 4387 8619
rect 5549 8585 5583 8619
rect 6009 8585 6043 8619
rect 11805 8585 11839 8619
rect 13461 8585 13495 8619
rect 14933 8585 14967 8619
rect 15301 8585 15335 8619
rect 17325 8585 17359 8619
rect 17877 8585 17911 8619
rect 19073 8585 19107 8619
rect 24777 8585 24811 8619
rect 2053 8517 2087 8551
rect 3065 8517 3099 8551
rect 18705 8517 18739 8551
rect 3709 8449 3743 8483
rect 9137 8449 9171 8483
rect 10333 8449 10367 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 13829 8449 13863 8483
rect 16497 8449 16531 8483
rect 18153 8449 18187 8483
rect 21327 8449 21361 8483
rect 2973 8381 3007 8415
rect 3249 8381 3283 8415
rect 4261 8381 4295 8415
rect 4537 8381 4571 8415
rect 4629 8381 4663 8415
rect 4813 8381 4847 8415
rect 6837 8381 6871 8415
rect 6929 8381 6963 8415
rect 7113 8381 7147 8415
rect 8401 8381 8435 8415
rect 8493 8381 8527 8415
rect 8677 8381 8711 8415
rect 12265 8381 12299 8415
rect 12725 8381 12759 8415
rect 13001 8381 13035 8415
rect 14013 8381 14047 8415
rect 16313 8381 16347 8415
rect 19625 8381 19659 8415
rect 20085 8381 20119 8415
rect 21224 8381 21258 8415
rect 21649 8381 21683 8415
rect 24593 8381 24627 8415
rect 25145 8381 25179 8415
rect 1501 8313 1535 8347
rect 1593 8313 1627 8347
rect 2513 8313 2547 8347
rect 10701 8313 10735 8347
rect 10977 8313 11011 8347
rect 14334 8313 14368 8347
rect 15669 8313 15703 8347
rect 18245 8313 18279 8347
rect 19441 8313 19475 8347
rect 3985 8245 4019 8279
rect 4261 8245 4295 8279
rect 4997 8245 5031 8279
rect 6561 8245 6595 8279
rect 7297 8245 7331 8279
rect 7941 8245 7975 8279
rect 8217 8245 8251 8279
rect 9781 8245 9815 8279
rect 12541 8245 12575 8279
rect 16957 8245 16991 8279
rect 19717 8245 19751 8279
rect 20913 8245 20947 8279
rect 1593 8041 1627 8075
rect 2881 8041 2915 8075
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 9137 8041 9171 8075
rect 10149 8041 10183 8075
rect 11161 8041 11195 8075
rect 11713 8041 11747 8075
rect 13001 8041 13035 8075
rect 14657 8041 14691 8075
rect 19947 8041 19981 8075
rect 21097 8041 21131 8075
rect 2329 7973 2363 8007
rect 12167 7973 12201 8007
rect 13737 7973 13771 8007
rect 15853 7973 15887 8007
rect 16818 7973 16852 8007
rect 18429 7973 18463 8007
rect 1409 7905 1443 7939
rect 2973 7905 3007 7939
rect 3801 7905 3835 7939
rect 4169 7905 4203 7939
rect 5825 7905 5859 7939
rect 7297 7905 7331 7939
rect 7573 7905 7607 7939
rect 8493 7905 8527 7939
rect 9689 7905 9723 7939
rect 9781 7905 9815 7939
rect 9965 7905 9999 7939
rect 11805 7905 11839 7939
rect 12725 7905 12759 7939
rect 15301 7905 15335 7939
rect 16497 7905 16531 7939
rect 19876 7905 19910 7939
rect 20913 7905 20947 7939
rect 4077 7837 4111 7871
rect 6469 7837 6503 7871
rect 7757 7837 7791 7871
rect 13645 7837 13679 7871
rect 14289 7837 14323 7871
rect 16129 7837 16163 7871
rect 18337 7837 18371 7871
rect 18981 7837 19015 7871
rect 7389 7769 7423 7803
rect 19625 7769 19659 7803
rect 1961 7701 1995 7735
rect 3433 7701 3467 7735
rect 6929 7701 6963 7735
rect 8769 7701 8803 7735
rect 10885 7701 10919 7735
rect 15485 7701 15519 7735
rect 17417 7701 17451 7735
rect 18153 7701 18187 7735
rect 1685 7497 1719 7531
rect 4169 7497 4203 7531
rect 5273 7497 5307 7531
rect 5825 7497 5859 7531
rect 7205 7497 7239 7531
rect 8769 7497 8803 7531
rect 10333 7497 10367 7531
rect 11897 7497 11931 7531
rect 13645 7497 13679 7531
rect 19349 7497 19383 7531
rect 21465 7497 21499 7531
rect 3065 7429 3099 7463
rect 9045 7429 9079 7463
rect 14657 7429 14691 7463
rect 17049 7429 17083 7463
rect 19073 7429 19107 7463
rect 3617 7361 3651 7395
rect 9689 7361 9723 7395
rect 12541 7361 12575 7395
rect 13185 7361 13219 7395
rect 14105 7361 14139 7395
rect 15301 7361 15335 7395
rect 16497 7361 16531 7395
rect 20775 7361 20809 7395
rect 2053 7293 2087 7327
rect 2973 7293 3007 7327
rect 3249 7293 3283 7327
rect 4721 7293 4755 7327
rect 4905 7293 4939 7327
rect 7665 7293 7699 7327
rect 7849 7293 7883 7327
rect 8953 7293 8987 7327
rect 9229 7293 9263 7327
rect 9965 7293 9999 7327
rect 11069 7293 11103 7327
rect 11345 7293 11379 7327
rect 17509 7293 17543 7327
rect 19349 7293 19383 7327
rect 19625 7293 19659 7327
rect 20672 7293 20706 7327
rect 21097 7293 21131 7327
rect 11529 7225 11563 7259
rect 12633 7225 12667 7259
rect 14197 7225 14231 7259
rect 16221 7225 16255 7259
rect 16589 7225 16623 7259
rect 17785 7225 17819 7259
rect 18153 7225 18187 7259
rect 18245 7225 18279 7259
rect 18797 7225 18831 7259
rect 2513 7157 2547 7191
rect 2881 7157 2915 7191
rect 6561 7157 6595 7191
rect 7665 7157 7699 7191
rect 8401 7157 8435 7191
rect 12265 7157 12299 7191
rect 15853 7157 15887 7191
rect 19441 7157 19475 7191
rect 20177 7157 20211 7191
rect 3801 6953 3835 6987
rect 5273 6953 5307 6987
rect 7297 6953 7331 6987
rect 9413 6953 9447 6987
rect 9781 6953 9815 6987
rect 10885 6953 10919 6987
rect 14105 6953 14139 6987
rect 14473 6953 14507 6987
rect 16681 6953 16715 6987
rect 19855 6953 19889 6987
rect 2145 6885 2179 6919
rect 2789 6885 2823 6919
rect 3433 6885 3467 6919
rect 6561 6885 6595 6919
rect 15806 6885 15840 6919
rect 18337 6885 18371 6919
rect 1593 6817 1627 6851
rect 3008 6817 3042 6851
rect 4813 6817 4847 6851
rect 6193 6817 6227 6851
rect 7389 6817 7423 6851
rect 7849 6817 7883 6851
rect 9965 6817 9999 6851
rect 10149 6817 10183 6851
rect 11805 6817 11839 6851
rect 11989 6817 12023 6851
rect 12541 6817 12575 6851
rect 13369 6817 13403 6851
rect 13553 6817 13587 6851
rect 19752 6817 19786 6851
rect 24593 6817 24627 6851
rect 4261 6749 4295 6783
rect 7113 6749 7147 6783
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 12081 6749 12115 6783
rect 13645 6749 13679 6783
rect 15485 6749 15519 6783
rect 18245 6749 18279 6783
rect 3111 6681 3145 6715
rect 14933 6681 14967 6715
rect 18061 6681 18095 6715
rect 18797 6681 18831 6715
rect 4997 6613 5031 6647
rect 6837 6613 6871 6647
rect 7113 6613 7147 6647
rect 8953 6613 8987 6647
rect 13001 6613 13035 6647
rect 16405 6613 16439 6647
rect 24731 6613 24765 6647
rect 4077 6409 4111 6443
rect 5365 6409 5399 6443
rect 5641 6409 5675 6443
rect 6653 6409 6687 6443
rect 9045 6409 9079 6443
rect 10609 6409 10643 6443
rect 17141 6409 17175 6443
rect 19257 6409 19291 6443
rect 19947 6409 19981 6443
rect 20361 6409 20395 6443
rect 1869 6341 1903 6375
rect 2605 6273 2639 6307
rect 3157 6273 3191 6307
rect 3709 6273 3743 6307
rect 4629 6273 4663 6307
rect 5273 6273 5307 6307
rect 1685 6205 1719 6239
rect 2697 6205 2731 6239
rect 2789 6205 2823 6239
rect 2973 6205 3007 6239
rect 7021 6341 7055 6375
rect 9505 6341 9539 6375
rect 11345 6341 11379 6375
rect 7849 6273 7883 6307
rect 9689 6273 9723 6307
rect 10149 6273 10183 6307
rect 11713 6273 11747 6307
rect 14197 6273 14231 6307
rect 18613 6273 18647 6307
rect 19625 6273 19659 6307
rect 5733 6205 5767 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 11161 6205 11195 6239
rect 12265 6205 12299 6239
rect 12725 6205 12759 6239
rect 12909 6205 12943 6239
rect 13829 6205 13863 6239
rect 14381 6205 14415 6239
rect 14841 6205 14875 6239
rect 15117 6205 15151 6239
rect 15945 6205 15979 6239
rect 19876 6205 19910 6239
rect 6193 6137 6227 6171
rect 8170 6137 8204 6171
rect 9781 6137 9815 6171
rect 10977 6137 11011 6171
rect 16266 6137 16300 6171
rect 17877 6137 17911 6171
rect 18337 6137 18371 6171
rect 18429 6137 18463 6171
rect 2145 6069 2179 6103
rect 4859 6069 4893 6103
rect 5365 6069 5399 6103
rect 5917 6069 5951 6103
rect 7757 6069 7791 6103
rect 8769 6069 8803 6103
rect 12541 6069 12575 6103
rect 13461 6069 13495 6103
rect 15485 6069 15519 6103
rect 15761 6069 15795 6103
rect 16865 6069 16899 6103
rect 24685 6069 24719 6103
rect 1685 5865 1719 5899
rect 1961 5865 1995 5899
rect 2329 5865 2363 5899
rect 2789 5865 2823 5899
rect 3157 5865 3191 5899
rect 4261 5865 4295 5899
rect 5089 5865 5123 5899
rect 7389 5865 7423 5899
rect 8769 5865 8803 5899
rect 11621 5865 11655 5899
rect 13967 5865 14001 5899
rect 14473 5865 14507 5899
rect 16497 5865 16531 5899
rect 18245 5865 18279 5899
rect 5502 5797 5536 5831
rect 8170 5797 8204 5831
rect 9413 5797 9447 5831
rect 9873 5797 9907 5831
rect 12402 5797 12436 5831
rect 15669 5797 15703 5831
rect 17370 5797 17404 5831
rect 18981 5797 19015 5831
rect 19533 5797 19567 5831
rect 1476 5729 1510 5763
rect 2973 5729 3007 5763
rect 4077 5729 4111 5763
rect 5181 5729 5215 5763
rect 7849 5729 7883 5763
rect 9045 5729 9079 5763
rect 12081 5729 12115 5763
rect 13829 5729 13863 5763
rect 16221 5729 16255 5763
rect 9781 5661 9815 5695
rect 10149 5661 10183 5695
rect 15577 5661 15611 5695
rect 17049 5661 17083 5695
rect 18889 5661 18923 5695
rect 13001 5593 13035 5627
rect 17969 5593 18003 5627
rect 6101 5525 6135 5559
rect 6929 5525 6963 5559
rect 14749 5525 14783 5559
rect 18613 5525 18647 5559
rect 1547 5321 1581 5355
rect 2237 5321 2271 5355
rect 3801 5321 3835 5355
rect 8217 5321 8251 5355
rect 10885 5321 10919 5355
rect 11437 5321 11471 5355
rect 13829 5321 13863 5355
rect 15393 5321 15427 5355
rect 19809 5321 19843 5355
rect 20131 5321 20165 5355
rect 3157 5253 3191 5287
rect 4721 5253 4755 5287
rect 6193 5253 6227 5287
rect 7849 5253 7883 5287
rect 9505 5253 9539 5287
rect 12173 5253 12207 5287
rect 20545 5253 20579 5287
rect 4537 5185 4571 5219
rect 1444 5117 1478 5151
rect 1869 5117 1903 5151
rect 2973 5117 3007 5151
rect 4020 5117 4054 5151
rect 6929 5185 6963 5219
rect 8677 5185 8711 5219
rect 9689 5185 9723 5219
rect 12817 5185 12851 5219
rect 14105 5185 14139 5219
rect 18797 5185 18831 5219
rect 4997 5117 5031 5151
rect 8468 5117 8502 5151
rect 10609 5117 10643 5151
rect 12265 5117 12299 5151
rect 15117 5117 15151 5151
rect 15945 5117 15979 5151
rect 20060 5117 20094 5151
rect 4721 5049 4755 5083
rect 4813 5049 4847 5083
rect 5338 5049 5372 5083
rect 6561 5049 6595 5083
rect 7014 5049 7048 5083
rect 7573 5049 7607 5083
rect 10010 5049 10044 5083
rect 12541 5049 12575 5083
rect 12633 5049 12667 5083
rect 13461 5049 13495 5083
rect 14197 5049 14231 5083
rect 14749 5049 14783 5083
rect 16266 5049 16300 5083
rect 17141 5049 17175 5083
rect 18521 5049 18555 5083
rect 18613 5049 18647 5083
rect 3433 4981 3467 5015
rect 4123 4981 4157 5015
rect 5917 4981 5951 5015
rect 8953 4981 8987 5015
rect 11713 4981 11747 5015
rect 12265 4981 12299 5015
rect 15761 4981 15795 5015
rect 16865 4981 16899 5015
rect 17601 4981 17635 5015
rect 18337 4981 18371 5015
rect 19441 4981 19475 5015
rect 1547 4777 1581 4811
rect 4353 4777 4387 4811
rect 5825 4777 5859 4811
rect 7481 4777 7515 4811
rect 10241 4777 10275 4811
rect 12173 4777 12207 4811
rect 12633 4777 12667 4811
rect 14473 4777 14507 4811
rect 15117 4777 15151 4811
rect 18521 4777 18555 4811
rect 5549 4709 5583 4743
rect 6561 4709 6595 4743
rect 7113 4709 7147 4743
rect 9873 4709 9907 4743
rect 10609 4709 10643 4743
rect 15714 4709 15748 4743
rect 17509 4709 17543 4743
rect 18889 4709 18923 4743
rect 1476 4641 1510 4675
rect 4905 4641 4939 4675
rect 8033 4641 8067 4675
rect 8309 4641 8343 4675
rect 8769 4641 8803 4675
rect 12265 4641 12299 4675
rect 14013 4641 14047 4675
rect 6469 4573 6503 4607
rect 10517 4573 10551 4607
rect 10793 4573 10827 4607
rect 15393 4573 15427 4607
rect 17417 4573 17451 4607
rect 17693 4573 17727 4607
rect 8125 4505 8159 4539
rect 13185 4505 13219 4539
rect 14151 4437 14185 4471
rect 16313 4437 16347 4471
rect 1685 4233 1719 4267
rect 4905 4233 4939 4267
rect 6469 4233 6503 4267
rect 9229 4233 9263 4267
rect 10793 4233 10827 4267
rect 12265 4233 12299 4267
rect 13645 4233 13679 4267
rect 16313 4233 16347 4267
rect 17417 4233 17451 4267
rect 17785 4233 17819 4267
rect 8769 4165 8803 4199
rect 15761 4165 15795 4199
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 8401 4097 8435 4131
rect 9413 4097 9447 4131
rect 12449 4097 12483 4131
rect 16497 4097 16531 4131
rect 17141 4097 17175 4131
rect 18429 4097 18463 4131
rect 24731 4097 24765 4131
rect 5825 4029 5859 4063
rect 11412 4029 11446 4063
rect 11805 4029 11839 4063
rect 24644 4029 24678 4063
rect 5917 3961 5951 3995
rect 7021 3961 7055 3995
rect 9505 3961 9539 3995
rect 10057 3961 10091 3995
rect 11621 3961 11655 3995
rect 12770 3961 12804 3995
rect 14289 3961 14323 3995
rect 14381 3961 14415 3995
rect 14933 3961 14967 3995
rect 16589 3961 16623 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 8125 3893 8159 3927
rect 10517 3893 10551 3927
rect 13369 3893 13403 3927
rect 14013 3893 14047 3927
rect 15393 3893 15427 3927
rect 25145 3893 25179 3927
rect 5273 3689 5307 3723
rect 5503 3689 5537 3723
rect 5825 3689 5859 3723
rect 7389 3689 7423 3723
rect 9413 3689 9447 3723
rect 12541 3689 12575 3723
rect 14289 3689 14323 3723
rect 15025 3689 15059 3723
rect 15393 3689 15427 3723
rect 16497 3689 16531 3723
rect 17969 3689 18003 3723
rect 18245 3689 18279 3723
rect 6561 3621 6595 3655
rect 7113 3621 7147 3655
rect 8217 3621 8251 3655
rect 9873 3621 9907 3655
rect 10425 3621 10459 3655
rect 11437 3621 11471 3655
rect 11989 3621 12023 3655
rect 12909 3621 12943 3655
rect 13001 3621 13035 3655
rect 13553 3621 13587 3655
rect 17601 3621 17635 3655
rect 1476 3553 1510 3587
rect 5365 3553 5399 3587
rect 8769 3553 8803 3587
rect 14565 3553 14599 3587
rect 15577 3553 15611 3587
rect 15761 3553 15795 3587
rect 17141 3553 17175 3587
rect 17325 3553 17359 3587
rect 18429 3553 18463 3587
rect 4353 3485 4387 3519
rect 6469 3485 6503 3519
rect 8125 3485 8159 3519
rect 9781 3485 9815 3519
rect 11345 3485 11379 3519
rect 1547 3417 1581 3451
rect 7757 3417 7791 3451
rect 6285 3349 6319 3383
rect 10701 3349 10735 3383
rect 18567 3349 18601 3383
rect 1869 3145 1903 3179
rect 5365 3145 5399 3179
rect 6469 3145 6503 3179
rect 7021 3145 7055 3179
rect 8861 3145 8895 3179
rect 10333 3145 10367 3179
rect 10701 3145 10735 3179
rect 11437 3145 11471 3179
rect 12173 3145 12207 3179
rect 13093 3145 13127 3179
rect 14841 3145 14875 3179
rect 16037 3145 16071 3179
rect 17141 3145 17175 3179
rect 17509 3145 17543 3179
rect 18429 3145 18463 3179
rect 4859 3077 4893 3111
rect 9965 3077 9999 3111
rect 12633 3077 12667 3111
rect 1547 3009 1581 3043
rect 7849 3009 7883 3043
rect 8493 3009 8527 3043
rect 9413 3009 9447 3043
rect 10885 3009 10919 3043
rect 11713 3009 11747 3043
rect 13369 3009 13403 3043
rect 1444 2941 1478 2975
rect 2237 2941 2271 2975
rect 4629 2941 4663 2975
rect 4756 2941 4790 2975
rect 5800 2941 5834 2975
rect 12449 2941 12483 2975
rect 13921 2941 13955 2975
rect 15025 2941 15059 2975
rect 15485 2941 15519 2975
rect 16405 2941 16439 2975
rect 16589 2941 16623 2975
rect 3847 2873 3881 2907
rect 7665 2873 7699 2907
rect 7941 2873 7975 2907
rect 9505 2873 9539 2907
rect 3617 2805 3651 2839
rect 4261 2805 4295 2839
rect 5871 2805 5905 2839
rect 9229 2805 9263 2839
rect 14105 2805 14139 2839
rect 14565 2805 14599 2839
rect 15301 2805 15335 2839
rect 16773 2805 16807 2839
rect 7297 2601 7331 2635
rect 7757 2601 7791 2635
rect 8769 2601 8803 2635
rect 11483 2601 11517 2635
rect 15669 2601 15703 2635
rect 18475 2601 18509 2635
rect 20223 2601 20257 2635
rect 4721 2533 4755 2567
rect 8170 2533 8204 2567
rect 9597 2533 9631 2567
rect 9965 2533 9999 2567
rect 12633 2533 12667 2567
rect 17509 2533 17543 2567
rect 23121 2533 23155 2567
rect 3040 2465 3074 2499
rect 4512 2465 4546 2499
rect 5733 2465 5767 2499
rect 6285 2465 6319 2499
rect 7849 2465 7883 2499
rect 11412 2465 11446 2499
rect 12449 2465 12483 2499
rect 12725 2465 12759 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15485 2465 15519 2499
rect 16656 2465 16690 2499
rect 17049 2465 17083 2499
rect 18404 2465 18438 2499
rect 20152 2465 20186 2499
rect 22569 2465 22603 2499
rect 9045 2397 9079 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 11805 2397 11839 2431
rect 18889 2397 18923 2431
rect 20637 2397 20671 2431
rect 3111 2329 3145 2363
rect 5917 2329 5951 2363
rect 16129 2329 16163 2363
rect 16727 2329 16761 2363
rect 22753 2329 22787 2363
rect 3525 2261 3559 2295
rect 4905 2261 4939 2295
rect 10793 2261 10827 2295
rect 14381 2261 14415 2295
<< metal1 >>
rect 3050 27480 3056 27532
rect 3108 27520 3114 27532
rect 3878 27520 3884 27532
rect 3108 27492 3884 27520
rect 3108 27480 3114 27492
rect 3878 27480 3884 27492
rect 3936 27480 3942 27532
rect 13906 27480 13912 27532
rect 13964 27520 13970 27532
rect 14550 27520 14556 27532
rect 13964 27492 14556 27520
rect 13964 27480 13970 27492
rect 14550 27480 14556 27492
rect 14608 27480 14614 27532
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 25958 27520 25964 27532
rect 24912 27492 25964 27520
rect 24912 27480 24918 27492
rect 25958 27480 25964 27492
rect 26016 27480 26022 27532
rect 6914 26596 6920 26648
rect 6972 26636 6978 26648
rect 8110 26636 8116 26648
rect 6972 26608 8116 26636
rect 6972 26596 6978 26608
rect 8110 26596 8116 26608
rect 8168 26596 8174 26648
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1464 24259 1522 24265
rect 1464 24225 1476 24259
rect 1510 24256 1522 24259
rect 1854 24256 1860 24268
rect 1510 24228 1860 24256
rect 1510 24225 1522 24228
rect 1464 24219 1522 24225
rect 1854 24216 1860 24228
rect 1912 24216 1918 24268
rect 5994 24216 6000 24268
rect 6052 24256 6058 24268
rect 8332 24259 8390 24265
rect 8332 24256 8344 24259
rect 6052 24228 8344 24256
rect 6052 24216 6058 24228
rect 8332 24225 8344 24228
rect 8378 24256 8390 24259
rect 8754 24256 8760 24268
rect 8378 24228 8760 24256
rect 8378 24225 8390 24228
rect 8332 24219 8390 24225
rect 8754 24216 8760 24228
rect 8812 24216 8818 24268
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 2682 24052 2688 24064
rect 1581 24024 2688 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 8435 24055 8493 24061
rect 8435 24021 8447 24055
rect 8481 24052 8493 24055
rect 9214 24052 9220 24064
rect 8481 24024 9220 24052
rect 8481 24021 8493 24024
rect 8435 24015 8493 24021
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1854 23848 1860 23860
rect 1815 23820 1860 23848
rect 1854 23808 1860 23820
rect 1912 23808 1918 23860
rect 8754 23848 8760 23860
rect 8715 23820 8760 23848
rect 8754 23808 8760 23820
rect 8812 23808 8818 23860
rect 9493 23851 9551 23857
rect 9493 23817 9505 23851
rect 9539 23848 9551 23851
rect 10686 23848 10692 23860
rect 9539 23820 10692 23848
rect 9539 23817 9551 23820
rect 9493 23811 9551 23817
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 14737 23851 14795 23857
rect 14737 23817 14749 23851
rect 14783 23848 14795 23851
rect 15746 23848 15752 23860
rect 14783 23820 15752 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 19889 23851 19947 23857
rect 19889 23817 19901 23851
rect 19935 23848 19947 23851
rect 20898 23848 20904 23860
rect 19935 23820 20904 23848
rect 19935 23817 19947 23820
rect 19889 23811 19947 23817
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21637 23851 21695 23857
rect 21637 23817 21649 23851
rect 21683 23848 21695 23851
rect 23382 23848 23388 23860
rect 21683 23820 23388 23848
rect 21683 23817 21695 23820
rect 21637 23811 21695 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 4338 23672 4344 23724
rect 4396 23712 4402 23724
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 4396 23684 9137 23712
rect 4396 23672 4402 23684
rect 1302 23604 1308 23656
rect 1360 23644 1366 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 1360 23616 1444 23644
rect 1360 23604 1366 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 2225 23647 2283 23653
rect 2225 23644 2237 23647
rect 1478 23616 2237 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 2225 23613 2237 23616
rect 2271 23613 2283 23647
rect 2225 23607 2283 23613
rect 6892 23647 6950 23653
rect 6892 23613 6904 23647
rect 6938 23644 6950 23647
rect 7190 23644 7196 23656
rect 6938 23616 7196 23644
rect 6938 23613 6950 23616
rect 6892 23607 6950 23613
rect 7190 23604 7196 23616
rect 7248 23644 7254 23656
rect 8347 23653 8375 23684
rect 9125 23681 9137 23684
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 7285 23647 7343 23653
rect 7285 23644 7297 23647
rect 7248 23616 7297 23644
rect 7248 23604 7254 23616
rect 7285 23613 7297 23616
rect 7331 23613 7343 23647
rect 7285 23607 7343 23613
rect 8332 23647 8390 23653
rect 8332 23613 8344 23647
rect 8378 23613 8390 23647
rect 8332 23607 8390 23613
rect 9309 23647 9367 23653
rect 9309 23613 9321 23647
rect 9355 23644 9367 23647
rect 9858 23644 9864 23656
rect 9355 23616 9864 23644
rect 9355 23613 9367 23616
rect 9309 23607 9367 23613
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23644 14611 23647
rect 16920 23647 16978 23653
rect 14599 23616 15240 23644
rect 14599 23613 14611 23616
rect 14553 23607 14611 23613
rect 1394 23468 1400 23520
rect 1452 23508 1458 23520
rect 1535 23511 1593 23517
rect 1535 23508 1547 23511
rect 1452 23480 1547 23508
rect 1452 23468 1458 23480
rect 1535 23477 1547 23480
rect 1581 23477 1593 23511
rect 1535 23471 1593 23477
rect 6963 23511 7021 23517
rect 6963 23477 6975 23511
rect 7009 23508 7021 23511
rect 7098 23508 7104 23520
rect 7009 23480 7104 23508
rect 7009 23477 7021 23480
rect 6963 23471 7021 23477
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 8435 23511 8493 23517
rect 8435 23477 8447 23511
rect 8481 23508 8493 23511
rect 8662 23508 8668 23520
rect 8481 23480 8668 23508
rect 8481 23477 8493 23480
rect 8435 23471 8493 23477
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 15212 23517 15240 23616
rect 16920 23613 16932 23647
rect 16966 23644 16978 23647
rect 17402 23644 17408 23656
rect 16966 23616 17408 23644
rect 16966 23613 16978 23616
rect 16920 23607 16978 23613
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 17494 23604 17500 23656
rect 17552 23644 17558 23656
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 17552 23616 19717 23644
rect 17552 23604 17558 23616
rect 19705 23613 19717 23616
rect 19751 23644 19763 23647
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 19751 23616 20269 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 21453 23647 21511 23653
rect 21453 23613 21465 23647
rect 21499 23644 21511 23647
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21499 23616 22017 23644
rect 21499 23613 21511 23616
rect 21453 23607 21511 23613
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 24648 23647 24706 23653
rect 24648 23613 24660 23647
rect 24694 23644 24706 23647
rect 25130 23644 25136 23656
rect 24694 23616 25136 23644
rect 24694 23613 24706 23616
rect 24648 23607 24706 23613
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 21468 23576 21496 23607
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 19484 23548 21496 23576
rect 19484 23536 19490 23548
rect 15197 23511 15255 23517
rect 15197 23477 15209 23511
rect 15243 23508 15255 23511
rect 15286 23508 15292 23520
rect 15243 23480 15292 23508
rect 15243 23477 15255 23480
rect 15197 23471 15255 23477
rect 15286 23468 15292 23480
rect 15344 23468 15350 23520
rect 16482 23468 16488 23520
rect 16540 23508 16546 23520
rect 16991 23511 17049 23517
rect 16991 23508 17003 23511
rect 16540 23480 17003 23508
rect 16540 23468 16546 23480
rect 16991 23477 17003 23480
rect 17037 23477 17049 23511
rect 17402 23508 17408 23520
rect 17363 23480 17408 23508
rect 16991 23471 17049 23477
rect 17402 23468 17408 23480
rect 17460 23468 17466 23520
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 24719 23511 24777 23517
rect 24719 23508 24731 23511
rect 22980 23480 24731 23508
rect 22980 23468 22986 23480
rect 24719 23477 24731 23480
rect 24765 23477 24777 23511
rect 24719 23471 24777 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 9858 23264 9864 23316
rect 9916 23304 9922 23316
rect 10091 23307 10149 23313
rect 10091 23304 10103 23307
rect 9916 23276 10103 23304
rect 9916 23264 9922 23276
rect 10091 23273 10103 23276
rect 10137 23273 10149 23307
rect 10091 23267 10149 23273
rect 1464 23171 1522 23177
rect 1464 23137 1476 23171
rect 1510 23168 1522 23171
rect 1578 23168 1584 23180
rect 1510 23140 1584 23168
rect 1510 23137 1522 23140
rect 1464 23131 1522 23137
rect 1578 23128 1584 23140
rect 1636 23128 1642 23180
rect 10020 23171 10078 23177
rect 10020 23137 10032 23171
rect 10066 23168 10078 23171
rect 10134 23168 10140 23180
rect 10066 23140 10140 23168
rect 10066 23137 10078 23140
rect 10020 23131 10078 23137
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 1535 22967 1593 22973
rect 1535 22933 1547 22967
rect 1581 22964 1593 22967
rect 3786 22964 3792 22976
rect 1581 22936 3792 22964
rect 1581 22933 1593 22936
rect 1535 22927 1593 22933
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 9033 22763 9091 22769
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 9398 22760 9404 22772
rect 9079 22732 9404 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10137 22763 10195 22769
rect 10137 22729 10149 22763
rect 10183 22760 10195 22763
rect 11974 22760 11980 22772
rect 10183 22732 11980 22760
rect 10183 22729 10195 22732
rect 10137 22723 10195 22729
rect 11974 22720 11980 22732
rect 12032 22720 12038 22772
rect 24762 22760 24768 22772
rect 24723 22732 24768 22760
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 8849 22559 8907 22565
rect 8849 22525 8861 22559
rect 8895 22556 8907 22559
rect 9953 22559 10011 22565
rect 9953 22556 9965 22559
rect 8895 22528 9536 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 9508 22432 9536 22528
rect 9784 22528 9965 22556
rect 9784 22432 9812 22528
rect 9953 22525 9965 22528
rect 9999 22525 10011 22559
rect 9953 22519 10011 22525
rect 23658 22516 23664 22568
rect 23716 22556 23722 22568
rect 24581 22559 24639 22565
rect 24581 22556 24593 22559
rect 23716 22528 24593 22556
rect 23716 22516 23722 22528
rect 24581 22525 24593 22528
rect 24627 22556 24639 22559
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24627 22528 25145 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 25133 22519 25191 22525
rect 9490 22420 9496 22432
rect 9451 22392 9496 22420
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10505 22423 10563 22429
rect 10505 22420 10517 22423
rect 10192 22392 10517 22420
rect 10192 22380 10198 22392
rect 10505 22389 10517 22392
rect 10551 22389 10563 22423
rect 10505 22383 10563 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 11379 22219 11437 22225
rect 11379 22216 11391 22219
rect 9548 22188 11391 22216
rect 9548 22176 9554 22188
rect 11379 22185 11391 22188
rect 11425 22185 11437 22219
rect 11379 22179 11437 22185
rect 8272 22083 8330 22089
rect 8272 22049 8284 22083
rect 8318 22080 8330 22083
rect 8754 22080 8760 22092
rect 8318 22052 8760 22080
rect 8318 22049 8330 22052
rect 8272 22043 8330 22049
rect 8754 22040 8760 22052
rect 8812 22040 8818 22092
rect 9858 22080 9864 22092
rect 9819 22052 9864 22080
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 11238 22080 11244 22092
rect 11199 22052 11244 22080
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 7834 21836 7840 21888
rect 7892 21876 7898 21888
rect 8343 21879 8401 21885
rect 8343 21876 8355 21879
rect 7892 21848 8355 21876
rect 7892 21836 7898 21848
rect 8343 21845 8355 21848
rect 8389 21845 8401 21879
rect 9950 21876 9956 21888
rect 9911 21848 9956 21876
rect 8343 21839 8401 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 9355 21675 9413 21681
rect 9355 21641 9367 21675
rect 9401 21672 9413 21675
rect 9766 21672 9772 21684
rect 9401 21644 9772 21672
rect 9401 21641 9413 21644
rect 9355 21635 9413 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 8754 21536 8760 21548
rect 8715 21508 8760 21536
rect 8754 21496 8760 21508
rect 8812 21496 8818 21548
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21536 10563 21539
rect 10686 21536 10692 21548
rect 10551 21508 10692 21536
rect 10551 21505 10563 21508
rect 10505 21499 10563 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 10870 21536 10876 21548
rect 10831 21508 10876 21536
rect 10870 21496 10876 21508
rect 10928 21496 10934 21548
rect 7561 21471 7619 21477
rect 7561 21437 7573 21471
rect 7607 21468 7619 21471
rect 8294 21468 8300 21480
rect 7607 21440 8300 21468
rect 7607 21437 7619 21440
rect 7561 21431 7619 21437
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 9252 21471 9310 21477
rect 9252 21468 9264 21471
rect 9048 21440 9264 21468
rect 8113 21335 8171 21341
rect 8113 21301 8125 21335
rect 8159 21332 8171 21335
rect 8202 21332 8208 21344
rect 8159 21304 8208 21332
rect 8159 21301 8171 21304
rect 8113 21295 8171 21301
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 8846 21292 8852 21344
rect 8904 21332 8910 21344
rect 9048 21341 9076 21440
rect 9252 21437 9264 21440
rect 9298 21437 9310 21471
rect 9252 21431 9310 21437
rect 9674 21360 9680 21412
rect 9732 21400 9738 21412
rect 10229 21403 10287 21409
rect 10229 21400 10241 21403
rect 9732 21372 10241 21400
rect 9732 21360 9738 21372
rect 10229 21369 10241 21372
rect 10275 21400 10287 21403
rect 10597 21403 10655 21409
rect 10597 21400 10609 21403
rect 10275 21372 10609 21400
rect 10275 21369 10287 21372
rect 10229 21363 10287 21369
rect 10597 21369 10609 21372
rect 10643 21400 10655 21403
rect 11698 21400 11704 21412
rect 10643 21372 11704 21400
rect 10643 21369 10655 21372
rect 10597 21363 10655 21369
rect 11698 21360 11704 21372
rect 11756 21360 11762 21412
rect 9033 21335 9091 21341
rect 9033 21332 9045 21335
rect 8904 21304 9045 21332
rect 8904 21292 8910 21304
rect 9033 21301 9045 21304
rect 9079 21301 9091 21335
rect 9766 21332 9772 21344
rect 9727 21304 9772 21332
rect 9033 21295 9091 21301
rect 9766 21292 9772 21304
rect 9824 21292 9830 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 11238 21332 11244 21344
rect 10744 21304 11244 21332
rect 10744 21292 10750 21304
rect 11238 21292 11244 21304
rect 11296 21332 11302 21344
rect 11425 21335 11483 21341
rect 11425 21332 11437 21335
rect 11296 21304 11437 21332
rect 11296 21292 11302 21304
rect 11425 21301 11437 21304
rect 11471 21301 11483 21335
rect 11425 21295 11483 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 10042 21128 10048 21140
rect 9955 21100 10048 21128
rect 10042 21088 10048 21100
rect 10100 21128 10106 21140
rect 10100 21100 10916 21128
rect 10100 21088 10106 21100
rect 10888 21072 10916 21100
rect 7653 21063 7711 21069
rect 7653 21029 7665 21063
rect 7699 21060 7711 21063
rect 7834 21060 7840 21072
rect 7699 21032 7840 21060
rect 7699 21029 7711 21032
rect 7653 21023 7711 21029
rect 7834 21020 7840 21032
rect 7892 21020 7898 21072
rect 7926 21020 7932 21072
rect 7984 21060 7990 21072
rect 10318 21060 10324 21072
rect 7984 21032 8029 21060
rect 10279 21032 10324 21060
rect 7984 21020 7990 21032
rect 10318 21020 10324 21032
rect 10376 21020 10382 21072
rect 10870 21060 10876 21072
rect 10831 21032 10876 21060
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1946 20992 1952 21004
rect 1443 20964 1952 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1946 20952 1952 20964
rect 2004 20952 2010 21004
rect 6365 20995 6423 21001
rect 6365 20961 6377 20995
rect 6411 20992 6423 20995
rect 6638 20992 6644 21004
rect 6411 20964 6644 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 11790 20992 11796 21004
rect 11751 20964 11796 20992
rect 11790 20952 11796 20964
rect 11848 20952 11854 21004
rect 22830 21001 22836 21004
rect 22808 20995 22836 21001
rect 22808 20992 22820 20995
rect 22743 20964 22820 20992
rect 22808 20961 22820 20964
rect 22888 20992 22894 21004
rect 24670 20992 24676 21004
rect 22888 20964 24676 20992
rect 22808 20955 22836 20961
rect 22830 20952 22836 20955
rect 22888 20952 22894 20964
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 8110 20924 8116 20936
rect 8071 20896 8116 20924
rect 8110 20884 8116 20896
rect 8168 20884 8174 20936
rect 10226 20924 10232 20936
rect 10187 20896 10232 20924
rect 10226 20884 10232 20896
rect 10284 20884 10290 20936
rect 10318 20884 10324 20936
rect 10376 20924 10382 20936
rect 11054 20924 11060 20936
rect 10376 20896 11060 20924
rect 10376 20884 10382 20896
rect 11054 20884 11060 20896
rect 11112 20924 11118 20936
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 11112 20896 11713 20924
rect 11112 20884 11118 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 6549 20791 6607 20797
rect 6549 20757 6561 20791
rect 6595 20788 6607 20791
rect 6822 20788 6828 20800
rect 6595 20760 6828 20788
rect 6595 20757 6607 20760
rect 6549 20751 6607 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 8754 20788 8760 20800
rect 8715 20760 8760 20788
rect 8754 20748 8760 20760
rect 8812 20748 8818 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 22879 20791 22937 20797
rect 22879 20788 22891 20791
rect 18380 20760 22891 20788
rect 18380 20748 18386 20760
rect 22879 20757 22891 20760
rect 22925 20757 22937 20791
rect 22879 20751 22937 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 9861 20587 9919 20593
rect 9861 20553 9873 20587
rect 9907 20584 9919 20587
rect 9950 20584 9956 20596
rect 9907 20556 9956 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 11054 20584 11060 20596
rect 11015 20556 11060 20584
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11698 20584 11704 20596
rect 11659 20556 11704 20584
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 14001 20587 14059 20593
rect 14001 20584 14013 20587
rect 13786 20556 14013 20584
rect 9493 20519 9551 20525
rect 9493 20485 9505 20519
rect 9539 20516 9551 20519
rect 9539 20488 10272 20516
rect 9539 20485 9551 20488
rect 9493 20479 9551 20485
rect 10244 20460 10272 20488
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20448 7067 20451
rect 8113 20451 8171 20457
rect 8113 20448 8125 20451
rect 7055 20420 8125 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 8113 20417 8125 20420
rect 8159 20448 8171 20451
rect 8754 20448 8760 20460
rect 8159 20420 8760 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 10042 20448 10048 20460
rect 10003 20420 10048 20448
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10226 20408 10232 20460
rect 10284 20448 10290 20460
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 10284 20420 12449 20448
rect 10284 20408 10290 20420
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 12437 20411 12495 20417
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20380 4767 20383
rect 5788 20383 5846 20389
rect 4755 20352 5304 20380
rect 4755 20349 4767 20352
rect 4709 20343 4767 20349
rect 5276 20256 5304 20352
rect 5788 20349 5800 20383
rect 5834 20380 5846 20383
rect 13516 20383 13574 20389
rect 5834 20352 6316 20380
rect 5834 20349 5846 20352
rect 5788 20343 5846 20349
rect 6288 20256 6316 20352
rect 13516 20349 13528 20383
rect 13562 20380 13574 20383
rect 13786 20380 13814 20556
rect 14001 20553 14013 20556
rect 14047 20584 14059 20587
rect 14274 20584 14280 20596
rect 14047 20556 14280 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14274 20544 14280 20556
rect 14332 20584 14338 20596
rect 17494 20584 17500 20596
rect 14332 20556 17500 20584
rect 14332 20544 14338 20556
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 22830 20584 22836 20596
rect 22791 20556 22836 20584
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 13562 20352 13814 20380
rect 13562 20349 13574 20352
rect 13516 20343 13574 20349
rect 8202 20312 8208 20324
rect 8163 20284 8208 20312
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 8754 20312 8760 20324
rect 8715 20284 8760 20312
rect 8754 20272 8760 20284
rect 8812 20272 8818 20324
rect 10137 20315 10195 20321
rect 10137 20281 10149 20315
rect 10183 20281 10195 20315
rect 10686 20312 10692 20324
rect 10647 20284 10692 20312
rect 10137 20275 10195 20281
rect 1673 20247 1731 20253
rect 1673 20213 1685 20247
rect 1719 20244 1731 20247
rect 1946 20244 1952 20256
rect 1719 20216 1952 20244
rect 1719 20213 1731 20216
rect 1673 20207 1731 20213
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 4893 20247 4951 20253
rect 4893 20244 4905 20247
rect 3752 20216 4905 20244
rect 3752 20204 3758 20216
rect 4893 20213 4905 20216
rect 4939 20213 4951 20247
rect 5258 20244 5264 20256
rect 5219 20216 5264 20244
rect 4893 20207 4951 20213
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5859 20247 5917 20253
rect 5859 20213 5871 20247
rect 5905 20244 5917 20247
rect 5994 20244 6000 20256
rect 5905 20216 6000 20244
rect 5905 20213 5917 20216
rect 5859 20207 5917 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6270 20244 6276 20256
rect 6231 20216 6276 20244
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 6638 20244 6644 20256
rect 6599 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 7745 20247 7803 20253
rect 7745 20244 7757 20247
rect 7248 20216 7757 20244
rect 7248 20204 7254 20216
rect 7745 20213 7757 20216
rect 7791 20244 7803 20247
rect 7926 20244 7932 20256
rect 7791 20216 7932 20244
rect 7791 20213 7803 20216
rect 7745 20207 7803 20213
rect 7926 20204 7932 20216
rect 7984 20204 7990 20256
rect 8220 20244 8248 20272
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 8220 20216 9045 20244
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 9033 20207 9091 20213
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10152 20244 10180 20275
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 10008 20216 10180 20244
rect 10008 20204 10014 20216
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13587 20247 13645 20253
rect 13587 20244 13599 20247
rect 13136 20216 13599 20244
rect 13136 20204 13142 20216
rect 13587 20213 13599 20216
rect 13633 20213 13645 20247
rect 13587 20207 13645 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 11756 20012 13216 20040
rect 11756 20000 11762 20012
rect 7190 19972 7196 19984
rect 7151 19944 7196 19972
rect 7190 19932 7196 19944
rect 7248 19932 7254 19984
rect 8110 19972 8116 19984
rect 8071 19944 8116 19972
rect 8110 19932 8116 19944
rect 8168 19932 8174 19984
rect 8202 19932 8208 19984
rect 8260 19972 8266 19984
rect 8754 19972 8760 19984
rect 8260 19944 8305 19972
rect 8715 19944 8760 19972
rect 8260 19932 8266 19944
rect 8754 19932 8760 19944
rect 8812 19932 8818 19984
rect 9766 19932 9772 19984
rect 9824 19972 9830 19984
rect 10045 19975 10103 19981
rect 10045 19972 10057 19975
rect 9824 19944 10057 19972
rect 9824 19932 9830 19944
rect 10045 19941 10057 19944
rect 10091 19941 10103 19975
rect 10045 19935 10103 19941
rect 10597 19975 10655 19981
rect 10597 19941 10609 19975
rect 10643 19972 10655 19975
rect 10686 19972 10692 19984
rect 10643 19944 10692 19972
rect 10643 19941 10655 19944
rect 10597 19935 10655 19941
rect 10686 19932 10692 19944
rect 10744 19932 10750 19984
rect 11606 19972 11612 19984
rect 11567 19944 11612 19972
rect 11606 19932 11612 19944
rect 11664 19932 11670 19984
rect 13078 19972 13084 19984
rect 13039 19944 13084 19972
rect 13078 19932 13084 19944
rect 13136 19932 13142 19984
rect 13188 19981 13216 20012
rect 13173 19975 13231 19981
rect 13173 19941 13185 19975
rect 13219 19972 13231 19975
rect 13262 19972 13268 19984
rect 13219 19944 13268 19972
rect 13219 19941 13231 19944
rect 13173 19935 13231 19941
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 4982 19904 4988 19916
rect 4943 19876 4988 19904
rect 4982 19864 4988 19876
rect 5040 19864 5046 19916
rect 6546 19904 6552 19916
rect 6507 19876 6552 19904
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 3970 19796 3976 19848
rect 4028 19836 4034 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 4028 19808 4353 19836
rect 4028 19796 4034 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 9950 19836 9956 19848
rect 9911 19808 9956 19836
rect 4341 19799 4399 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 11422 19728 11428 19780
rect 11480 19768 11486 19780
rect 11532 19768 11560 19799
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11756 19808 11805 19836
rect 11756 19796 11762 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 11793 19799 11851 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 11480 19740 11560 19768
rect 11480 19728 11486 19740
rect 7650 19700 7656 19712
rect 7611 19672 7656 19700
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 13722 19660 13728 19712
rect 13780 19700 13786 19712
rect 14001 19703 14059 19709
rect 14001 19700 14013 19703
rect 13780 19672 14013 19700
rect 13780 19660 13786 19672
rect 14001 19669 14013 19672
rect 14047 19669 14059 19703
rect 14001 19663 14059 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 4062 19496 4068 19508
rect 3927 19468 4068 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 4062 19456 4068 19468
rect 4120 19496 4126 19508
rect 4982 19496 4988 19508
rect 4120 19468 4988 19496
rect 4120 19456 4126 19468
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 6546 19496 6552 19508
rect 6507 19468 6552 19496
rect 6546 19456 6552 19468
rect 6604 19496 6610 19508
rect 7377 19499 7435 19505
rect 7377 19496 7389 19499
rect 6604 19468 7389 19496
rect 6604 19456 6610 19468
rect 7377 19465 7389 19468
rect 7423 19496 7435 19499
rect 7742 19496 7748 19508
rect 7423 19468 7748 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 10134 19496 10140 19508
rect 10095 19468 10140 19496
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 13262 19496 13268 19508
rect 13223 19468 13268 19496
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 5721 19431 5779 19437
rect 5721 19397 5733 19431
rect 5767 19428 5779 19431
rect 7190 19428 7196 19440
rect 5767 19400 7196 19428
rect 5767 19397 5779 19400
rect 5721 19391 5779 19397
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 9490 19388 9496 19440
rect 9548 19428 9554 19440
rect 12713 19431 12771 19437
rect 12713 19428 12725 19431
rect 9548 19400 12725 19428
rect 9548 19388 9554 19400
rect 12713 19397 12725 19400
rect 12759 19428 12771 19431
rect 12897 19431 12955 19437
rect 12897 19428 12909 19431
rect 12759 19400 12909 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 12897 19397 12909 19400
rect 12943 19397 12955 19431
rect 12897 19391 12955 19397
rect 4338 19360 4344 19372
rect 4299 19332 4344 19360
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 8110 19360 8116 19372
rect 8071 19332 8116 19360
rect 8110 19320 8116 19332
rect 8168 19320 8174 19372
rect 9033 19363 9091 19369
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9950 19360 9956 19372
rect 9079 19332 9956 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9950 19320 9956 19332
rect 10008 19360 10014 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10008 19332 10977 19360
rect 10008 19320 10014 19332
rect 10965 19329 10977 19332
rect 11011 19360 11023 19363
rect 13354 19360 13360 19372
rect 11011 19332 13360 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 1118 19252 1124 19304
rect 1176 19292 1182 19304
rect 1397 19295 1455 19301
rect 1397 19292 1409 19295
rect 1176 19264 1409 19292
rect 1176 19252 1182 19264
rect 1397 19261 1409 19264
rect 1443 19292 1455 19295
rect 1949 19295 2007 19301
rect 1949 19292 1961 19295
rect 1443 19264 1961 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1949 19261 1961 19264
rect 1995 19261 2007 19295
rect 1949 19255 2007 19261
rect 2568 19295 2626 19301
rect 2568 19261 2580 19295
rect 2614 19292 2626 19295
rect 2614 19264 3096 19292
rect 2614 19261 2626 19264
rect 2568 19255 2626 19261
rect 3068 19168 3096 19264
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5537 19295 5595 19301
rect 5537 19292 5549 19295
rect 5316 19264 5549 19292
rect 5316 19252 5322 19264
rect 5537 19261 5549 19264
rect 5583 19292 5595 19295
rect 5583 19264 6132 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 4065 19227 4123 19233
rect 4065 19193 4077 19227
rect 4111 19193 4123 19227
rect 4065 19187 4123 19193
rect 2038 19116 2044 19168
rect 2096 19156 2102 19168
rect 2639 19159 2697 19165
rect 2639 19156 2651 19159
rect 2096 19128 2651 19156
rect 2096 19116 2102 19128
rect 2639 19125 2651 19128
rect 2685 19125 2697 19159
rect 3050 19156 3056 19168
rect 3011 19128 3056 19156
rect 2639 19119 2697 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3418 19156 3424 19168
rect 3379 19128 3424 19156
rect 3418 19116 3424 19128
rect 3476 19156 3482 19168
rect 4080 19156 4108 19187
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 4212 19196 4257 19224
rect 4212 19184 4218 19196
rect 6104 19165 6132 19264
rect 8570 19252 8576 19304
rect 8628 19292 8634 19304
rect 9125 19295 9183 19301
rect 9125 19292 9137 19295
rect 8628 19264 9137 19292
rect 8628 19252 8634 19264
rect 9125 19261 9137 19264
rect 9171 19292 9183 19295
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 9171 19264 9597 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 12504 19295 12562 19301
rect 12504 19261 12516 19295
rect 12550 19292 12562 19295
rect 12713 19295 12771 19301
rect 12713 19292 12725 19295
rect 12550 19264 12725 19292
rect 12550 19261 12562 19264
rect 12504 19255 12562 19261
rect 12713 19261 12725 19264
rect 12759 19261 12771 19295
rect 12713 19255 12771 19261
rect 7650 19224 7656 19236
rect 7611 19196 7656 19224
rect 7650 19184 7656 19196
rect 7708 19184 7714 19236
rect 7742 19184 7748 19236
rect 7800 19224 7806 19236
rect 7800 19196 7845 19224
rect 7800 19184 7806 19196
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10321 19227 10379 19233
rect 10321 19224 10333 19227
rect 10008 19196 10333 19224
rect 10008 19184 10014 19196
rect 10321 19193 10333 19196
rect 10367 19193 10379 19227
rect 10321 19187 10379 19193
rect 10413 19227 10471 19233
rect 10413 19193 10425 19227
rect 10459 19193 10471 19227
rect 11606 19224 11612 19236
rect 10413 19187 10471 19193
rect 11302 19196 11612 19224
rect 3476 19128 4108 19156
rect 6089 19159 6147 19165
rect 3476 19116 3482 19128
rect 6089 19125 6101 19159
rect 6135 19156 6147 19159
rect 6730 19156 6736 19168
rect 6135 19128 6736 19156
rect 6135 19125 6147 19128
rect 6089 19119 6147 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 8202 19156 8208 19168
rect 7892 19128 8208 19156
rect 7892 19116 7898 19128
rect 8202 19116 8208 19128
rect 8260 19156 8266 19168
rect 8573 19159 8631 19165
rect 8573 19156 8585 19159
rect 8260 19128 8585 19156
rect 8260 19116 8266 19128
rect 8573 19125 8585 19128
rect 8619 19125 8631 19159
rect 8573 19119 8631 19125
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 9309 19159 9367 19165
rect 9309 19156 9321 19159
rect 9180 19128 9321 19156
rect 9180 19116 9186 19128
rect 9309 19125 9321 19128
rect 9355 19125 9367 19159
rect 9309 19119 9367 19125
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10428 19156 10456 19187
rect 10192 19128 10456 19156
rect 10192 19116 10198 19128
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11302 19156 11330 19196
rect 11606 19184 11612 19196
rect 11664 19224 11670 19236
rect 11793 19227 11851 19233
rect 11793 19224 11805 19227
rect 11664 19196 11805 19224
rect 11664 19184 11670 19196
rect 11793 19193 11805 19196
rect 11839 19193 11851 19227
rect 11793 19187 11851 19193
rect 13725 19227 13783 19233
rect 13725 19193 13737 19227
rect 13771 19193 13783 19227
rect 13725 19187 13783 19193
rect 13817 19227 13875 19233
rect 13817 19193 13829 19227
rect 13863 19224 13875 19227
rect 13998 19224 14004 19236
rect 13863 19196 14004 19224
rect 13863 19193 13875 19196
rect 13817 19187 13875 19193
rect 11422 19156 11428 19168
rect 10928 19128 11330 19156
rect 11383 19128 11428 19156
rect 10928 19116 10934 19128
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 12575 19159 12633 19165
rect 12575 19156 12587 19159
rect 12308 19128 12587 19156
rect 12308 19116 12314 19128
rect 12575 19125 12587 19128
rect 12621 19125 12633 19159
rect 12575 19119 12633 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13740 19156 13768 19187
rect 13998 19184 14004 19196
rect 14056 19184 14062 19236
rect 14366 19224 14372 19236
rect 14327 19196 14372 19224
rect 14366 19184 14372 19196
rect 14424 19184 14430 19236
rect 14645 19159 14703 19165
rect 14645 19156 14657 19159
rect 13412 19128 14657 19156
rect 13412 19116 13418 19128
rect 14645 19125 14657 19128
rect 14691 19125 14703 19159
rect 14645 19119 14703 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1535 18955 1593 18961
rect 1535 18921 1547 18955
rect 1581 18952 1593 18955
rect 3418 18952 3424 18964
rect 1581 18924 3424 18952
rect 1581 18921 1593 18924
rect 1535 18915 1593 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 6914 18912 6920 18964
rect 6972 18952 6978 18964
rect 7653 18955 7711 18961
rect 6972 18924 7281 18952
rect 6972 18912 6978 18924
rect 5074 18884 5080 18896
rect 5035 18856 5080 18884
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 7098 18893 7104 18896
rect 7095 18884 7104 18893
rect 7059 18856 7104 18884
rect 7095 18847 7104 18856
rect 7098 18844 7104 18847
rect 7156 18844 7162 18896
rect 7253 18884 7281 18924
rect 7653 18921 7665 18955
rect 7699 18952 7711 18955
rect 7742 18952 7748 18964
rect 7699 18924 7748 18952
rect 7699 18921 7711 18924
rect 7653 18915 7711 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8110 18912 8116 18964
rect 8168 18952 8174 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8168 18924 8309 18952
rect 8168 18912 8174 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 13078 18952 13084 18964
rect 13039 18924 13084 18952
rect 8297 18915 8355 18921
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 13998 18952 14004 18964
rect 13780 18924 14004 18952
rect 13780 18912 13786 18924
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 9490 18884 9496 18896
rect 7253 18856 9496 18884
rect 9490 18844 9496 18856
rect 9548 18884 9554 18896
rect 10870 18884 10876 18896
rect 9548 18856 9720 18884
rect 10831 18856 10876 18884
rect 9548 18844 9554 18856
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 8478 18816 8484 18828
rect 8439 18788 8484 18816
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 9692 18825 9720 18856
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 13814 18844 13820 18896
rect 13872 18884 13878 18896
rect 14366 18884 14372 18896
rect 13872 18856 13917 18884
rect 14327 18856 14372 18884
rect 13872 18844 13878 18856
rect 14366 18844 14372 18856
rect 14424 18884 14430 18896
rect 16482 18884 16488 18896
rect 14424 18856 16252 18884
rect 16443 18856 16488 18884
rect 14424 18844 14430 18856
rect 9692 18819 9770 18825
rect 9692 18788 9724 18819
rect 9712 18785 9724 18788
rect 9758 18785 9770 18819
rect 12618 18816 12624 18828
rect 12579 18788 12624 18816
rect 9712 18779 9770 18785
rect 12618 18776 12624 18788
rect 12676 18776 12682 18828
rect 15356 18819 15414 18825
rect 15356 18785 15368 18819
rect 15402 18816 15414 18819
rect 15470 18816 15476 18828
rect 15402 18788 15476 18816
rect 15402 18785 15414 18788
rect 15356 18779 15414 18785
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 2958 18748 2964 18760
rect 2919 18720 2964 18748
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 5350 18748 5356 18760
rect 5031 18720 5356 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18748 6791 18751
rect 6914 18748 6920 18760
rect 6779 18720 6920 18748
rect 6779 18717 6791 18720
rect 6733 18711 6791 18717
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 9815 18751 9873 18757
rect 9815 18717 9827 18751
rect 9861 18748 9873 18751
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 9861 18720 10793 18748
rect 9861 18717 9873 18720
rect 9815 18711 9873 18717
rect 10781 18717 10793 18720
rect 10827 18748 10839 18751
rect 11146 18748 11152 18760
rect 10827 18720 11152 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11296 18720 11341 18748
rect 11296 18708 11302 18720
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13504 18720 13737 18748
rect 13504 18708 13510 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 13725 18711 13783 18717
rect 14200 18720 15945 18748
rect 5534 18680 5540 18692
rect 5495 18652 5540 18680
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 9306 18640 9312 18692
rect 9364 18680 9370 18692
rect 9950 18680 9956 18692
rect 9364 18652 9956 18680
rect 9364 18640 9370 18652
rect 9950 18640 9956 18652
rect 10008 18680 10014 18692
rect 10505 18683 10563 18689
rect 10505 18680 10517 18683
rect 10008 18652 10517 18680
rect 10008 18640 10014 18652
rect 10505 18649 10517 18652
rect 10551 18649 10563 18683
rect 10505 18643 10563 18649
rect 12759 18683 12817 18689
rect 12759 18649 12771 18683
rect 12805 18680 12817 18683
rect 14200 18680 14228 18720
rect 15933 18717 15945 18720
rect 15979 18748 15991 18751
rect 16022 18748 16028 18760
rect 15979 18720 16028 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16224 18748 16252 18856
rect 16482 18844 16488 18856
rect 16540 18844 16546 18896
rect 16574 18844 16580 18896
rect 16632 18884 16638 18896
rect 16632 18856 16677 18884
rect 16632 18844 16638 18856
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 16224 18720 16773 18748
rect 16761 18717 16773 18720
rect 16807 18748 16819 18751
rect 17678 18748 17684 18760
rect 16807 18720 17684 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 12805 18652 14228 18680
rect 12805 18649 12817 18652
rect 12759 18643 12817 18649
rect 7926 18612 7932 18624
rect 7887 18584 7932 18612
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 8665 18615 8723 18621
rect 8665 18612 8677 18615
rect 8260 18584 8677 18612
rect 8260 18572 8266 18584
rect 8665 18581 8677 18584
rect 8711 18581 8723 18615
rect 8665 18575 8723 18581
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 9766 18612 9772 18624
rect 8812 18584 9772 18612
rect 8812 18572 8818 18584
rect 9766 18572 9772 18584
rect 9824 18612 9830 18624
rect 10137 18615 10195 18621
rect 10137 18612 10149 18615
rect 9824 18584 10149 18612
rect 9824 18572 9830 18584
rect 10137 18581 10149 18584
rect 10183 18581 10195 18615
rect 13446 18612 13452 18624
rect 13407 18584 13452 18612
rect 10137 18575 10195 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14642 18612 14648 18624
rect 13780 18584 14648 18612
rect 13780 18572 13786 18584
rect 14642 18572 14648 18584
rect 14700 18612 14706 18624
rect 15427 18615 15485 18621
rect 15427 18612 15439 18615
rect 14700 18584 15439 18612
rect 14700 18572 14706 18584
rect 15427 18581 15439 18584
rect 15473 18581 15485 18615
rect 15427 18575 15485 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 2317 18411 2375 18417
rect 2317 18408 2329 18411
rect 1452 18380 2329 18408
rect 1452 18368 1458 18380
rect 2317 18377 2329 18380
rect 2363 18377 2375 18411
rect 4798 18408 4804 18420
rect 2317 18371 2375 18377
rect 4126 18380 4804 18408
rect 2041 18343 2099 18349
rect 2041 18309 2053 18343
rect 2087 18340 2099 18343
rect 4126 18340 4154 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5074 18408 5080 18420
rect 4939 18380 5080 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 2087 18312 4154 18340
rect 2087 18309 2099 18312
rect 2041 18303 2099 18309
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2056 18204 2084 18303
rect 2958 18232 2964 18284
rect 3016 18272 3022 18284
rect 3510 18272 3516 18284
rect 3016 18244 3516 18272
rect 3016 18232 3022 18244
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 4338 18272 4344 18284
rect 4203 18244 4344 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 1443 18176 2084 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 3329 18139 3387 18145
rect 3329 18105 3341 18139
rect 3375 18136 3387 18139
rect 3605 18139 3663 18145
rect 3605 18136 3617 18139
rect 3375 18108 3617 18136
rect 3375 18105 3387 18108
rect 3329 18099 3387 18105
rect 3605 18105 3617 18108
rect 3651 18136 3663 18139
rect 3970 18136 3976 18148
rect 3651 18108 3976 18136
rect 3651 18105 3663 18108
rect 3605 18099 3663 18105
rect 3970 18096 3976 18108
rect 4028 18136 4034 18148
rect 4908 18136 4936 18371
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6963 18411 7021 18417
rect 6963 18377 6975 18411
rect 7009 18408 7021 18411
rect 7650 18408 7656 18420
rect 7009 18380 7656 18408
rect 7009 18377 7021 18380
rect 6963 18371 7021 18377
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 8757 18411 8815 18417
rect 8757 18377 8769 18411
rect 8803 18408 8815 18411
rect 9674 18408 9680 18420
rect 8803 18380 9680 18408
rect 8803 18377 8815 18380
rect 8757 18371 8815 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 11701 18411 11759 18417
rect 11701 18377 11713 18411
rect 11747 18408 11759 18411
rect 11790 18408 11796 18420
rect 11747 18380 11796 18408
rect 11747 18377 11759 18380
rect 11701 18371 11759 18377
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12618 18368 12624 18420
rect 12676 18408 12682 18420
rect 14826 18408 14832 18420
rect 12676 18380 14832 18408
rect 12676 18368 12682 18380
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 15470 18408 15476 18420
rect 15383 18380 15476 18408
rect 15470 18368 15476 18380
rect 15528 18408 15534 18420
rect 19426 18408 19432 18420
rect 15528 18380 19432 18408
rect 15528 18368 15534 18380
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 25130 18408 25136 18420
rect 25091 18380 25136 18408
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 6012 18340 6040 18368
rect 5092 18312 6040 18340
rect 5092 18281 5120 18312
rect 8478 18300 8484 18352
rect 8536 18340 8542 18352
rect 8846 18340 8852 18352
rect 8536 18312 8852 18340
rect 8536 18300 8542 18312
rect 8846 18300 8852 18312
rect 8904 18340 8910 18352
rect 9033 18343 9091 18349
rect 9033 18340 9045 18343
rect 8904 18312 9045 18340
rect 8904 18300 8910 18312
rect 9033 18309 9045 18312
rect 9079 18309 9091 18343
rect 9033 18303 9091 18309
rect 9134 18312 11259 18340
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5534 18272 5540 18284
rect 5495 18244 5540 18272
rect 5077 18235 5135 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 6270 18232 6276 18284
rect 6328 18272 6334 18284
rect 9134 18272 9162 18312
rect 6328 18244 9162 18272
rect 6328 18232 6334 18244
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9272 18244 9689 18272
rect 9272 18232 9278 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 6892 18207 6950 18213
rect 6892 18204 6904 18207
rect 5776 18176 6904 18204
rect 5776 18164 5782 18176
rect 6892 18173 6904 18176
rect 6938 18204 6950 18207
rect 7837 18207 7895 18213
rect 6938 18176 7328 18204
rect 6938 18173 6950 18176
rect 6892 18167 6950 18173
rect 4028 18108 4936 18136
rect 5169 18139 5227 18145
rect 4028 18096 4034 18108
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 5258 18136 5264 18148
rect 5215 18108 5264 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 106 18028 112 18080
rect 164 18068 170 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 164 18040 1593 18068
rect 164 18028 170 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4212 18040 4537 18068
rect 4212 18028 4218 18040
rect 4525 18037 4537 18040
rect 4571 18068 4583 18071
rect 5184 18068 5212 18099
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 7300 18080 7328 18176
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7926 18204 7932 18216
rect 7883 18176 7932 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9490 18204 9496 18216
rect 9451 18176 9496 18204
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 11231 18213 11259 18312
rect 12268 18272 12296 18368
rect 13449 18343 13507 18349
rect 13449 18309 13461 18343
rect 13495 18340 13507 18343
rect 13630 18340 13636 18352
rect 13495 18312 13636 18340
rect 13495 18309 13507 18312
rect 13449 18303 13507 18309
rect 13630 18300 13636 18312
rect 13688 18340 13694 18352
rect 13688 18312 16344 18340
rect 13688 18300 13694 18312
rect 16316 18284 16344 18312
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12268 18244 12909 18272
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 12897 18235 12955 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16298 18272 16304 18284
rect 16211 18244 16304 18272
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 11216 18207 11274 18213
rect 11216 18173 11228 18207
rect 11262 18204 11274 18207
rect 11790 18204 11796 18216
rect 11262 18176 11796 18204
rect 11262 18173 11274 18176
rect 11216 18167 11274 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 24648 18207 24706 18213
rect 24648 18173 24660 18207
rect 24694 18204 24706 18207
rect 25130 18204 25136 18216
rect 24694 18176 25136 18204
rect 24694 18173 24706 18176
rect 24648 18167 24706 18173
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 8158 18139 8216 18145
rect 8158 18105 8170 18139
rect 8204 18105 8216 18139
rect 8158 18099 8216 18105
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18105 9827 18139
rect 9769 18099 9827 18105
rect 10321 18139 10379 18145
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 10686 18136 10692 18148
rect 10367 18108 10692 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 4571 18040 5212 18068
rect 6641 18071 6699 18077
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 6641 18037 6653 18071
rect 6687 18068 6699 18071
rect 7098 18068 7104 18080
rect 6687 18040 7104 18068
rect 6687 18037 6699 18040
rect 6641 18031 6699 18037
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7742 18068 7748 18080
rect 7703 18040 7748 18068
rect 7742 18028 7748 18040
rect 7800 18068 7806 18080
rect 8173 18068 8201 18099
rect 7800 18040 8201 18068
rect 9784 18068 9812 18099
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18136 13047 18139
rect 14277 18139 14335 18145
rect 13035 18108 13584 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 13556 18080 13584 18108
rect 14277 18105 14289 18139
rect 14323 18136 14335 18139
rect 14458 18136 14464 18148
rect 14323 18108 14464 18136
rect 14323 18105 14335 18108
rect 14277 18099 14335 18105
rect 14458 18096 14464 18108
rect 14516 18096 14522 18148
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 16117 18139 16175 18145
rect 14608 18108 14653 18136
rect 14608 18096 14614 18108
rect 16117 18105 16129 18139
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 9784 18040 10609 18068
rect 7800 18028 7806 18040
rect 10597 18037 10609 18040
rect 10643 18068 10655 18071
rect 10778 18068 10784 18080
rect 10643 18040 10784 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 10965 18071 11023 18077
rect 10965 18068 10977 18071
rect 10928 18040 10977 18068
rect 10928 18028 10934 18040
rect 10965 18037 10977 18040
rect 11011 18037 11023 18071
rect 10965 18031 11023 18037
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11287 18071 11345 18077
rect 11287 18068 11299 18071
rect 11112 18040 11299 18068
rect 11112 18028 11118 18040
rect 11287 18037 11299 18040
rect 11333 18037 11345 18071
rect 12618 18068 12624 18080
rect 12579 18040 12624 18068
rect 11287 18031 11345 18037
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 13814 18068 13820 18080
rect 13596 18040 13820 18068
rect 13596 18028 13602 18040
rect 13814 18028 13820 18040
rect 13872 18068 13878 18080
rect 13909 18071 13967 18077
rect 13909 18068 13921 18071
rect 13872 18040 13921 18068
rect 13872 18028 13878 18040
rect 13909 18037 13921 18040
rect 13955 18068 13967 18071
rect 14568 18068 14596 18096
rect 15746 18068 15752 18080
rect 13955 18040 14596 18068
rect 15707 18040 15752 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 16132 18068 16160 18099
rect 16574 18068 16580 18080
rect 15804 18040 16580 18068
rect 15804 18028 15810 18040
rect 16574 18028 16580 18040
rect 16632 18068 16638 18080
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16632 18040 16957 18068
rect 16632 18028 16638 18040
rect 16945 18037 16957 18040
rect 16991 18037 17003 18071
rect 16945 18031 17003 18037
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 24719 18071 24777 18077
rect 24719 18068 24731 18071
rect 18656 18040 24731 18068
rect 18656 18028 18662 18040
rect 24719 18037 24731 18040
rect 24765 18037 24777 18071
rect 24719 18031 24777 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2038 17864 2044 17876
rect 1999 17836 2044 17864
rect 2038 17824 2044 17836
rect 2096 17824 2102 17876
rect 3510 17864 3516 17876
rect 3471 17836 3516 17864
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4338 17864 4344 17876
rect 4299 17836 4344 17864
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 7834 17864 7840 17876
rect 7795 17836 7840 17864
rect 7834 17824 7840 17836
rect 7892 17824 7898 17876
rect 9214 17824 9220 17876
rect 9272 17864 9278 17876
rect 9401 17867 9459 17873
rect 9401 17864 9413 17867
rect 9272 17836 9413 17864
rect 9272 17824 9278 17836
rect 9401 17833 9413 17836
rect 9447 17833 9459 17867
rect 9401 17827 9459 17833
rect 10873 17867 10931 17873
rect 10873 17833 10885 17867
rect 10919 17864 10931 17867
rect 11054 17864 11060 17876
rect 10919 17836 11060 17864
rect 10919 17833 10931 17836
rect 10873 17827 10931 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 12897 17867 12955 17873
rect 11204 17836 11249 17864
rect 11204 17824 11210 17836
rect 12897 17833 12909 17867
rect 12943 17864 12955 17867
rect 13538 17864 13544 17876
rect 12943 17836 13544 17864
rect 12943 17833 12955 17836
rect 12897 17827 12955 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 16482 17864 16488 17876
rect 16443 17836 16488 17864
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 4356 17796 4384 17824
rect 4617 17799 4675 17805
rect 4617 17796 4629 17799
rect 4356 17768 4629 17796
rect 4617 17765 4629 17768
rect 4663 17765 4675 17799
rect 4617 17759 4675 17765
rect 4706 17756 4712 17808
rect 4764 17796 4770 17808
rect 4764 17768 4809 17796
rect 4764 17756 4770 17768
rect 7098 17756 7104 17808
rect 7156 17796 7162 17808
rect 7279 17799 7337 17805
rect 7279 17796 7291 17799
rect 7156 17768 7291 17796
rect 7156 17756 7162 17768
rect 7279 17765 7291 17768
rect 7325 17796 7337 17799
rect 7742 17796 7748 17808
rect 7325 17768 7748 17796
rect 7325 17765 7337 17768
rect 7279 17759 7337 17765
rect 7742 17756 7748 17768
rect 7800 17756 7806 17808
rect 9858 17796 9864 17808
rect 9819 17768 9864 17796
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 10778 17756 10784 17808
rect 10836 17796 10842 17808
rect 11517 17799 11575 17805
rect 11517 17796 11529 17799
rect 10836 17768 11529 17796
rect 10836 17756 10842 17768
rect 11517 17765 11529 17768
rect 11563 17796 11575 17799
rect 11790 17796 11796 17808
rect 11563 17768 11796 17796
rect 11563 17765 11575 17768
rect 11517 17759 11575 17765
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 13722 17796 13728 17808
rect 13683 17768 13728 17796
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 13817 17799 13875 17805
rect 13817 17765 13829 17799
rect 13863 17796 13875 17799
rect 13998 17796 14004 17808
rect 13863 17768 14004 17796
rect 13863 17765 13875 17768
rect 13817 17759 13875 17765
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 14458 17756 14464 17808
rect 14516 17796 14522 17808
rect 16853 17799 16911 17805
rect 16853 17796 16865 17799
rect 14516 17768 16865 17796
rect 14516 17756 14522 17768
rect 16853 17765 16865 17768
rect 16899 17765 16911 17799
rect 16853 17759 16911 17765
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1578 17728 1584 17740
rect 1443 17700 1584 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2498 17728 2504 17740
rect 2459 17700 2504 17728
rect 2498 17688 2504 17700
rect 2556 17688 2562 17740
rect 5350 17688 5356 17740
rect 5408 17728 5414 17740
rect 5626 17728 5632 17740
rect 5408 17700 5632 17728
rect 5408 17688 5414 17700
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 15562 17688 15568 17740
rect 15620 17728 15626 17740
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 15620 17700 15761 17728
rect 15620 17688 15626 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 2639 17663 2697 17669
rect 2639 17629 2651 17663
rect 2685 17660 2697 17663
rect 3418 17660 3424 17672
rect 2685 17632 3424 17660
rect 2685 17629 2697 17632
rect 2639 17623 2697 17629
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 4908 17592 4936 17623
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 6236 17632 6929 17660
rect 6236 17620 6242 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 8662 17620 8668 17672
rect 8720 17660 8726 17672
rect 9582 17660 9588 17672
rect 8720 17632 9588 17660
rect 8720 17620 8726 17632
rect 9582 17620 9588 17632
rect 9640 17660 9646 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9640 17632 9781 17660
rect 9640 17620 9646 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17660 10471 17663
rect 10686 17660 10692 17672
rect 10459 17632 10692 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 10686 17620 10692 17632
rect 10744 17660 10750 17672
rect 11238 17660 11244 17672
rect 10744 17632 11244 17660
rect 10744 17620 10750 17632
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 12250 17660 12256 17672
rect 11471 17632 12256 17660
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 14001 17663 14059 17669
rect 14001 17660 14013 17663
rect 13786 17632 14013 17660
rect 5166 17592 5172 17604
rect 3108 17564 5172 17592
rect 3108 17552 3114 17564
rect 5166 17552 5172 17564
rect 5224 17552 5230 17604
rect 11974 17592 11980 17604
rect 11935 17564 11980 17592
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 13786 17592 13814 17632
rect 14001 17629 14013 17632
rect 14047 17629 14059 17663
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 14001 17623 14059 17629
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 13688 17564 13814 17592
rect 13688 17552 13694 17564
rect 2314 17524 2320 17536
rect 2275 17496 2320 17524
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 2958 17524 2964 17536
rect 2919 17496 2964 17524
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 6825 17527 6883 17533
rect 6825 17493 6837 17527
rect 6871 17524 6883 17527
rect 6914 17524 6920 17536
rect 6871 17496 6920 17524
rect 6871 17493 6883 17496
rect 6825 17487 6883 17493
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 4617 17323 4675 17329
rect 4617 17320 4629 17323
rect 4126 17292 4629 17320
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17184 4031 17187
rect 4126 17184 4154 17292
rect 4617 17289 4629 17292
rect 4663 17320 4675 17323
rect 4706 17320 4712 17332
rect 4663 17292 4712 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 8754 17320 8760 17332
rect 8715 17292 8760 17320
rect 8754 17280 8760 17292
rect 8812 17280 8818 17332
rect 9582 17320 9588 17332
rect 9543 17292 9588 17320
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10229 17323 10287 17329
rect 10229 17320 10241 17323
rect 9916 17292 10241 17320
rect 9916 17280 9922 17292
rect 10229 17289 10241 17292
rect 10275 17320 10287 17323
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 10275 17292 10425 17320
rect 10275 17289 10287 17292
rect 10229 17283 10287 17289
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 10413 17283 10471 17289
rect 10520 17292 13001 17320
rect 5534 17252 5540 17264
rect 4908 17224 5540 17252
rect 4908 17193 4936 17224
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 7377 17255 7435 17261
rect 7377 17221 7389 17255
rect 7423 17252 7435 17255
rect 10520 17252 10548 17292
rect 7423 17224 10548 17252
rect 7423 17221 7435 17224
rect 7377 17215 7435 17221
rect 4019 17156 4154 17184
rect 4893 17187 4951 17193
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 4893 17153 4905 17187
rect 4939 17153 4951 17187
rect 5166 17184 5172 17196
rect 5127 17156 5172 17184
rect 4893 17147 4951 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2038 17116 2044 17128
rect 1443 17088 2044 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17116 3203 17119
rect 3329 17119 3387 17125
rect 3329 17116 3341 17119
rect 3191 17088 3341 17116
rect 3191 17085 3203 17088
rect 3145 17079 3203 17085
rect 3329 17085 3341 17088
rect 3375 17116 3387 17119
rect 6892 17119 6950 17125
rect 3375 17088 4154 17116
rect 3375 17085 3387 17088
rect 3329 17079 3387 17085
rect 4126 17048 4154 17088
rect 6892 17085 6904 17119
rect 6938 17116 6950 17119
rect 7392 17116 7420 17215
rect 8772 17196 8800 17224
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 8110 17184 8116 17196
rect 7883 17156 8116 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10459 17156 10609 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11054 17184 11060 17196
rect 10919 17156 11060 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 6938 17088 7420 17116
rect 6938 17085 6950 17088
rect 6892 17079 6950 17085
rect 4985 17051 5043 17057
rect 4985 17048 4997 17051
rect 4126 17020 4997 17048
rect 4985 17017 4997 17020
rect 5031 17048 5043 17051
rect 5350 17048 5356 17060
rect 5031 17020 5356 17048
rect 5031 17017 5043 17020
rect 4985 17011 5043 17017
rect 5350 17008 5356 17020
rect 5408 17048 5414 17060
rect 5813 17051 5871 17057
rect 5813 17048 5825 17051
rect 5408 17020 5825 17048
rect 5408 17008 5414 17020
rect 5813 17017 5825 17020
rect 5859 17017 5871 17051
rect 5813 17011 5871 17017
rect 6362 17008 6368 17060
rect 6420 17048 6426 17060
rect 6641 17051 6699 17057
rect 6641 17048 6653 17051
rect 6420 17020 6653 17048
rect 6420 17008 6426 17020
rect 6641 17017 6653 17020
rect 6687 17048 6699 17051
rect 7742 17048 7748 17060
rect 6687 17020 7748 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 7742 17008 7748 17020
rect 7800 17048 7806 17060
rect 8199 17051 8257 17057
rect 8199 17048 8211 17051
rect 7800 17020 8211 17048
rect 7800 17008 7806 17020
rect 8199 17017 8211 17020
rect 8245 17048 8257 17051
rect 8662 17048 8668 17060
rect 8245 17020 8668 17048
rect 8245 17017 8257 17020
rect 8199 17011 8257 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 10612 17048 10640 17147
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11974 17184 11980 17196
rect 11563 17156 11980 17184
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12590 17125 12618 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14550 17320 14556 17332
rect 14507 17292 14556 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 14366 17252 14372 17264
rect 14056 17224 14372 17252
rect 14056 17212 14062 17224
rect 14366 17212 14372 17224
rect 14424 17252 14430 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 14424 17224 14749 17252
rect 14424 17212 14430 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 24762 17252 24768 17264
rect 24723 17224 24768 17252
rect 14737 17215 14795 17221
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 16298 17184 16304 17196
rect 16259 17156 16304 17184
rect 16298 17144 16304 17156
rect 16356 17184 16362 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 16356 17156 17233 17184
rect 16356 17144 16362 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 12575 17119 12633 17125
rect 12575 17085 12587 17119
rect 12621 17085 12633 17119
rect 12575 17079 12633 17085
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13541 17119 13599 17125
rect 13541 17116 13553 17119
rect 13228 17088 13553 17116
rect 13228 17076 13234 17088
rect 13541 17085 13553 17088
rect 13587 17085 13599 17119
rect 13541 17079 13599 17085
rect 13786 17088 13952 17116
rect 10686 17048 10692 17060
rect 10599 17020 10692 17048
rect 10686 17008 10692 17020
rect 10744 17048 10750 17060
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 10744 17020 10977 17048
rect 10744 17008 10750 17020
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 12250 17048 12256 17060
rect 12163 17020 12256 17048
rect 10965 17011 11023 17017
rect 12250 17008 12256 17020
rect 12308 17048 12314 17060
rect 13630 17048 13636 17060
rect 12308 17020 13636 17048
rect 12308 17008 12314 17020
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 106 16940 112 16992
rect 164 16980 170 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 164 16952 1593 16980
rect 164 16940 170 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 1949 16983 2007 16989
rect 1949 16980 1961 16983
rect 1728 16952 1961 16980
rect 1728 16940 1734 16952
rect 1949 16949 1961 16952
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 2498 16980 2504 16992
rect 2096 16952 2504 16980
rect 2096 16940 2102 16952
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 6178 16980 6184 16992
rect 6139 16952 6184 16980
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6963 16983 7021 16989
rect 6963 16949 6975 16983
rect 7009 16980 7021 16983
rect 7098 16980 7104 16992
rect 7009 16952 7104 16980
rect 7009 16949 7021 16952
rect 6963 16943 7021 16949
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 9769 16983 9827 16989
rect 9769 16949 9781 16983
rect 9815 16980 9827 16983
rect 11422 16980 11428 16992
rect 9815 16952 11428 16980
rect 9815 16949 9827 16952
rect 9769 16943 9827 16949
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 11790 16980 11796 16992
rect 11751 16952 11796 16980
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 12667 16983 12725 16989
rect 12667 16949 12679 16983
rect 12713 16980 12725 16983
rect 12894 16980 12900 16992
rect 12713 16952 12900 16980
rect 12713 16949 12725 16952
rect 12667 16943 12725 16949
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13354 16980 13360 16992
rect 13315 16952 13360 16980
rect 13354 16940 13360 16952
rect 13412 16980 13418 16992
rect 13786 16980 13814 17088
rect 13924 17057 13952 17088
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 15286 17116 15292 17128
rect 14056 17088 15292 17116
rect 14056 17076 14062 17088
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24268 17088 24593 17116
rect 24268 17076 24274 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 13903 17051 13961 17057
rect 13903 17017 13915 17051
rect 13949 17017 13961 17051
rect 13903 17011 13961 17017
rect 16390 17008 16396 17060
rect 16448 17048 16454 17060
rect 16942 17048 16948 17060
rect 16448 17020 16493 17048
rect 16903 17020 16948 17048
rect 16448 17008 16454 17020
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 15378 16980 15384 16992
rect 13412 16952 13814 16980
rect 15339 16952 15384 16980
rect 13412 16940 13418 16952
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15620 16952 15669 16980
rect 15620 16940 15626 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 16117 16983 16175 16989
rect 16117 16949 16129 16983
rect 16163 16980 16175 16983
rect 16408 16980 16436 17008
rect 16163 16952 16436 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1535 16779 1593 16785
rect 1535 16745 1547 16779
rect 1581 16776 1593 16779
rect 1762 16776 1768 16788
rect 1581 16748 1768 16776
rect 1581 16745 1593 16748
rect 1535 16739 1593 16745
rect 1762 16736 1768 16748
rect 1820 16776 1826 16788
rect 2314 16776 2320 16788
rect 1820 16748 2320 16776
rect 1820 16736 1826 16748
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 5258 16736 5264 16788
rect 5316 16776 5322 16788
rect 5353 16779 5411 16785
rect 5353 16776 5365 16779
rect 5316 16748 5365 16776
rect 5316 16736 5322 16748
rect 5353 16745 5365 16748
rect 5399 16745 5411 16779
rect 5353 16739 5411 16745
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5592 16748 5641 16776
rect 5592 16736 5598 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 5629 16739 5687 16745
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 10008 16748 10057 16776
rect 10008 16736 10014 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 10045 16739 10103 16745
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16776 10655 16779
rect 11790 16776 11796 16788
rect 10643 16748 11796 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 14642 16776 14648 16788
rect 14603 16748 14648 16776
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 4798 16717 4804 16720
rect 4795 16708 4804 16717
rect 4711 16680 4804 16708
rect 4795 16671 4804 16680
rect 4856 16708 4862 16720
rect 6362 16708 6368 16720
rect 4856 16680 6368 16708
rect 4798 16668 4804 16671
rect 4856 16668 4862 16680
rect 6362 16668 6368 16680
rect 6420 16668 6426 16720
rect 7193 16711 7251 16717
rect 7193 16677 7205 16711
rect 7239 16708 7251 16711
rect 9398 16708 9404 16720
rect 7239 16680 9404 16708
rect 7239 16677 7251 16680
rect 7193 16671 7251 16677
rect 9398 16668 9404 16680
rect 9456 16708 9462 16720
rect 12250 16708 12256 16720
rect 9456 16680 9720 16708
rect 12211 16680 12256 16708
rect 9456 16668 9462 16680
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1854 16640 1860 16652
rect 1510 16612 1860 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2498 16640 2504 16652
rect 2459 16612 2504 16640
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2924 16612 2973 16640
rect 2924 16600 2930 16612
rect 2961 16609 2973 16612
rect 3007 16640 3019 16643
rect 6086 16640 6092 16652
rect 3007 16612 6092 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6454 16640 6460 16652
rect 6415 16612 6460 16640
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16609 6975 16643
rect 8294 16640 8300 16652
rect 8255 16612 8300 16640
rect 6917 16603 6975 16609
rect 3142 16572 3148 16584
rect 3103 16544 3148 16572
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16572 4491 16575
rect 5534 16572 5540 16584
rect 4479 16544 5540 16572
rect 4479 16541 4491 16544
rect 4433 16535 4491 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 6104 16572 6132 16600
rect 6932 16572 6960 16603
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 9692 16649 9720 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12894 16668 12900 16720
rect 12952 16708 12958 16720
rect 13722 16708 13728 16720
rect 12952 16680 13728 16708
rect 12952 16668 12958 16680
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 13817 16711 13875 16717
rect 13817 16677 13829 16711
rect 13863 16708 13875 16711
rect 14182 16708 14188 16720
rect 13863 16680 14188 16708
rect 13863 16677 13875 16680
rect 13817 16671 13875 16677
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 14369 16711 14427 16717
rect 14369 16677 14381 16711
rect 14415 16708 14427 16711
rect 14734 16708 14740 16720
rect 14415 16680 14740 16708
rect 14415 16677 14427 16680
rect 14369 16671 14427 16677
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 6104 16544 7481 16572
rect 7469 16541 7481 16544
rect 7515 16572 7527 16575
rect 7650 16572 7656 16584
rect 7515 16544 7656 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7650 16532 7656 16544
rect 7708 16572 7714 16584
rect 8496 16572 8524 16603
rect 7708 16544 8524 16572
rect 8757 16575 8815 16581
rect 7708 16532 7714 16544
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 9490 16572 9496 16584
rect 8803 16544 9496 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 12158 16572 12164 16584
rect 12119 16544 12164 16572
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12713 16507 12771 16513
rect 12713 16473 12725 16507
rect 12759 16504 12771 16507
rect 14384 16504 14412 16671
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 15654 16668 15660 16720
rect 15712 16708 15718 16720
rect 16162 16711 16220 16717
rect 16162 16708 16174 16711
rect 15712 16680 16174 16708
rect 15712 16668 15718 16680
rect 16162 16677 16174 16680
rect 16208 16677 16220 16711
rect 17770 16708 17776 16720
rect 17731 16680 17776 16708
rect 16162 16671 16220 16677
rect 17770 16668 17776 16680
rect 17828 16668 17834 16720
rect 15838 16640 15844 16652
rect 15799 16612 15844 16640
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 24118 16600 24124 16652
rect 24176 16640 24182 16652
rect 24581 16643 24639 16649
rect 24581 16640 24593 16643
rect 24176 16612 24593 16640
rect 24176 16600 24182 16612
rect 24581 16609 24593 16612
rect 24627 16609 24639 16643
rect 24581 16603 24639 16609
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 17037 16575 17095 16581
rect 17037 16572 17049 16575
rect 16356 16544 17049 16572
rect 16356 16532 16362 16544
rect 17037 16541 17049 16544
rect 17083 16541 17095 16575
rect 17678 16572 17684 16584
rect 17639 16544 17684 16572
rect 17037 16535 17095 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 12759 16476 14412 16504
rect 18233 16507 18291 16513
rect 12759 16473 12771 16476
rect 12713 16467 12771 16473
rect 18233 16473 18245 16507
rect 18279 16473 18291 16507
rect 18233 16467 18291 16473
rect 1854 16436 1860 16448
rect 1815 16408 1860 16436
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 2314 16436 2320 16448
rect 2275 16408 2320 16436
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 3418 16436 3424 16448
rect 3379 16408 3424 16436
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 4341 16439 4399 16445
rect 4341 16405 4353 16439
rect 4387 16436 4399 16439
rect 4430 16436 4436 16448
rect 4387 16408 4436 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8110 16436 8116 16448
rect 7975 16408 8116 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 10873 16439 10931 16445
rect 10873 16436 10885 16439
rect 10836 16408 10885 16436
rect 10836 16396 10842 16408
rect 10873 16405 10885 16408
rect 10919 16405 10931 16439
rect 13170 16436 13176 16448
rect 13131 16408 13176 16436
rect 10873 16399 10931 16405
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13446 16436 13452 16448
rect 13407 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 14182 16396 14188 16448
rect 14240 16436 14246 16448
rect 15746 16436 15752 16448
rect 14240 16408 15752 16436
rect 14240 16396 14246 16408
rect 15746 16396 15752 16408
rect 15804 16436 15810 16448
rect 16761 16439 16819 16445
rect 16761 16436 16773 16439
rect 15804 16408 16773 16436
rect 15804 16396 15810 16408
rect 16761 16405 16773 16408
rect 16807 16405 16819 16439
rect 16761 16399 16819 16405
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 18248 16436 18276 16467
rect 18506 16436 18512 16448
rect 17000 16408 18512 16436
rect 17000 16396 17006 16408
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 24765 16439 24823 16445
rect 24765 16405 24777 16439
rect 24811 16436 24823 16439
rect 27614 16436 27620 16448
rect 24811 16408 27620 16436
rect 24811 16405 24823 16408
rect 24765 16399 24823 16405
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3878 16232 3884 16244
rect 3839 16204 3884 16232
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 6086 16232 6092 16244
rect 6047 16204 6092 16232
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 9677 16235 9735 16241
rect 9677 16201 9689 16235
rect 9723 16232 9735 16235
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 9723 16204 10609 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 10597 16201 10609 16204
rect 10643 16232 10655 16235
rect 10686 16232 10692 16244
rect 10643 16204 10692 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11793 16235 11851 16241
rect 11793 16201 11805 16235
rect 11839 16232 11851 16235
rect 12158 16232 12164 16244
rect 11839 16204 12164 16232
rect 11839 16201 11851 16204
rect 11793 16195 11851 16201
rect 12158 16192 12164 16204
rect 12216 16232 12222 16244
rect 12575 16235 12633 16241
rect 12575 16232 12587 16235
rect 12216 16204 12587 16232
rect 12216 16192 12222 16204
rect 12575 16201 12587 16204
rect 12621 16201 12633 16235
rect 12575 16195 12633 16201
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 13780 16204 15025 16232
rect 13780 16192 13786 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 15473 16235 15531 16241
rect 15473 16201 15485 16235
rect 15519 16232 15531 16235
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15519 16204 15761 16232
rect 15519 16201 15531 16204
rect 15473 16195 15531 16201
rect 15749 16201 15761 16204
rect 15795 16232 15807 16235
rect 15930 16232 15936 16244
rect 15795 16204 15936 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 17770 16232 17776 16244
rect 17727 16204 17776 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24581 16235 24639 16241
rect 24581 16232 24593 16235
rect 24176 16204 24593 16232
rect 24176 16192 24182 16204
rect 24581 16201 24593 16204
rect 24627 16201 24639 16235
rect 24581 16195 24639 16201
rect 3605 16167 3663 16173
rect 3605 16133 3617 16167
rect 3651 16164 3663 16167
rect 4614 16164 4620 16176
rect 3651 16136 4620 16164
rect 3651 16133 3663 16136
rect 3605 16127 3663 16133
rect 4614 16124 4620 16136
rect 4672 16124 4678 16176
rect 9950 16124 9956 16176
rect 10008 16164 10014 16176
rect 13265 16167 13323 16173
rect 13265 16164 13277 16167
rect 10008 16136 13277 16164
rect 10008 16124 10014 16136
rect 13265 16133 13277 16136
rect 13311 16164 13323 16167
rect 13354 16164 13360 16176
rect 13311 16136 13360 16164
rect 13311 16133 13323 16136
rect 13265 16127 13323 16133
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 18046 16164 18052 16176
rect 13464 16136 18052 16164
rect 13464 16108 13492 16136
rect 18046 16124 18052 16136
rect 18104 16124 18110 16176
rect 3142 16056 3148 16108
rect 3200 16096 3206 16108
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 3200 16068 8769 16096
rect 3200 16056 3206 16068
rect 8757 16065 8769 16068
rect 8803 16096 8815 16099
rect 9030 16096 9036 16108
rect 8803 16068 9036 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 10962 16096 10968 16108
rect 10612 16068 10968 16096
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 2314 16028 2320 16040
rect 2087 16000 2320 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3384 16000 3433 16028
rect 3384 15988 3390 16000
rect 3421 15997 3433 16000
rect 3467 16028 3479 16031
rect 3878 16028 3884 16040
rect 3467 16000 3884 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 4430 16028 4436 16040
rect 4391 16000 4436 16028
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 16028 7159 16031
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 7147 16000 7205 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 7193 15997 7205 16000
rect 7239 15997 7251 16031
rect 7650 16028 7656 16040
rect 7611 16000 7656 16028
rect 7193 15991 7251 15997
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 6454 15960 6460 15972
rect 5132 15932 6460 15960
rect 5132 15920 5138 15932
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 7208 15960 7236 15991
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 10612 16028 10640 16068
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11425 16099 11483 16105
rect 11425 16065 11437 16099
rect 11471 16096 11483 16099
rect 11698 16096 11704 16108
rect 11471 16068 11704 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12250 16096 12256 16108
rect 12207 16068 12256 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12250 16056 12256 16068
rect 12308 16096 12314 16108
rect 13446 16096 13452 16108
rect 12308 16068 12756 16096
rect 13407 16068 13452 16096
rect 12308 16056 12314 16068
rect 7852 16000 10640 16028
rect 7852 15960 7880 16000
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12472 16031 12530 16037
rect 12472 16028 12484 16031
rect 12400 16000 12484 16028
rect 12400 15988 12406 16000
rect 12472 15997 12484 16000
rect 12518 15997 12530 16031
rect 12728 16028 12756 16068
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 15335 16099 15393 16105
rect 15335 16096 15347 16099
rect 13688 16068 15347 16096
rect 13688 16056 13694 16068
rect 15335 16065 15347 16068
rect 15381 16065 15393 16099
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 15335 16059 15393 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 14366 16028 14372 16040
rect 12728 16000 14372 16028
rect 12472 15991 12530 15997
rect 7208 15932 7880 15960
rect 7929 15963 7987 15969
rect 7929 15929 7941 15963
rect 7975 15960 7987 15963
rect 8938 15960 8944 15972
rect 7975 15932 8944 15960
rect 7975 15929 7987 15932
rect 7929 15923 7987 15929
rect 8938 15920 8944 15932
rect 8996 15920 9002 15972
rect 9119 15963 9177 15969
rect 9119 15929 9131 15963
rect 9165 15960 9177 15963
rect 10778 15960 10784 15972
rect 9165 15932 9674 15960
rect 10739 15932 10784 15960
rect 9165 15929 9177 15932
rect 9119 15923 9177 15929
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2498 15892 2504 15904
rect 2459 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 3234 15892 3240 15904
rect 3195 15864 3240 15892
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15892 4399 15895
rect 4798 15892 4804 15904
rect 4387 15864 4804 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 5629 15895 5687 15901
rect 5629 15892 5641 15895
rect 5592 15864 5641 15892
rect 5592 15852 5598 15864
rect 5629 15861 5641 15864
rect 5675 15861 5687 15895
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 5629 15855 5687 15861
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8662 15892 8668 15904
rect 8575 15864 8668 15892
rect 8662 15852 8668 15864
rect 8720 15892 8726 15904
rect 9134 15892 9162 15923
rect 8720 15864 9162 15892
rect 9646 15892 9674 15932
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 10873 15963 10931 15969
rect 10873 15929 10885 15963
rect 10919 15929 10931 15963
rect 12487 15960 12515 15991
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15248 16031 15306 16037
rect 15248 16028 15260 16031
rect 15160 16000 15260 16028
rect 15160 15988 15166 16000
rect 15248 15997 15260 16000
rect 15294 16028 15306 16031
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15294 16000 15485 16028
rect 15294 15997 15306 16000
rect 15248 15991 15306 15997
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 18100 16031 18158 16037
rect 18100 15997 18112 16031
rect 18146 16028 18158 16031
rect 18506 16028 18512 16040
rect 18146 16000 18512 16028
rect 18146 15997 18158 16000
rect 18100 15991 18158 15997
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 12487 15932 12909 15960
rect 10873 15923 10931 15929
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 9950 15892 9956 15904
rect 9646 15864 9956 15892
rect 8720 15852 8726 15864
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10888 15892 10916 15923
rect 13354 15920 13360 15972
rect 13412 15960 13418 15972
rect 13770 15963 13828 15969
rect 13770 15960 13782 15963
rect 13412 15932 13782 15960
rect 13412 15920 13418 15932
rect 13770 15929 13782 15932
rect 13816 15960 13828 15963
rect 14090 15960 14096 15972
rect 13816 15932 14096 15960
rect 13816 15929 13828 15932
rect 13770 15923 13828 15929
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 14182 15920 14188 15972
rect 14240 15960 14246 15972
rect 14645 15963 14703 15969
rect 14645 15960 14657 15963
rect 14240 15932 14657 15960
rect 14240 15920 14246 15932
rect 14645 15929 14657 15932
rect 14691 15929 14703 15963
rect 14645 15923 14703 15929
rect 14734 15920 14740 15972
rect 14792 15960 14798 15972
rect 16298 15960 16304 15972
rect 14792 15932 16304 15960
rect 14792 15920 14798 15932
rect 16298 15920 16304 15932
rect 16356 15920 16362 15972
rect 16393 15963 16451 15969
rect 16393 15929 16405 15963
rect 16439 15929 16451 15963
rect 16393 15923 16451 15929
rect 18187 15963 18245 15969
rect 18187 15929 18199 15963
rect 18233 15960 18245 15963
rect 18782 15960 18788 15972
rect 18233 15932 18788 15960
rect 18233 15929 18245 15932
rect 18187 15923 18245 15929
rect 10744 15864 10916 15892
rect 10744 15852 10750 15864
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15712 15864 16037 15892
rect 15712 15852 15718 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16408 15892 16436 15923
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 16574 15892 16580 15904
rect 16408 15864 16580 15892
rect 16025 15855 16083 15861
rect 16574 15852 16580 15864
rect 16632 15892 16638 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 16632 15864 17233 15892
rect 16632 15852 16638 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4488 15660 4721 15688
rect 4488 15648 4494 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 4709 15651 4767 15657
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 9030 15688 9036 15700
rect 8991 15660 9036 15688
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10008 15660 10317 15688
rect 10008 15648 10014 15660
rect 1670 15620 1676 15632
rect 1631 15592 1676 15620
rect 1670 15580 1676 15592
rect 1728 15580 1734 15632
rect 2225 15623 2283 15629
rect 2225 15589 2237 15623
rect 2271 15620 2283 15623
rect 2406 15620 2412 15632
rect 2271 15592 2412 15620
rect 2271 15589 2283 15592
rect 2225 15583 2283 15589
rect 2406 15580 2412 15592
rect 2464 15620 2470 15632
rect 3786 15620 3792 15632
rect 2464 15592 3792 15620
rect 2464 15580 2470 15592
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 4525 15623 4583 15629
rect 4525 15589 4537 15623
rect 4571 15620 4583 15623
rect 4798 15620 4804 15632
rect 4571 15592 4804 15620
rect 4571 15589 4583 15592
rect 4525 15583 4583 15589
rect 4798 15580 4804 15592
rect 4856 15580 4862 15632
rect 6840 15620 6868 15648
rect 5276 15592 7420 15620
rect 4614 15552 4620 15564
rect 4575 15524 4620 15552
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 5276 15561 5304 15592
rect 7392 15564 7420 15592
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 8665 15623 8723 15629
rect 8665 15620 8677 15623
rect 7708 15592 8677 15620
rect 7708 15580 7714 15592
rect 8665 15589 8677 15592
rect 8711 15589 8723 15623
rect 9122 15620 9128 15632
rect 8665 15583 8723 15589
rect 8772 15592 9128 15620
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5224 15524 5273 15552
rect 5224 15512 5230 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 5350 15512 5356 15564
rect 5408 15552 5414 15564
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 5408 15524 5457 15552
rect 5408 15512 5414 15524
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6043 15524 6500 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 3418 15484 3424 15496
rect 1627 15456 3424 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 3881 15419 3939 15425
rect 3881 15385 3893 15419
rect 3927 15416 3939 15419
rect 4982 15416 4988 15428
rect 3927 15388 4988 15416
rect 3927 15385 3939 15388
rect 3881 15379 3939 15385
rect 4982 15376 4988 15388
rect 5040 15416 5046 15428
rect 6012 15416 6040 15515
rect 6472 15425 6500 15524
rect 6822 15512 6828 15564
rect 6880 15552 6886 15564
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 6880 15524 6929 15552
rect 6880 15512 6886 15524
rect 6917 15521 6929 15524
rect 6963 15521 6975 15555
rect 7374 15552 7380 15564
rect 7287 15524 7380 15552
rect 6917 15515 6975 15521
rect 7374 15512 7380 15524
rect 7432 15512 7438 15564
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 7616 15524 7757 15552
rect 7616 15512 7622 15524
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 8343 15524 8493 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8481 15521 8493 15524
rect 8527 15552 8539 15555
rect 8772 15552 8800 15592
rect 9122 15580 9128 15592
rect 9180 15580 9186 15632
rect 10289 15629 10317 15660
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11020 15660 12480 15688
rect 11020 15648 11026 15660
rect 10274 15623 10332 15629
rect 10274 15589 10286 15623
rect 10320 15589 10332 15623
rect 10274 15583 10332 15589
rect 11790 15580 11796 15632
rect 11848 15620 11854 15632
rect 11885 15623 11943 15629
rect 11885 15620 11897 15623
rect 11848 15592 11897 15620
rect 11848 15580 11854 15592
rect 11885 15589 11897 15592
rect 11931 15589 11943 15623
rect 11885 15583 11943 15589
rect 8527 15524 8800 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 9858 15552 9864 15564
rect 8996 15524 9864 15552
rect 8996 15512 9002 15524
rect 9858 15512 9864 15524
rect 9916 15552 9922 15564
rect 9953 15555 10011 15561
rect 9953 15552 9965 15555
rect 9916 15524 9965 15552
rect 9916 15512 9922 15524
rect 9953 15521 9965 15524
rect 9999 15521 10011 15555
rect 12452 15552 12480 15660
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13357 15691 13415 15697
rect 13357 15688 13369 15691
rect 13228 15660 13369 15688
rect 13228 15648 13234 15660
rect 13357 15657 13369 15660
rect 13403 15657 13415 15691
rect 15838 15688 15844 15700
rect 15799 15660 15844 15688
rect 13357 15651 13415 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17770 15688 17776 15700
rect 17175 15660 17776 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17770 15648 17776 15660
rect 17828 15648 17834 15700
rect 18046 15688 18052 15700
rect 18007 15660 18052 15688
rect 18046 15648 18052 15660
rect 18104 15648 18110 15700
rect 15654 15580 15660 15632
rect 15712 15620 15718 15632
rect 16530 15623 16588 15629
rect 16530 15620 16542 15623
rect 15712 15592 16542 15620
rect 15712 15580 15718 15592
rect 16530 15589 16542 15592
rect 16576 15589 16588 15623
rect 17678 15620 17684 15632
rect 17639 15592 17684 15620
rect 16530 15583 16588 15589
rect 17678 15580 17684 15592
rect 17736 15580 17742 15632
rect 13262 15552 13268 15564
rect 12452 15524 13268 15552
rect 9953 15515 10011 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 13872 15524 14289 15552
rect 13872 15512 13878 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 17954 15552 17960 15564
rect 17915 15524 17960 15552
rect 14277 15515 14335 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 18417 15555 18475 15561
rect 18417 15521 18429 15555
rect 18463 15521 18475 15555
rect 18417 15515 18475 15521
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 11606 15484 11612 15496
rect 7156 15456 11612 15484
rect 7156 15444 7162 15456
rect 11606 15444 11612 15456
rect 11664 15484 11670 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11664 15456 11805 15484
rect 11664 15444 11670 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15484 16267 15487
rect 16850 15484 16856 15496
rect 16255 15456 16856 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 5040 15388 6040 15416
rect 6457 15419 6515 15425
rect 5040 15376 5046 15388
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 8481 15419 8539 15425
rect 8481 15416 8493 15419
rect 6503 15388 8493 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 8481 15385 8493 15388
rect 8527 15385 8539 15419
rect 8481 15379 8539 15385
rect 10134 15376 10140 15428
rect 10192 15416 10198 15428
rect 11149 15419 11207 15425
rect 11149 15416 11161 15419
rect 10192 15388 11161 15416
rect 10192 15376 10198 15388
rect 11149 15385 11161 15388
rect 11195 15385 11207 15419
rect 11149 15379 11207 15385
rect 11698 15376 11704 15428
rect 11756 15416 11762 15428
rect 12084 15416 12112 15447
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 17862 15444 17868 15496
rect 17920 15484 17926 15496
rect 18432 15484 18460 15515
rect 17920 15456 18460 15484
rect 17920 15444 17926 15456
rect 13446 15416 13452 15428
rect 11756 15388 13452 15416
rect 11756 15376 11762 15388
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 2590 15348 2596 15360
rect 2551 15320 2596 15348
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2740 15320 2881 15348
rect 2740 15308 2746 15320
rect 2869 15317 2881 15320
rect 2915 15348 2927 15351
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 2915 15320 3433 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 10870 15348 10876 15360
rect 10831 15320 10876 15348
rect 3421 15311 3479 15317
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 12710 15348 12716 15360
rect 12671 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1544 15116 1593 15144
rect 1544 15104 1550 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1728 15116 1961 15144
rect 1728 15104 1734 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 4341 15147 4399 15153
rect 4341 15113 4353 15147
rect 4387 15144 4399 15147
rect 4614 15144 4620 15156
rect 4387 15116 4620 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 9539 15147 9597 15153
rect 9539 15113 9551 15147
rect 9585 15144 9597 15147
rect 10778 15144 10784 15156
rect 9585 15116 10784 15144
rect 9585 15113 9597 15116
rect 9539 15107 9597 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13320 15116 13461 15144
rect 13320 15104 13326 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 14148 15116 15485 15144
rect 14148 15104 14154 15116
rect 15473 15113 15485 15116
rect 15519 15144 15531 15147
rect 15654 15144 15660 15156
rect 15519 15116 15660 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 16577 15147 16635 15153
rect 16577 15144 16589 15147
rect 16448 15116 16589 15144
rect 16448 15104 16454 15116
rect 16577 15113 16589 15116
rect 16623 15113 16635 15147
rect 17494 15144 17500 15156
rect 17407 15116 17500 15144
rect 16577 15107 16635 15113
rect 17494 15104 17500 15116
rect 17552 15144 17558 15156
rect 17954 15144 17960 15156
rect 17552 15116 17960 15144
rect 17552 15104 17558 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 22094 15144 22100 15156
rect 20211 15116 22100 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 3142 15076 3148 15088
rect 3103 15048 3148 15076
rect 3142 15036 3148 15048
rect 3200 15036 3206 15088
rect 5534 15036 5540 15088
rect 5592 15076 5598 15088
rect 5813 15079 5871 15085
rect 5813 15076 5825 15079
rect 5592 15048 5825 15076
rect 5592 15036 5598 15048
rect 5813 15045 5825 15048
rect 5859 15045 5871 15079
rect 5813 15039 5871 15045
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 8205 15079 8263 15085
rect 8205 15076 8217 15079
rect 7984 15048 8217 15076
rect 7984 15036 7990 15048
rect 8205 15045 8217 15048
rect 8251 15045 8263 15079
rect 8205 15039 8263 15045
rect 9309 15079 9367 15085
rect 9309 15045 9321 15079
rect 9355 15076 9367 15079
rect 9950 15076 9956 15088
rect 9355 15048 9956 15076
rect 9355 15045 9367 15048
rect 9309 15039 9367 15045
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 11940 15048 12848 15076
rect 11940 15036 11946 15048
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2464 14980 2605 15008
rect 2464 14968 2470 14980
rect 2593 14977 2605 14980
rect 2639 14977 2651 15011
rect 8018 15008 8024 15020
rect 2593 14971 2651 14977
rect 7392 14980 8024 15008
rect 7392 14952 7420 14980
rect 8018 14968 8024 14980
rect 8076 15008 8082 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8076 14980 8585 15008
rect 8076 14968 8082 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 12342 15008 12348 15020
rect 8573 14971 8631 14977
rect 9876 14980 12348 15008
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 4614 14940 4620 14952
rect 4575 14912 4620 14940
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5166 14940 5172 14952
rect 5127 14912 5172 14940
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5810 14940 5816 14952
rect 5316 14912 5361 14940
rect 5771 14912 5816 14940
rect 5316 14900 5322 14912
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7374 14940 7380 14952
rect 7335 14912 7380 14940
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 7616 14912 7665 14940
rect 7616 14900 7622 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 8202 14940 8208 14952
rect 8163 14912 8208 14940
rect 7653 14903 7711 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9876 14949 9904 14980
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12710 15008 12716 15020
rect 12575 14980 12716 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12820 15017 12848 15048
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 15562 15008 15568 15020
rect 13780 14980 15568 15008
rect 13780 14968 13786 14980
rect 9436 14943 9494 14949
rect 9436 14940 9448 14943
rect 9324 14912 9448 14940
rect 2682 14832 2688 14884
rect 2740 14872 2746 14884
rect 3973 14875 4031 14881
rect 2740 14844 2785 14872
rect 2740 14832 2746 14844
rect 3973 14841 3985 14875
rect 4019 14872 4031 14875
rect 4338 14872 4344 14884
rect 4019 14844 4344 14872
rect 4019 14841 4031 14844
rect 3973 14835 4031 14841
rect 4338 14832 4344 14844
rect 4396 14872 4402 14884
rect 5184 14872 5212 14900
rect 4396 14844 5212 14872
rect 4396 14832 4402 14844
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 9324 14872 9352 14912
rect 9436 14909 9448 14912
rect 9482 14940 9494 14943
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9482 14912 9873 14940
rect 9482 14909 9494 14912
rect 9436 14903 9494 14909
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 14568 14949 14596 14980
rect 15562 14968 15568 14980
rect 15620 15008 15626 15020
rect 15620 14980 15884 15008
rect 15620 14968 15626 14980
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 10192 14912 10425 14940
rect 10192 14900 10198 14912
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 14001 14943 14059 14949
rect 14001 14940 14013 14943
rect 10413 14903 10471 14909
rect 13786 14912 14013 14940
rect 7524 14844 9352 14872
rect 10734 14875 10792 14881
rect 7524 14832 7530 14844
rect 10734 14841 10746 14875
rect 10780 14841 10792 14875
rect 10734 14835 10792 14841
rect 2314 14804 2320 14816
rect 2275 14776 2320 14804
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 4856 14776 6193 14804
rect 4856 14764 4862 14776
rect 6181 14773 6193 14776
rect 6227 14804 6239 14807
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6227 14776 6561 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 7558 14804 7564 14816
rect 6595 14776 7564 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10008 14776 10241 14804
rect 10008 14764 10014 14776
rect 10229 14773 10241 14776
rect 10275 14804 10287 14807
rect 10749 14804 10777 14835
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 12253 14875 12311 14881
rect 12253 14872 12265 14875
rect 10928 14844 12265 14872
rect 10928 14832 10934 14844
rect 12253 14841 12265 14844
rect 12299 14872 12311 14875
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 12299 14844 12633 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12621 14841 12633 14844
rect 12667 14841 12679 14875
rect 12621 14835 12679 14841
rect 11330 14804 11336 14816
rect 10275 14776 10777 14804
rect 11291 14776 11336 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 13786 14804 13814 14912
rect 14001 14909 14013 14912
rect 14047 14940 14059 14943
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 14047 14912 14105 14940
rect 14047 14909 14059 14912
rect 14001 14903 14059 14909
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14909 14611 14943
rect 14553 14903 14611 14909
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15856 14940 15884 14980
rect 15930 14968 15936 15020
rect 15988 15008 15994 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 15988 14980 17785 15008
rect 15988 14968 15994 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 16482 14940 16488 14952
rect 15856 14912 16488 14940
rect 15657 14903 15715 14909
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14872 14887 14875
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14875 14844 15117 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 15105 14841 15117 14844
rect 15151 14872 15163 14875
rect 15672 14872 15700 14903
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 17788 14940 17816 14971
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 21545 15011 21603 15017
rect 21545 15008 21557 15011
rect 19484 14980 21557 15008
rect 19484 14968 19490 14980
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17788 14912 18061 14940
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18506 14940 18512 14952
rect 18467 14912 18512 14940
rect 18049 14903 18107 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 21167 14949 21195 14980
rect 21545 14977 21557 14980
rect 21591 14977 21603 15011
rect 21545 14971 21603 14977
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14940 20039 14943
rect 21152 14943 21210 14949
rect 20027 14912 20668 14940
rect 20027 14909 20039 14912
rect 19981 14903 20039 14909
rect 15151 14844 15700 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 15746 14832 15752 14884
rect 15804 14872 15810 14884
rect 15978 14875 16036 14881
rect 15978 14872 15990 14875
rect 15804 14844 15990 14872
rect 15804 14832 15810 14844
rect 15978 14841 15990 14844
rect 16024 14872 16036 14875
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 16024 14844 16865 14872
rect 16024 14841 16036 14844
rect 15978 14835 16036 14841
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 16853 14835 16911 14841
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 17920 14844 19073 14872
rect 17920 14832 17926 14844
rect 19061 14841 19073 14844
rect 19107 14841 19119 14875
rect 19061 14835 19119 14841
rect 18138 14804 18144 14816
rect 13688 14776 13814 14804
rect 18099 14776 18144 14804
rect 13688 14764 13694 14776
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 20640 14813 20668 14912
rect 21152 14909 21164 14943
rect 21198 14909 21210 14943
rect 21152 14903 21210 14909
rect 20625 14807 20683 14813
rect 20625 14773 20637 14807
rect 20671 14804 20683 14807
rect 20898 14804 20904 14816
rect 20671 14776 20904 14804
rect 20671 14773 20683 14776
rect 20625 14767 20683 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21223 14807 21281 14813
rect 21223 14773 21235 14807
rect 21269 14804 21281 14807
rect 21358 14804 21364 14816
rect 21269 14776 21364 14804
rect 21269 14773 21281 14776
rect 21223 14767 21281 14773
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 4338 14600 4344 14612
rect 4299 14572 4344 14600
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 4614 14600 4620 14612
rect 4575 14572 4620 14600
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 7193 14603 7251 14609
rect 7193 14569 7205 14603
rect 7239 14600 7251 14603
rect 7650 14600 7656 14612
rect 7239 14572 7656 14600
rect 7239 14569 7251 14572
rect 7193 14563 7251 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10008 14572 10272 14600
rect 10008 14560 10014 14572
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2774 14532 2780 14544
rect 2639 14504 2780 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2774 14492 2780 14504
rect 2832 14492 2838 14544
rect 3142 14532 3148 14544
rect 3103 14504 3148 14532
rect 3142 14492 3148 14504
rect 3200 14532 3206 14544
rect 5994 14532 6000 14544
rect 3200 14504 6000 14532
rect 3200 14492 3206 14504
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 7469 14535 7527 14541
rect 7469 14532 7481 14535
rect 6840 14504 7481 14532
rect 6840 14476 6868 14504
rect 7469 14501 7481 14504
rect 7515 14501 7527 14535
rect 7668 14532 7696 14560
rect 10244 14544 10272 14572
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 15565 14603 15623 14609
rect 11388 14572 13584 14600
rect 11388 14560 11394 14572
rect 8202 14532 8208 14544
rect 7668 14504 8208 14532
rect 7469 14495 7527 14501
rect 8202 14492 8208 14504
rect 8260 14532 8266 14544
rect 8757 14535 8815 14541
rect 8260 14504 8524 14532
rect 8260 14492 8266 14504
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4672 14436 5089 14464
rect 4672 14424 4678 14436
rect 5077 14433 5089 14436
rect 5123 14464 5135 14467
rect 6086 14464 6092 14476
rect 5123 14436 6092 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 6086 14424 6092 14436
rect 6144 14464 6150 14476
rect 6822 14464 6828 14476
rect 6144 14436 6828 14464
rect 6144 14424 6150 14436
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7098 14464 7104 14476
rect 7055 14436 7104 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 8496 14473 8524 14504
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 10134 14532 10140 14544
rect 8803 14504 10140 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 10366 14535 10424 14541
rect 10366 14532 10378 14535
rect 10284 14504 10378 14532
rect 10284 14492 10290 14504
rect 10366 14501 10378 14504
rect 10412 14501 10424 14535
rect 11606 14532 11612 14544
rect 11567 14504 11612 14532
rect 10366 14495 10424 14501
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 11974 14532 11980 14544
rect 11935 14504 11980 14532
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13446 14532 13452 14544
rect 13407 14504 13452 14532
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 13556 14541 13584 14572
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 15611 14572 17509 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 13814 14532 13820 14544
rect 13587 14504 13820 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 15672 14473 15700 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 17497 14563 17555 14569
rect 17586 14560 17592 14612
rect 17644 14600 17650 14612
rect 19061 14603 19119 14609
rect 19061 14600 19073 14603
rect 17644 14572 19073 14600
rect 17644 14560 17650 14572
rect 19061 14569 19073 14572
rect 19107 14569 19119 14603
rect 19061 14563 19119 14569
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 20254 14600 20260 14612
rect 19392 14572 20260 14600
rect 19392 14560 19398 14572
rect 20254 14560 20260 14572
rect 20312 14560 20318 14612
rect 15746 14492 15752 14544
rect 15804 14532 15810 14544
rect 15978 14535 16036 14541
rect 15978 14532 15990 14535
rect 15804 14504 15990 14532
rect 15804 14492 15810 14504
rect 15978 14501 15990 14504
rect 16024 14501 16036 14535
rect 16850 14532 16856 14544
rect 16811 14504 16856 14532
rect 15978 14495 16036 14501
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 18506 14492 18512 14544
rect 18564 14532 18570 14544
rect 18564 14504 19472 14532
rect 18564 14492 18570 14504
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14433 15715 14467
rect 16574 14464 16580 14476
rect 16535 14436 16580 14464
rect 15657 14427 15715 14433
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 1443 14368 2237 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2225 14365 2237 14368
rect 2271 14396 2283 14399
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 2271 14368 2513 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5500 14368 5733 14396
rect 5500 14356 5506 14368
rect 5721 14365 5733 14368
rect 5767 14396 5779 14399
rect 6730 14396 6736 14408
rect 5767 14368 6736 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 8312 14396 8340 14427
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 17402 14464 17408 14476
rect 17363 14436 17408 14464
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17862 14464 17868 14476
rect 17823 14436 17868 14464
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 19444 14473 19472 14504
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14464 19487 14467
rect 19794 14464 19800 14476
rect 19475 14436 19800 14464
rect 19475 14433 19487 14436
rect 19429 14427 19487 14433
rect 8662 14396 8668 14408
rect 8312 14368 8668 14396
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 9824 14368 10057 14396
rect 9824 14356 9830 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 11882 14396 11888 14408
rect 11843 14368 11888 14396
rect 10045 14359 10103 14365
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 12161 14359 12219 14365
rect 13556 14368 13737 14396
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 3881 14331 3939 14337
rect 3881 14328 3893 14331
rect 3660 14300 3893 14328
rect 3660 14288 3666 14300
rect 3881 14297 3893 14300
rect 3927 14328 3939 14331
rect 5258 14328 5264 14340
rect 3927 14300 5264 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 5810 14288 5816 14340
rect 5868 14328 5874 14340
rect 6181 14331 6239 14337
rect 6181 14328 6193 14331
rect 5868 14300 6193 14328
rect 5868 14288 5874 14300
rect 6181 14297 6193 14300
rect 6227 14328 6239 14331
rect 6362 14328 6368 14340
rect 6227 14300 6368 14328
rect 6227 14297 6239 14300
rect 6181 14291 6239 14297
rect 6362 14288 6368 14300
rect 6420 14328 6426 14340
rect 8110 14328 8116 14340
rect 6420 14300 8116 14328
rect 6420 14288 6426 14300
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 12176 14328 12204 14359
rect 13556 14328 13584 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 11756 14300 13584 14328
rect 11756 14288 11762 14300
rect 13630 14288 13636 14340
rect 13688 14328 13694 14340
rect 18984 14328 19012 14427
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 21082 14464 21088 14476
rect 21043 14436 21088 14464
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 21818 14396 21824 14408
rect 21775 14368 21824 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 19334 14328 19340 14340
rect 13688 14300 19340 14328
rect 13688 14288 13694 14300
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2222 14260 2228 14272
rect 1995 14232 2228 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 3694 14260 3700 14272
rect 3559 14232 3700 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 3694 14220 3700 14232
rect 3752 14260 3758 14272
rect 4154 14260 4160 14272
rect 3752 14232 4160 14260
rect 3752 14220 3758 14232
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 6546 14260 6552 14272
rect 6507 14232 6552 14260
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 10965 14263 11023 14269
rect 10965 14229 10977 14263
rect 11011 14260 11023 14263
rect 11146 14260 11152 14272
rect 11011 14232 11152 14260
rect 11011 14229 11023 14232
rect 10965 14223 11023 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 12676 14232 13185 14260
rect 12676 14220 12682 14232
rect 13173 14229 13185 14232
rect 13219 14260 13231 14263
rect 13722 14260 13728 14272
rect 13219 14232 13728 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 18417 14263 18475 14269
rect 18417 14260 18429 14263
rect 16172 14232 18429 14260
rect 16172 14220 16178 14232
rect 18417 14229 18429 14232
rect 18463 14260 18475 14263
rect 18506 14260 18512 14272
rect 18463 14232 18512 14260
rect 18463 14229 18475 14232
rect 18417 14223 18475 14229
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 20070 14260 20076 14272
rect 20031 14232 20076 14260
rect 20070 14220 20076 14232
rect 20128 14220 20134 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 6273 14059 6331 14065
rect 6273 14025 6285 14059
rect 6319 14056 6331 14059
rect 7098 14056 7104 14068
rect 6319 14028 7104 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 7098 14016 7104 14028
rect 7156 14056 7162 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 7156 14028 9413 14056
rect 7156 14016 7162 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11563 14028 11897 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11885 14025 11897 14028
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13872 14028 13921 14056
rect 13872 14016 13878 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 17402 14056 17408 14068
rect 15620 14028 17408 14056
rect 15620 14016 15626 14028
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 19794 14056 19800 14068
rect 19755 14028 19800 14056
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20119 14059 20177 14065
rect 20119 14056 20131 14059
rect 20036 14028 20131 14056
rect 20036 14016 20042 14028
rect 20119 14025 20131 14028
rect 20165 14025 20177 14059
rect 20119 14019 20177 14025
rect 20625 14059 20683 14065
rect 20625 14025 20637 14059
rect 20671 14056 20683 14059
rect 20993 14059 21051 14065
rect 20993 14056 21005 14059
rect 20671 14028 21005 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 20993 14025 21005 14028
rect 21039 14056 21051 14059
rect 21082 14056 21088 14068
rect 21039 14028 21088 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 25130 14056 25136 14068
rect 25091 14028 25136 14056
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 3200 13960 3249 13988
rect 3200 13948 3206 13960
rect 3237 13957 3249 13960
rect 3283 13988 3295 13991
rect 3878 13988 3884 14000
rect 3283 13960 3884 13988
rect 3283 13957 3295 13960
rect 3237 13951 3295 13957
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 4154 13948 4160 14000
rect 4212 13988 4218 14000
rect 6641 13991 6699 13997
rect 4212 13960 4660 13988
rect 4212 13948 4218 13960
rect 1489 13923 1547 13929
rect 1489 13889 1501 13923
rect 1535 13920 1547 13923
rect 2590 13920 2596 13932
rect 1535 13892 2596 13920
rect 1535 13889 1547 13892
rect 1489 13883 1547 13889
rect 2590 13880 2596 13892
rect 2648 13920 2654 13932
rect 2648 13892 3280 13920
rect 2648 13880 2654 13892
rect 3252 13852 3280 13892
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3568 13892 4476 13920
rect 3568 13880 3574 13892
rect 3878 13852 3884 13864
rect 3252 13824 3648 13852
rect 3839 13824 3884 13852
rect 1851 13787 1909 13793
rect 1851 13753 1863 13787
rect 1897 13784 1909 13787
rect 1946 13784 1952 13796
rect 1897 13756 1952 13784
rect 1897 13753 1909 13756
rect 1851 13747 1909 13753
rect 1946 13744 1952 13756
rect 2004 13744 2010 13796
rect 2130 13676 2136 13728
rect 2188 13716 2194 13728
rect 2314 13716 2320 13728
rect 2188 13688 2320 13716
rect 2188 13676 2194 13688
rect 2314 13676 2320 13688
rect 2372 13716 2378 13728
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 2372 13688 2421 13716
rect 2372 13676 2378 13688
rect 2409 13685 2421 13688
rect 2455 13685 2467 13719
rect 2774 13716 2780 13728
rect 2735 13688 2780 13716
rect 2409 13679 2467 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 3510 13716 3516 13728
rect 3471 13688 3516 13716
rect 3510 13676 3516 13688
rect 3568 13676 3574 13728
rect 3620 13716 3648 13824
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 4246 13852 4252 13864
rect 4207 13824 4252 13852
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4448 13852 4476 13892
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4448 13824 4537 13852
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4632 13852 4660 13960
rect 6641 13957 6653 13991
rect 6687 13988 6699 13991
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 6687 13960 7972 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 7944 13864 7972 13960
rect 13786 13960 14749 13988
rect 8662 13920 8668 13932
rect 8623 13892 8668 13920
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9122 13920 9128 13932
rect 9079 13892 9128 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 9548 13892 10609 13920
rect 9548 13880 9554 13892
rect 10597 13889 10609 13892
rect 10643 13920 10655 13923
rect 10686 13920 10692 13932
rect 10643 13892 10692 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 11940 13892 12173 13920
rect 11940 13880 11946 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13786 13920 13814 13960
rect 14737 13957 14749 13960
rect 14783 13957 14795 13991
rect 15654 13988 15660 14000
rect 15615 13960 15660 13988
rect 14737 13951 14795 13957
rect 15654 13948 15660 13960
rect 15712 13948 15718 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16040 13960 17049 13988
rect 13228 13892 13814 13920
rect 14292 13892 14596 13920
rect 13228 13880 13234 13892
rect 5077 13855 5135 13861
rect 5077 13852 5089 13855
rect 4632 13824 5089 13852
rect 4525 13815 4583 13821
rect 5077 13821 5089 13824
rect 5123 13852 5135 13855
rect 6362 13852 6368 13864
rect 5123 13824 6368 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6788 13824 6837 13852
rect 6788 13812 6794 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6825 13815 6883 13821
rect 7116 13824 7297 13852
rect 5537 13787 5595 13793
rect 5537 13753 5549 13787
rect 5583 13784 5595 13787
rect 6086 13784 6092 13796
rect 5583 13756 6092 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 7116 13784 7144 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 6604 13756 7144 13784
rect 6604 13744 6610 13756
rect 3789 13719 3847 13725
rect 3789 13716 3801 13719
rect 3620 13688 3801 13716
rect 3789 13685 3801 13688
rect 3835 13685 3847 13719
rect 3789 13679 3847 13685
rect 5258 13676 5264 13728
rect 5316 13716 5322 13728
rect 5813 13719 5871 13725
rect 5813 13716 5825 13719
rect 5316 13688 5825 13716
rect 5316 13676 5322 13688
rect 5813 13685 5825 13688
rect 5859 13685 5871 13719
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 5813 13679 5871 13685
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7760 13716 7788 13815
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7984 13824 8217 13852
rect 7984 13812 7990 13824
rect 8205 13821 8217 13824
rect 8251 13852 8263 13855
rect 8846 13852 8852 13864
rect 8251 13824 8852 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9134 13852 9162 13880
rect 9309 13855 9367 13861
rect 9309 13852 9321 13855
rect 9134 13824 9321 13852
rect 9309 13821 9321 13824
rect 9355 13821 9367 13855
rect 9309 13815 9367 13821
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 9122 13787 9180 13793
rect 9122 13784 9134 13787
rect 9088 13756 9134 13784
rect 9088 13744 9094 13756
rect 9122 13753 9134 13756
rect 9168 13753 9180 13787
rect 9122 13747 9180 13753
rect 10959 13787 11017 13793
rect 10959 13753 10971 13787
rect 11005 13753 11017 13787
rect 10959 13747 11017 13753
rect 10134 13716 10140 13728
rect 7248 13688 7788 13716
rect 10095 13688 10140 13716
rect 7248 13676 7254 13688
rect 10134 13676 10140 13688
rect 10192 13716 10198 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 10192 13688 10425 13716
rect 10192 13676 10198 13688
rect 10413 13685 10425 13688
rect 10459 13716 10471 13719
rect 10980 13716 11008 13747
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 12989 13787 13047 13793
rect 12989 13784 13001 13787
rect 12860 13756 13001 13784
rect 12860 13744 12866 13756
rect 12989 13753 13001 13756
rect 13035 13753 13047 13787
rect 12989 13747 13047 13753
rect 13081 13787 13139 13793
rect 13081 13753 13093 13787
rect 13127 13753 13139 13787
rect 13081 13747 13139 13753
rect 13633 13787 13691 13793
rect 13633 13753 13645 13787
rect 13679 13784 13691 13787
rect 13722 13784 13728 13796
rect 13679 13756 13728 13784
rect 13679 13753 13691 13756
rect 13633 13747 13691 13753
rect 10459 13688 11008 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12713 13719 12771 13725
rect 12713 13716 12725 13719
rect 11664 13688 12725 13716
rect 11664 13676 11670 13688
rect 12713 13685 12725 13688
rect 12759 13716 12771 13719
rect 13096 13716 13124 13747
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 14292 13793 14320 13892
rect 14568 13861 14596 13892
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 15930 13812 15936 13864
rect 15988 13852 15994 13864
rect 16040 13861 16068 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 16850 13920 16856 13932
rect 16807 13892 16856 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 21358 13920 21364 13932
rect 21223 13892 21364 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15988 13824 16037 13852
rect 15988 13812 15994 13824
rect 16025 13821 16037 13824
rect 16071 13821 16083 13855
rect 16482 13852 16488 13864
rect 16443 13824 16488 13852
rect 16025 13815 16083 13821
rect 16482 13812 16488 13824
rect 16540 13852 16546 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 16540 13824 17785 13852
rect 16540 13812 16546 13824
rect 17773 13821 17785 13824
rect 17819 13852 17831 13855
rect 17862 13852 17868 13864
rect 17819 13824 17868 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 19978 13852 19984 13864
rect 19939 13824 19984 13852
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 24648 13855 24706 13861
rect 24648 13821 24660 13855
rect 24694 13852 24706 13855
rect 25130 13852 25136 13864
rect 24694 13824 25136 13852
rect 24694 13821 24706 13824
rect 24648 13815 24706 13821
rect 25130 13812 25136 13824
rect 25188 13812 25194 13864
rect 14277 13787 14335 13793
rect 14277 13784 14289 13787
rect 14255 13756 14289 13784
rect 14277 13753 14289 13756
rect 14323 13753 14335 13787
rect 18506 13784 18512 13796
rect 18467 13756 18512 13784
rect 14277 13747 14335 13753
rect 14292 13716 14320 13747
rect 18506 13744 18512 13756
rect 18564 13744 18570 13796
rect 18601 13787 18659 13793
rect 18601 13753 18613 13787
rect 18647 13753 18659 13787
rect 21266 13784 21272 13796
rect 21227 13756 21272 13784
rect 18601 13747 18659 13753
rect 18230 13716 18236 13728
rect 12759 13688 14320 13716
rect 18191 13688 18236 13716
rect 12759 13685 12771 13688
rect 12713 13679 12771 13685
rect 18230 13676 18236 13688
rect 18288 13716 18294 13728
rect 18616 13716 18644 13747
rect 21266 13744 21272 13756
rect 21324 13744 21330 13796
rect 21821 13787 21879 13793
rect 21821 13753 21833 13787
rect 21867 13784 21879 13787
rect 22002 13784 22008 13796
rect 21867 13756 22008 13784
rect 21867 13753 21879 13756
rect 21821 13747 21879 13753
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 18288 13688 18644 13716
rect 18288 13676 18294 13688
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19521 13719 19579 13725
rect 19521 13716 19533 13719
rect 19392 13688 19533 13716
rect 19392 13676 19398 13688
rect 19521 13685 19533 13688
rect 19567 13716 19579 13719
rect 21174 13716 21180 13728
rect 19567 13688 21180 13716
rect 19567 13685 19579 13688
rect 19521 13679 19579 13685
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 21726 13676 21732 13728
rect 21784 13716 21790 13728
rect 24719 13719 24777 13725
rect 24719 13716 24731 13719
rect 21784 13688 24731 13716
rect 21784 13676 21790 13688
rect 24719 13685 24731 13688
rect 24765 13685 24777 13719
rect 24719 13679 24777 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 2740 13484 3157 13512
rect 2740 13472 2746 13484
rect 3145 13481 3157 13484
rect 3191 13512 3203 13515
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 3191 13484 3617 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 3786 13512 3792 13524
rect 3747 13484 3792 13512
rect 3605 13475 3663 13481
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 5500 13484 5917 13512
rect 5500 13472 5506 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 6178 13512 6184 13524
rect 6139 13484 6184 13512
rect 5905 13475 5963 13481
rect 1946 13404 1952 13456
rect 2004 13444 2010 13456
rect 2546 13447 2604 13453
rect 2546 13444 2558 13447
rect 2004 13416 2558 13444
rect 2004 13404 2010 13416
rect 2546 13413 2558 13416
rect 2592 13413 2604 13447
rect 2546 13407 2604 13413
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 4065 13447 4123 13453
rect 4065 13444 4077 13447
rect 2832 13416 4077 13444
rect 2832 13404 2838 13416
rect 4065 13413 4077 13416
rect 4111 13413 4123 13447
rect 4065 13407 4123 13413
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 2314 13376 2320 13388
rect 2096 13348 2320 13376
rect 2096 13336 2102 13348
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13376 3663 13379
rect 4157 13379 4215 13385
rect 4157 13376 4169 13379
rect 3651 13348 4169 13376
rect 3651 13345 3663 13348
rect 3605 13339 3663 13345
rect 4157 13345 4169 13348
rect 4203 13345 4215 13379
rect 5920 13376 5948 13475
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 8202 13512 8208 13524
rect 8163 13484 8208 13512
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9030 13512 9036 13524
rect 8404 13484 9036 13512
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 8404 13444 8432 13484
rect 9030 13472 9036 13484
rect 9088 13512 9094 13524
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 9088 13484 9137 13512
rect 9088 13472 9094 13484
rect 9125 13481 9137 13484
rect 9171 13481 9183 13515
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 9125 13475 9183 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 12802 13512 12808 13524
rect 10933 13484 12808 13512
rect 7616 13416 8432 13444
rect 8711 13447 8769 13453
rect 7616 13404 7622 13416
rect 8711 13413 8723 13447
rect 8757 13444 8769 13447
rect 10933 13444 10961 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 14001 13515 14059 13521
rect 14001 13512 14013 13515
rect 13504 13484 14013 13512
rect 13504 13472 13510 13484
rect 14001 13481 14013 13484
rect 14047 13481 14059 13515
rect 14001 13475 14059 13481
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 16577 13515 16635 13521
rect 16577 13512 16589 13515
rect 16540 13484 16589 13512
rect 16540 13472 16546 13484
rect 16577 13481 16589 13484
rect 16623 13481 16635 13515
rect 16577 13475 16635 13481
rect 18049 13515 18107 13521
rect 18049 13481 18061 13515
rect 18095 13512 18107 13515
rect 18230 13512 18236 13524
rect 18095 13484 18236 13512
rect 18095 13481 18107 13484
rect 18049 13475 18107 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18506 13512 18512 13524
rect 18467 13484 18512 13512
rect 18506 13472 18512 13484
rect 18564 13512 18570 13524
rect 19797 13515 19855 13521
rect 18564 13484 19748 13512
rect 18564 13472 18570 13484
rect 11146 13444 11152 13456
rect 8757 13416 10961 13444
rect 11059 13416 11152 13444
rect 8757 13413 8769 13416
rect 8711 13407 8769 13413
rect 11146 13404 11152 13416
rect 11204 13444 11210 13456
rect 11790 13444 11796 13456
rect 11204 13416 11796 13444
rect 11204 13404 11210 13416
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 13170 13444 13176 13456
rect 13131 13416 13176 13444
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 13722 13444 13728 13456
rect 13683 13416 13728 13444
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 17310 13404 17316 13456
rect 17368 13444 17374 13456
rect 17450 13447 17508 13453
rect 17450 13444 17462 13447
rect 17368 13416 17462 13444
rect 17368 13404 17374 13416
rect 17450 13413 17462 13416
rect 17496 13413 17508 13447
rect 19150 13444 19156 13456
rect 19111 13416 19156 13444
rect 17450 13407 17508 13413
rect 19150 13404 19156 13416
rect 19208 13404 19214 13456
rect 19720 13444 19748 13484
rect 19797 13481 19809 13515
rect 19843 13512 19855 13515
rect 21082 13512 21088 13524
rect 19843 13484 21088 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21177 13515 21235 13521
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 21358 13512 21364 13524
rect 21223 13484 21364 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 21542 13444 21548 13456
rect 19720 13416 21548 13444
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 21818 13444 21824 13456
rect 21779 13416 21824 13444
rect 21818 13404 21824 13416
rect 21876 13404 21882 13456
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5920 13348 6101 13376
rect 4157 13339 4215 13345
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6546 13376 6552 13388
rect 6507 13348 6552 13376
rect 6089 13339 6147 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7190 13376 7196 13388
rect 7147 13348 7196 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 7374 13376 7380 13388
rect 7335 13348 7380 13376
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 8624 13379 8682 13385
rect 8624 13345 8636 13379
rect 8670 13376 8682 13379
rect 9490 13376 9496 13388
rect 8670 13348 9496 13376
rect 8670 13345 8682 13348
rect 8624 13339 8682 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 15562 13376 15568 13388
rect 15523 13348 15568 13376
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16025 13379 16083 13385
rect 16025 13376 16037 13379
rect 15896 13348 16037 13376
rect 15896 13336 15902 13348
rect 16025 13345 16037 13348
rect 16071 13376 16083 13379
rect 16114 13376 16120 13388
rect 16071 13348 16120 13376
rect 16071 13345 16083 13348
rect 16025 13339 16083 13345
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 22370 13336 22376 13388
rect 22428 13376 22434 13388
rect 23382 13376 23388 13388
rect 22428 13348 23388 13376
rect 22428 13336 22434 13348
rect 23382 13336 23388 13348
rect 23440 13376 23446 13388
rect 23604 13379 23662 13385
rect 23604 13376 23616 13379
rect 23440 13348 23616 13376
rect 23440 13336 23446 13348
rect 23604 13345 23616 13348
rect 23650 13345 23662 13379
rect 23604 13339 23662 13345
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 3234 13308 3240 13320
rect 2271 13280 3240 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 3234 13268 3240 13280
rect 3292 13308 3298 13320
rect 3694 13308 3700 13320
rect 3292 13280 3700 13308
rect 3292 13268 3298 13280
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11238 13308 11244 13320
rect 11103 13280 11244 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11238 13268 11244 13280
rect 11296 13308 11302 13320
rect 11514 13308 11520 13320
rect 11296 13280 11520 13308
rect 11296 13268 11302 13280
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 13078 13308 13084 13320
rect 13039 13280 13084 13308
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13308 17187 13311
rect 18138 13308 18144 13320
rect 17175 13280 18144 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 18138 13268 18144 13280
rect 18196 13268 18202 13320
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13308 18935 13311
rect 19518 13308 19524 13320
rect 18923 13280 19524 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 21726 13308 21732 13320
rect 21687 13280 21732 13308
rect 21726 13268 21732 13280
rect 21784 13268 21790 13320
rect 22002 13308 22008 13320
rect 21963 13280 22008 13308
rect 22002 13268 22008 13280
rect 22060 13268 22066 13320
rect 1673 13243 1731 13249
rect 1673 13209 1685 13243
rect 1719 13240 1731 13243
rect 1946 13240 1952 13252
rect 1719 13212 1952 13240
rect 1719 13209 1731 13212
rect 1673 13203 1731 13209
rect 1946 13200 1952 13212
rect 2004 13200 2010 13252
rect 9950 13200 9956 13252
rect 10008 13240 10014 13252
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 10008 13212 11621 13240
rect 10008 13200 10014 13212
rect 11609 13209 11621 13212
rect 11655 13240 11667 13243
rect 11698 13240 11704 13252
rect 11655 13212 11704 13240
rect 11655 13209 11667 13212
rect 11609 13203 11667 13209
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 2038 13172 2044 13184
rect 1999 13144 2044 13172
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 5166 13172 5172 13184
rect 5127 13144 5172 13172
rect 5166 13132 5172 13144
rect 5224 13172 5230 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 5224 13144 5457 13172
rect 5224 13132 5230 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 7834 13172 7840 13184
rect 7795 13144 7840 13172
rect 5445 13135 5503 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 10091 13175 10149 13181
rect 10091 13141 10103 13175
rect 10137 13172 10149 13175
rect 11422 13172 11428 13184
rect 10137 13144 11428 13172
rect 10137 13141 10149 13144
rect 10091 13135 10149 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 19426 13132 19432 13184
rect 19484 13172 19490 13184
rect 20073 13175 20131 13181
rect 20073 13172 20085 13175
rect 19484 13144 20085 13172
rect 19484 13132 19490 13144
rect 20073 13141 20085 13144
rect 20119 13141 20131 13175
rect 20073 13135 20131 13141
rect 23707 13175 23765 13181
rect 23707 13141 23719 13175
rect 23753 13172 23765 13175
rect 24210 13172 24216 13184
rect 23753 13144 24216 13172
rect 23753 13141 23765 13144
rect 23707 13135 23765 13141
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3142 12968 3148 12980
rect 3103 12940 3148 12968
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13170 12968 13176 12980
rect 13127 12940 13176 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12968 15626 12980
rect 16390 12968 16396 12980
rect 15620 12940 16396 12968
rect 15620 12928 15626 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 17865 12971 17923 12977
rect 17865 12937 17877 12971
rect 17911 12968 17923 12971
rect 18138 12968 18144 12980
rect 17911 12940 18144 12968
rect 17911 12937 17923 12940
rect 17865 12931 17923 12937
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 21818 12928 21824 12980
rect 21876 12968 21882 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 21876 12940 22293 12968
rect 21876 12928 21882 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 22281 12931 22339 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 4430 12900 4436 12912
rect 4126 12872 4436 12900
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 1762 12832 1768 12844
rect 1719 12804 1768 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2406 12832 2412 12844
rect 2363 12804 2412 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3510 12832 3516 12844
rect 3375 12804 3516 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3510 12792 3516 12804
rect 3568 12832 3574 12844
rect 4126 12832 4154 12872
rect 4430 12860 4436 12872
rect 4488 12900 4494 12912
rect 7285 12903 7343 12909
rect 7285 12900 7297 12903
rect 4488 12872 7297 12900
rect 4488 12860 4494 12872
rect 7285 12869 7297 12872
rect 7331 12869 7343 12903
rect 7285 12863 7343 12869
rect 8849 12903 8907 12909
rect 8849 12869 8861 12903
rect 8895 12900 8907 12903
rect 9677 12903 9735 12909
rect 9677 12900 9689 12903
rect 8895 12872 9689 12900
rect 8895 12869 8907 12872
rect 8849 12863 8907 12869
rect 9677 12869 9689 12872
rect 9723 12900 9735 12903
rect 9723 12872 10640 12900
rect 9723 12869 9735 12872
rect 9677 12863 9735 12869
rect 3568 12804 4154 12832
rect 7300 12832 7328 12863
rect 9309 12835 9367 12841
rect 7300 12804 8340 12832
rect 3568 12792 3574 12804
rect 8312 12776 8340 12804
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 9490 12832 9496 12844
rect 9355 12804 9496 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 10612 12841 10640 12872
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15712 12872 16037 12900
rect 15712 12860 15718 12872
rect 16025 12869 16037 12872
rect 16071 12869 16083 12903
rect 16025 12863 16083 12869
rect 17129 12903 17187 12909
rect 17129 12869 17141 12903
rect 17175 12900 17187 12903
rect 19886 12900 19892 12912
rect 17175 12872 19892 12900
rect 17175 12869 17187 12872
rect 17129 12863 17187 12869
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 13722 12832 13728 12844
rect 13679 12804 13728 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 13722 12792 13728 12804
rect 13780 12832 13786 12844
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 13780 12804 14565 12832
rect 13780 12792 13786 12804
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3418 12764 3424 12776
rect 3200 12736 3424 12764
rect 3200 12724 3206 12736
rect 3418 12724 3424 12736
rect 3476 12764 3482 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3476 12736 3617 12764
rect 3476 12724 3482 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 4246 12764 4252 12776
rect 4159 12736 4252 12764
rect 3605 12727 3663 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 4430 12724 4436 12776
rect 4488 12764 4494 12776
rect 4982 12764 4988 12776
rect 4488 12736 4533 12764
rect 4943 12736 4988 12764
rect 4488 12724 4494 12736
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7156 12736 7481 12764
rect 7156 12724 7162 12736
rect 7469 12733 7481 12736
rect 7515 12733 7527 12767
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 7469 12727 7527 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8849 12767 8907 12773
rect 8352 12736 8445 12764
rect 8352 12724 8358 12736
rect 8849 12733 8861 12767
rect 8895 12764 8907 12767
rect 8938 12764 8944 12776
rect 8895 12736 8944 12764
rect 8895 12733 8907 12736
rect 8849 12727 8907 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12216 12736 12449 12764
rect 12216 12724 12222 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15838 12764 15844 12776
rect 15059 12736 15844 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 2130 12696 2136 12708
rect 1811 12668 2136 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 2130 12656 2136 12668
rect 2188 12656 2194 12708
rect 4264 12696 4292 12724
rect 5166 12696 5172 12708
rect 4264 12668 5172 12696
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 6181 12699 6239 12705
rect 6181 12665 6193 12699
rect 6227 12696 6239 12699
rect 7374 12696 7380 12708
rect 6227 12668 7380 12696
rect 6227 12665 6239 12668
rect 6181 12659 6239 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 10918 12699 10976 12705
rect 10918 12696 10930 12699
rect 10520 12668 10930 12696
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 2004 12600 2605 12628
rect 2004 12588 2010 12600
rect 2593 12597 2605 12600
rect 2639 12597 2651 12631
rect 2593 12591 2651 12597
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3329 12631 3387 12637
rect 3329 12628 3341 12631
rect 3200 12600 3341 12628
rect 3200 12588 3206 12600
rect 3329 12597 3341 12600
rect 3375 12628 3387 12631
rect 3421 12631 3479 12637
rect 3421 12628 3433 12631
rect 3375 12600 3433 12628
rect 3375 12597 3387 12600
rect 3329 12591 3387 12597
rect 3421 12597 3433 12600
rect 3467 12597 3479 12631
rect 3694 12628 3700 12640
rect 3655 12600 3700 12628
rect 3421 12591 3479 12597
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 5258 12588 5264 12640
rect 5316 12628 5322 12640
rect 5721 12631 5779 12637
rect 5721 12628 5733 12631
rect 5316 12600 5733 12628
rect 5316 12588 5322 12600
rect 5721 12597 5733 12600
rect 5767 12597 5779 12631
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 5721 12591 5779 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 9766 12628 9772 12640
rect 8720 12600 9772 12628
rect 8720 12588 8726 12600
rect 9766 12588 9772 12600
rect 9824 12628 9830 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9824 12600 10057 12628
rect 9824 12588 9830 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 10045 12591 10103 12597
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 10520 12637 10548 12668
rect 10918 12665 10930 12668
rect 10964 12665 10976 12699
rect 10918 12659 10976 12665
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 13449 12699 13507 12705
rect 13449 12696 13461 12699
rect 12952 12668 13461 12696
rect 12952 12656 12958 12668
rect 13449 12665 13461 12668
rect 13495 12696 13507 12699
rect 13725 12699 13783 12705
rect 13725 12696 13737 12699
rect 13495 12668 13737 12696
rect 13495 12665 13507 12668
rect 13449 12659 13507 12665
rect 13725 12665 13737 12668
rect 13771 12665 13783 12699
rect 14274 12696 14280 12708
rect 14235 12668 14280 12696
rect 13725 12659 13783 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14366 12656 14372 12708
rect 14424 12696 14430 12708
rect 15105 12699 15163 12705
rect 15105 12696 15117 12699
rect 14424 12668 15117 12696
rect 14424 12656 14430 12668
rect 15105 12665 15117 12668
rect 15151 12665 15163 12699
rect 16040 12696 16068 12863
rect 19886 12860 19892 12872
rect 19944 12860 19950 12912
rect 23799 12903 23857 12909
rect 23799 12900 23811 12903
rect 21376 12872 23811 12900
rect 16206 12832 16212 12844
rect 16119 12804 16212 12832
rect 16206 12792 16212 12804
rect 16264 12832 16270 12844
rect 17586 12832 17592 12844
rect 16264 12804 17592 12832
rect 16264 12792 16270 12804
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 18874 12832 18880 12844
rect 18787 12804 18880 12832
rect 18874 12792 18880 12804
rect 18932 12832 18938 12844
rect 20070 12832 20076 12844
rect 18932 12804 20076 12832
rect 18932 12792 18938 12804
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 21376 12841 21404 12872
rect 23799 12869 23811 12872
rect 23845 12869 23857 12903
rect 23799 12863 23857 12869
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 20855 12804 21373 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 21542 12792 21548 12844
rect 21600 12832 21606 12844
rect 21637 12835 21695 12841
rect 21637 12832 21649 12835
rect 21600 12804 21649 12832
rect 21600 12792 21606 12804
rect 21637 12801 21649 12804
rect 21683 12801 21695 12835
rect 21637 12795 21695 12801
rect 23750 12773 23756 12776
rect 23728 12767 23756 12773
rect 23728 12764 23740 12767
rect 23663 12736 23740 12764
rect 23728 12733 23740 12736
rect 23808 12764 23814 12776
rect 24121 12767 24179 12773
rect 24121 12764 24133 12767
rect 23808 12736 24133 12764
rect 23728 12727 23756 12733
rect 23750 12724 23756 12727
rect 23808 12724 23814 12736
rect 24121 12733 24133 12736
rect 24167 12733 24179 12767
rect 24121 12727 24179 12733
rect 16530 12699 16588 12705
rect 16530 12696 16542 12699
rect 16040 12668 16542 12696
rect 15105 12659 15163 12665
rect 16530 12665 16542 12668
rect 16576 12696 16588 12699
rect 16758 12696 16764 12708
rect 16576 12668 16764 12696
rect 16576 12665 16588 12668
rect 16530 12659 16588 12665
rect 16758 12656 16764 12668
rect 16816 12696 16822 12708
rect 17310 12696 17316 12708
rect 16816 12668 17316 12696
rect 16816 12656 16822 12668
rect 17310 12656 17316 12668
rect 17368 12696 17374 12708
rect 17405 12699 17463 12705
rect 17405 12696 17417 12699
rect 17368 12668 17417 12696
rect 17368 12656 17374 12668
rect 17405 12665 17417 12668
rect 17451 12665 17463 12699
rect 18230 12696 18236 12708
rect 18191 12668 18236 12696
rect 17405 12659 17463 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 18322 12656 18328 12708
rect 18380 12696 18386 12708
rect 18380 12668 18425 12696
rect 18380 12656 18386 12668
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19484 12668 19809 12696
rect 19484 12656 19490 12668
rect 19797 12665 19809 12668
rect 19843 12665 19855 12699
rect 19797 12659 19855 12665
rect 19886 12656 19892 12708
rect 19944 12696 19950 12708
rect 19944 12668 19989 12696
rect 19944 12656 19950 12668
rect 20070 12656 20076 12708
rect 20128 12696 20134 12708
rect 21177 12699 21235 12705
rect 21177 12696 21189 12699
rect 20128 12668 21189 12696
rect 20128 12656 20134 12668
rect 21177 12665 21189 12668
rect 21223 12696 21235 12699
rect 21453 12699 21511 12705
rect 21453 12696 21465 12699
rect 21223 12668 21465 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 21453 12665 21465 12668
rect 21499 12665 21511 12699
rect 21453 12659 21511 12665
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10192 12600 10517 12628
rect 10192 12588 10198 12600
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 12158 12628 12164 12640
rect 12119 12600 12164 12628
rect 10505 12591 10563 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 19150 12628 19156 12640
rect 19111 12600 19156 12628
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 19518 12628 19524 12640
rect 19479 12600 19524 12628
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 3329 12427 3387 12433
rect 3329 12424 3341 12427
rect 2455 12396 3341 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 3329 12393 3341 12396
rect 3375 12424 3387 12427
rect 4246 12424 4252 12436
rect 3375 12396 4252 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 8846 12424 8852 12436
rect 7340 12396 8852 12424
rect 7340 12384 7346 12396
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 9950 12424 9956 12436
rect 9539 12396 9956 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 11514 12424 11520 12436
rect 11475 12396 11520 12424
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 13078 12384 13084 12396
rect 13136 12424 13142 12436
rect 15427 12427 15485 12433
rect 15427 12424 15439 12427
rect 13136 12396 15439 12424
rect 13136 12384 13142 12396
rect 15427 12393 15439 12396
rect 15473 12393 15485 12427
rect 16206 12424 16212 12436
rect 16167 12396 16212 12424
rect 15427 12387 15485 12393
rect 16206 12384 16212 12396
rect 16264 12384 16270 12436
rect 17681 12427 17739 12433
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 18233 12427 18291 12433
rect 18233 12424 18245 12427
rect 17727 12396 18245 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 18233 12393 18245 12396
rect 18279 12424 18291 12427
rect 18322 12424 18328 12436
rect 18279 12396 18328 12424
rect 18279 12393 18291 12396
rect 18233 12387 18291 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 19208 12396 19257 12424
rect 19208 12384 19214 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 19978 12384 19984 12436
rect 20036 12424 20042 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 20036 12396 20085 12424
rect 20036 12384 20042 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 21726 12424 21732 12436
rect 21687 12396 21732 12424
rect 20073 12387 20131 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 3697 12359 3755 12365
rect 3697 12325 3709 12359
rect 3743 12356 3755 12359
rect 3878 12356 3884 12368
rect 3743 12328 3884 12356
rect 3743 12325 3755 12328
rect 3697 12319 3755 12325
rect 3878 12316 3884 12328
rect 3936 12356 3942 12368
rect 4890 12356 4896 12368
rect 3936 12328 4896 12356
rect 3936 12316 3942 12328
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 6457 12359 6515 12365
rect 6457 12325 6469 12359
rect 6503 12356 6515 12359
rect 10318 12356 10324 12368
rect 6503 12328 10324 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 10318 12316 10324 12328
rect 10376 12316 10382 12368
rect 10642 12359 10700 12365
rect 10642 12356 10654 12359
rect 10422 12328 10654 12356
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 1397 12291 1455 12297
rect 1397 12288 1409 12291
rect 1360 12260 1409 12288
rect 1360 12248 1366 12260
rect 1397 12257 1409 12260
rect 1443 12257 1455 12291
rect 1397 12251 1455 12257
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4488 12260 4997 12288
rect 4488 12248 4494 12260
rect 4985 12257 4997 12260
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5224 12260 5457 12288
rect 5224 12248 5230 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5592 12260 5825 12288
rect 5592 12248 5598 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 5813 12251 5871 12257
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 7156 12260 7297 12288
rect 7156 12248 7162 12260
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 7285 12251 7343 12257
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8628 12260 8677 12288
rect 8628 12248 8634 12260
rect 8665 12257 8677 12260
rect 8711 12288 8723 12291
rect 8938 12288 8944 12300
rect 8711 12260 8944 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10422 12288 10450 12328
rect 10642 12325 10654 12328
rect 10688 12325 10700 12359
rect 10642 12319 10700 12325
rect 12805 12359 12863 12365
rect 12805 12325 12817 12359
rect 12851 12356 12863 12359
rect 13814 12356 13820 12368
rect 12851 12328 13820 12356
rect 12851 12325 12863 12328
rect 12805 12319 12863 12325
rect 13814 12316 13820 12328
rect 13872 12356 13878 12368
rect 13872 12328 13917 12356
rect 13872 12316 13878 12328
rect 16850 12316 16856 12368
rect 16908 12356 16914 12368
rect 17082 12359 17140 12365
rect 17082 12356 17094 12359
rect 16908 12328 17094 12356
rect 16908 12316 16914 12328
rect 17082 12325 17094 12328
rect 17128 12325 17140 12359
rect 17082 12319 17140 12325
rect 21818 12316 21824 12368
rect 21876 12356 21882 12368
rect 22097 12359 22155 12365
rect 22097 12356 22109 12359
rect 21876 12328 22109 12356
rect 21876 12316 21882 12328
rect 22097 12325 22109 12328
rect 22143 12325 22155 12359
rect 22097 12319 22155 12325
rect 10192 12260 10450 12288
rect 11241 12291 11299 12297
rect 10192 12248 10198 12260
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 11287 12260 12725 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 12713 12257 12725 12260
rect 12759 12288 12771 12291
rect 12894 12288 12900 12300
rect 12759 12260 12900 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 15286 12288 15292 12300
rect 15344 12297 15350 12300
rect 15344 12291 15382 12297
rect 14884 12260 15292 12288
rect 14884 12248 14890 12260
rect 15286 12248 15292 12260
rect 15370 12257 15382 12291
rect 15344 12251 15382 12257
rect 15344 12248 15350 12251
rect 16298 12248 16304 12300
rect 16356 12288 16362 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16356 12260 16773 12288
rect 16356 12248 16362 12260
rect 16761 12257 16773 12260
rect 16807 12288 16819 12291
rect 16942 12288 16948 12300
rect 16807 12260 16948 12288
rect 16807 12257 16819 12260
rect 16761 12251 16819 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 18230 12248 18236 12300
rect 18288 12288 18294 12300
rect 18509 12291 18567 12297
rect 18509 12288 18521 12291
rect 18288 12260 18521 12288
rect 18288 12248 18294 12260
rect 18509 12257 18521 12260
rect 18555 12288 18567 12291
rect 19334 12288 19340 12300
rect 18555 12260 19340 12288
rect 18555 12257 18567 12260
rect 18509 12251 18567 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 20809 12291 20867 12297
rect 20809 12257 20821 12291
rect 20855 12288 20867 12291
rect 20898 12288 20904 12300
rect 20855 12260 20904 12288
rect 20855 12257 20867 12260
rect 20809 12251 20867 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 24556 12291 24614 12297
rect 24556 12257 24568 12291
rect 24602 12288 24614 12291
rect 24946 12288 24952 12300
rect 24602 12260 24952 12288
rect 24602 12257 24614 12260
rect 24556 12251 24614 12257
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 1544 12192 2053 12220
rect 1544 12180 1550 12192
rect 2041 12189 2053 12192
rect 2087 12220 2099 12223
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 2087 12192 2513 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6696 12192 7205 12220
rect 6696 12180 6702 12192
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 8036 12220 8064 12248
rect 7239 12192 8064 12220
rect 8757 12223 8815 12229
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 8757 12189 8769 12223
rect 8803 12220 8815 12223
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 8803 12192 10333 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 10321 12189 10333 12192
rect 10367 12220 10379 12223
rect 10870 12220 10876 12232
rect 10367 12192 10876 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14366 12220 14372 12232
rect 13771 12192 14372 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 22002 12220 22008 12232
rect 21963 12192 22008 12220
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22649 12223 22707 12229
rect 22649 12189 22661 12223
rect 22695 12220 22707 12223
rect 22738 12220 22744 12232
rect 22695 12192 22744 12220
rect 22695 12189 22707 12192
rect 22649 12183 22707 12189
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 22888 12192 23489 12220
rect 22888 12180 22894 12192
rect 23477 12189 23489 12192
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 14274 12152 14280 12164
rect 14235 12124 14280 12152
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 4522 12084 4528 12096
rect 4483 12056 4528 12084
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12084 4951 12087
rect 4982 12084 4988 12096
rect 4939 12056 4988 12084
rect 4939 12053 4951 12056
rect 4893 12047 4951 12053
rect 4982 12044 4988 12056
rect 5040 12084 5046 12096
rect 5534 12084 5540 12096
rect 5040 12056 5540 12084
rect 5040 12044 5046 12056
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 6730 12084 6736 12096
rect 6691 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 9030 12084 9036 12096
rect 8991 12056 9036 12084
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 9732 12056 9873 12084
rect 9732 12044 9738 12056
rect 9861 12053 9873 12056
rect 9907 12053 9919 12087
rect 13538 12084 13544 12096
rect 13499 12056 13544 12084
rect 9861 12047 9919 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 15838 12084 15844 12096
rect 15799 12056 15844 12084
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 19794 12084 19800 12096
rect 19755 12056 19800 12084
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 20346 12044 20352 12096
rect 20404 12084 20410 12096
rect 21039 12087 21097 12093
rect 21039 12084 21051 12087
rect 20404 12056 21051 12084
rect 20404 12044 20410 12056
rect 21039 12053 21051 12056
rect 21085 12053 21097 12087
rect 21039 12047 21097 12053
rect 24627 12087 24685 12093
rect 24627 12053 24639 12087
rect 24673 12084 24685 12087
rect 24854 12084 24860 12096
rect 24673 12056 24860 12084
rect 24673 12053 24685 12056
rect 24627 12047 24685 12053
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7742 11880 7748 11892
rect 7064 11852 7748 11880
rect 7064 11840 7070 11852
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 8294 11880 8300 11892
rect 7883 11852 8300 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 10870 11880 10876 11892
rect 10831 11852 10876 11880
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12894 11880 12900 11892
rect 12299 11852 12900 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14277 11883 14335 11889
rect 13872 11852 13917 11880
rect 13872 11840 13878 11852
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14366 11880 14372 11892
rect 14323 11852 14372 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 16758 11880 16764 11892
rect 16719 11852 16764 11880
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17129 11883 17187 11889
rect 17129 11880 17141 11883
rect 17000 11852 17141 11880
rect 17000 11840 17006 11852
rect 17129 11849 17141 11852
rect 17175 11849 17187 11883
rect 17129 11843 17187 11849
rect 19794 11840 19800 11892
rect 19852 11880 19858 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 19852 11852 21465 11880
rect 19852 11840 19858 11852
rect 21453 11849 21465 11852
rect 21499 11880 21511 11883
rect 21818 11880 21824 11892
rect 21499 11852 21824 11880
rect 21499 11849 21511 11852
rect 21453 11843 21511 11849
rect 21818 11840 21824 11852
rect 21876 11840 21882 11892
rect 22002 11840 22008 11892
rect 22060 11880 22066 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22060 11852 23029 11880
rect 22060 11840 22066 11852
rect 23017 11849 23029 11852
rect 23063 11849 23075 11883
rect 23017 11843 23075 11849
rect 24673 11883 24731 11889
rect 24673 11849 24685 11883
rect 24719 11880 24731 11883
rect 24762 11880 24768 11892
rect 24719 11852 24768 11880
rect 24719 11849 24731 11852
rect 24673 11843 24731 11849
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 11885 11815 11943 11821
rect 3476 11784 4200 11812
rect 3476 11772 3482 11784
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 3602 11744 3608 11756
rect 3563 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11676 3295 11679
rect 3326 11676 3332 11688
rect 3283 11648 3332 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3326 11636 3332 11648
rect 3384 11676 3390 11688
rect 4172 11676 4200 11784
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 12342 11812 12348 11824
rect 11931 11784 12348 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4341 11747 4399 11753
rect 4341 11744 4353 11747
rect 4304 11716 4353 11744
rect 4304 11704 4310 11716
rect 4341 11713 4353 11716
rect 4387 11744 4399 11747
rect 4522 11744 4528 11756
rect 4387 11716 4528 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4522 11704 4528 11716
rect 4580 11744 4586 11756
rect 5902 11744 5908 11756
rect 4580 11716 5488 11744
rect 5863 11716 5908 11744
rect 4580 11704 4586 11716
rect 5460 11688 5488 11716
rect 5902 11704 5908 11716
rect 5960 11704 5966 11756
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 10042 11744 10048 11756
rect 10003 11716 10048 11744
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 4430 11676 4436 11688
rect 3384 11648 4016 11676
rect 4172 11648 4436 11676
rect 3384 11636 3390 11648
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11577 1639 11611
rect 2130 11608 2136 11620
rect 2091 11580 2136 11608
rect 1581 11571 1639 11577
rect 1596 11540 1624 11571
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 2961 11611 3019 11617
rect 2961 11577 2973 11611
rect 3007 11608 3019 11611
rect 3053 11611 3111 11617
rect 3053 11608 3065 11611
rect 3007 11580 3065 11608
rect 3007 11577 3019 11580
rect 2961 11571 3019 11577
rect 3053 11577 3065 11580
rect 3099 11608 3111 11611
rect 3602 11608 3608 11620
rect 3099 11580 3608 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 3988 11617 4016 11648
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5442 11676 5448 11688
rect 5403 11648 5448 11676
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 8110 11676 8116 11688
rect 8071 11648 8116 11676
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8260 11648 8401 11676
rect 8260 11636 8266 11648
rect 8389 11645 8401 11648
rect 8435 11676 8447 11679
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8435 11648 8953 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 11400 11679 11458 11685
rect 11400 11645 11412 11679
rect 11446 11676 11458 11679
rect 11900 11676 11928 11775
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 16776 11812 16804 11840
rect 17773 11815 17831 11821
rect 17773 11812 17785 11815
rect 16776 11784 17785 11812
rect 17773 11781 17785 11784
rect 17819 11781 17831 11815
rect 17773 11775 17831 11781
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 13538 11744 13544 11756
rect 12943 11716 13544 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 17402 11744 17408 11756
rect 15764 11716 17408 11744
rect 14458 11676 14464 11688
rect 11446 11648 11928 11676
rect 14419 11648 14464 11676
rect 11446 11645 11458 11648
rect 11400 11639 11458 11645
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14516 11648 14933 11676
rect 14516 11636 14522 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 15764 11685 15792 11716
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 15620 11648 15761 11676
rect 15620 11636 15626 11648
rect 15749 11645 15761 11648
rect 15795 11645 15807 11679
rect 15749 11639 15807 11645
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 15896 11648 15945 11676
rect 15896 11636 15902 11648
rect 15933 11645 15945 11648
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 3973 11611 4031 11617
rect 3973 11577 3985 11611
rect 4019 11608 4031 11611
rect 9122 11608 9128 11620
rect 4019 11580 9128 11608
rect 4019 11577 4031 11580
rect 3973 11571 4031 11577
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9582 11608 9588 11620
rect 9543 11580 9588 11608
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 9732 11580 9777 11608
rect 12636 11580 13001 11608
rect 9732 11568 9738 11580
rect 1854 11540 1860 11552
rect 1596 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11540 1918 11552
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 1912 11512 2421 11540
rect 1912 11500 1918 11512
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 2409 11503 2467 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9088 11512 9321 11540
rect 9088 11500 9094 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10192 11512 10517 11540
rect 10192 11500 10198 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11471 11543 11529 11549
rect 11471 11509 11483 11543
rect 11517 11540 11529 11543
rect 11698 11540 11704 11552
rect 11517 11512 11704 11540
rect 11517 11509 11529 11512
rect 11471 11503 11529 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12636 11549 12664 11580
rect 12989 11577 13001 11580
rect 13035 11577 13047 11611
rect 12989 11571 13047 11577
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 13541 11611 13599 11617
rect 13541 11608 13553 11611
rect 13412 11580 13553 11608
rect 13412 11568 13418 11580
rect 13541 11577 13553 11580
rect 13587 11577 13599 11611
rect 16206 11608 16212 11620
rect 16167 11580 16212 11608
rect 13541 11571 13599 11577
rect 16206 11568 16212 11580
rect 16264 11568 16270 11620
rect 17788 11608 17816 11775
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 19613 11815 19671 11821
rect 19613 11812 19625 11815
rect 18932 11784 19625 11812
rect 18932 11772 18938 11784
rect 19613 11781 19625 11784
rect 19659 11781 19671 11815
rect 20898 11812 20904 11824
rect 20859 11784 20904 11812
rect 19613 11775 19671 11781
rect 20898 11772 20904 11784
rect 20956 11772 20962 11824
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11744 19947 11747
rect 20346 11744 20352 11756
rect 19935 11716 20352 11744
rect 19935 11713 19947 11716
rect 19889 11707 19947 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 22094 11744 22100 11756
rect 22007 11716 22100 11744
rect 22094 11704 22100 11716
rect 22152 11744 22158 11756
rect 22830 11744 22836 11756
rect 22152 11716 22836 11744
rect 22152 11704 22158 11716
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 24188 11679 24246 11685
rect 24188 11645 24200 11679
rect 24234 11676 24246 11679
rect 24688 11676 24716 11843
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 24234 11648 24716 11676
rect 24234 11645 24246 11648
rect 24188 11639 24246 11645
rect 18370 11611 18428 11617
rect 18370 11608 18382 11611
rect 17788 11580 18382 11608
rect 18370 11577 18382 11580
rect 18416 11608 18428 11611
rect 19150 11608 19156 11620
rect 18416 11580 19156 11608
rect 18416 11577 18428 11580
rect 18370 11571 18428 11577
rect 19150 11568 19156 11580
rect 19208 11608 19214 11620
rect 19245 11611 19303 11617
rect 19245 11608 19257 11611
rect 19208 11580 19257 11608
rect 19208 11568 19214 11580
rect 19245 11577 19257 11580
rect 19291 11577 19303 11611
rect 19978 11608 19984 11620
rect 19939 11580 19984 11608
rect 19245 11571 19303 11577
rect 19978 11568 19984 11580
rect 20036 11568 20042 11620
rect 20533 11611 20591 11617
rect 20533 11577 20545 11611
rect 20579 11577 20591 11611
rect 20533 11571 20591 11577
rect 12621 11543 12679 11549
rect 12621 11540 12633 11543
rect 12492 11512 12633 11540
rect 12492 11500 12498 11512
rect 12621 11509 12633 11512
rect 12667 11509 12679 11543
rect 12621 11503 12679 11509
rect 14645 11543 14703 11549
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 15838 11540 15844 11552
rect 14691 11512 15844 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 18966 11540 18972 11552
rect 18927 11512 18972 11540
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 20548 11540 20576 11571
rect 22186 11568 22192 11620
rect 22244 11608 22250 11620
rect 22738 11608 22744 11620
rect 22244 11580 22289 11608
rect 22699 11580 22744 11608
rect 22244 11568 22250 11580
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 19576 11512 20576 11540
rect 21913 11543 21971 11549
rect 19576 11500 19582 11512
rect 21913 11509 21925 11543
rect 21959 11540 21971 11543
rect 22204 11540 22232 11568
rect 21959 11512 22232 11540
rect 21959 11509 21971 11512
rect 21913 11503 21971 11509
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 24259 11543 24317 11549
rect 24259 11540 24271 11543
rect 22336 11512 24271 11540
rect 22336 11500 22342 11512
rect 24259 11509 24271 11512
rect 24305 11509 24317 11543
rect 24946 11540 24952 11552
rect 24907 11512 24952 11540
rect 24259 11503 24317 11509
rect 24946 11500 24952 11512
rect 25004 11500 25010 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3234 11336 3240 11348
rect 3191 11308 3240 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11305 4399 11339
rect 4341 11299 4399 11305
rect 1759 11271 1817 11277
rect 1759 11237 1771 11271
rect 1805 11268 1817 11271
rect 1946 11268 1952 11280
rect 1805 11240 1952 11268
rect 1805 11237 1817 11240
rect 1759 11231 1817 11237
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 4356 11268 4384 11299
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 4488 11308 5733 11336
rect 4488 11296 4494 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 5905 11339 5963 11345
rect 5905 11305 5917 11339
rect 5951 11336 5963 11339
rect 6270 11336 6276 11348
rect 5951 11308 6276 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 6270 11296 6276 11308
rect 6328 11296 6334 11348
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 8481 11339 8539 11345
rect 8481 11336 8493 11339
rect 6840 11308 8493 11336
rect 2240 11240 4384 11268
rect 2240 11212 2268 11240
rect 5166 11228 5172 11280
rect 5224 11268 5230 11280
rect 6840 11268 6868 11308
rect 8481 11305 8493 11308
rect 8527 11305 8539 11339
rect 8481 11299 8539 11305
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 8720 11308 9904 11336
rect 8720 11296 8726 11308
rect 5224 11240 6868 11268
rect 5224 11228 5230 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2222 11200 2228 11212
rect 1443 11172 2228 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 4154 11200 4160 11212
rect 2823 11172 4160 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 4154 11160 4160 11172
rect 4212 11200 4218 11212
rect 4522 11200 4528 11212
rect 4212 11172 4305 11200
rect 4483 11172 4528 11200
rect 4212 11160 4218 11172
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4890 11200 4896 11212
rect 4851 11172 4896 11200
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5626 11200 5632 11212
rect 5491 11172 5632 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5721 11203 5779 11209
rect 5721 11169 5733 11203
rect 5767 11200 5779 11203
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 5767 11172 6377 11200
rect 5767 11169 5779 11172
rect 5721 11163 5779 11169
rect 6365 11169 6377 11172
rect 6411 11200 6423 11203
rect 6730 11200 6736 11212
rect 6411 11172 6736 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 6840 11209 6868 11240
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 9766 11268 9772 11280
rect 6972 11240 9772 11268
rect 6972 11228 6978 11240
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 9876 11277 9904 11308
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12069 11339 12127 11345
rect 12069 11336 12081 11339
rect 11756 11308 12081 11336
rect 11756 11296 11762 11308
rect 12069 11305 12081 11308
rect 12115 11336 12127 11339
rect 12115 11308 12388 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12360 11277 12388 11308
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15562 11336 15568 11348
rect 14792 11308 15568 11336
rect 14792 11296 14798 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 22094 11336 22100 11348
rect 22055 11308 22100 11336
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 9861 11271 9919 11277
rect 9861 11237 9873 11271
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11237 12403 11271
rect 12345 11231 12403 11237
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 12492 11240 12537 11268
rect 12492 11228 12498 11240
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 17082 11271 17140 11277
rect 17082 11268 17094 11271
rect 16908 11240 17094 11268
rect 16908 11228 16914 11240
rect 17082 11237 17094 11240
rect 17128 11237 17140 11271
rect 17082 11231 17140 11237
rect 18966 11228 18972 11280
rect 19024 11268 19030 11280
rect 19061 11271 19119 11277
rect 19061 11268 19073 11271
rect 19024 11240 19073 11268
rect 19024 11228 19030 11240
rect 19061 11237 19073 11240
rect 19107 11268 19119 11271
rect 19150 11268 19156 11280
rect 19107 11240 19156 11268
rect 19107 11237 19119 11240
rect 19061 11231 19119 11237
rect 19150 11228 19156 11240
rect 19208 11268 19214 11280
rect 20070 11268 20076 11280
rect 19208 11240 20076 11268
rect 19208 11228 19214 11240
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 21082 11268 21088 11280
rect 21043 11240 21088 11268
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 22186 11228 22192 11280
rect 22244 11268 22250 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22244 11240 22477 11268
rect 22244 11228 22250 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11169 6883 11203
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 6825 11163 6883 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7558 11200 7564 11212
rect 7519 11172 7564 11200
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 11308 11203 11366 11209
rect 11308 11169 11320 11203
rect 11354 11200 11366 11203
rect 11974 11200 11980 11212
rect 11354 11172 11980 11200
rect 11354 11169 11366 11172
rect 11308 11163 11366 11169
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 15657 11203 15715 11209
rect 13872 11172 13917 11200
rect 13872 11160 13878 11172
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 15746 11200 15752 11212
rect 15703 11172 15752 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 21818 11160 21824 11212
rect 21876 11200 21882 11212
rect 22554 11200 22560 11212
rect 21876 11172 22560 11200
rect 21876 11160 21882 11172
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 24854 11200 24860 11212
rect 24627 11172 24860 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 5000 11104 9229 11132
rect 1302 11024 1308 11076
rect 1360 11064 1366 11076
rect 5000 11064 5028 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 10042 11132 10048 11144
rect 10003 11104 10048 11132
rect 9217 11095 9275 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11132 11851 11135
rect 12526 11132 12532 11144
rect 11839 11104 12532 11132
rect 11839 11101 11851 11104
rect 11793 11095 11851 11101
rect 12526 11092 12532 11104
rect 12584 11132 12590 11144
rect 13955 11135 14013 11141
rect 13955 11132 13967 11135
rect 12584 11104 13967 11132
rect 12584 11092 12590 11104
rect 13955 11101 13967 11104
rect 14001 11101 14013 11135
rect 16758 11132 16764 11144
rect 16719 11104 16764 11132
rect 13955 11095 14013 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 18969 11135 19027 11141
rect 18969 11101 18981 11135
rect 19015 11132 19027 11135
rect 19058 11132 19064 11144
rect 19015 11104 19064 11132
rect 19015 11101 19027 11104
rect 18969 11095 19027 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19334 11132 19340 11144
rect 19295 11104 19340 11132
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 20990 11132 20996 11144
rect 20951 11104 20996 11132
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 1360 11036 5028 11064
rect 5629 11067 5687 11073
rect 1360 11024 1366 11036
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 5675 11036 6285 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 6273 11033 6285 11036
rect 6319 11064 6331 11067
rect 7558 11064 7564 11076
rect 6319 11036 7564 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 8849 11067 8907 11073
rect 8849 11064 8861 11067
rect 8036 11036 8861 11064
rect 2038 10956 2044 11008
rect 2096 10996 2102 11008
rect 2222 10996 2228 11008
rect 2096 10968 2228 10996
rect 2096 10956 2102 10968
rect 2222 10956 2228 10968
rect 2280 10996 2286 11008
rect 2317 10999 2375 11005
rect 2317 10996 2329 10999
rect 2280 10968 2329 10996
rect 2280 10956 2286 10968
rect 2317 10965 2329 10968
rect 2363 10965 2375 10999
rect 2317 10959 2375 10965
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 8036 10996 8064 11036
rect 8849 11033 8861 11036
rect 8895 11064 8907 11067
rect 9030 11064 9036 11076
rect 8895 11036 9036 11064
rect 8895 11033 8907 11036
rect 8849 11027 8907 11033
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 12897 11067 12955 11073
rect 12897 11033 12909 11067
rect 12943 11064 12955 11067
rect 13170 11064 13176 11076
rect 12943 11036 13176 11064
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 21542 11064 21548 11076
rect 21503 11036 21548 11064
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 24762 11064 24768 11076
rect 24723 11036 24768 11064
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 7156 10968 8064 10996
rect 7156 10956 7162 10968
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8205 10999 8263 11005
rect 8205 10996 8217 10999
rect 8168 10968 8217 10996
rect 8168 10956 8174 10968
rect 8205 10965 8217 10968
rect 8251 10996 8263 10999
rect 8478 10996 8484 11008
rect 8251 10968 8484 10996
rect 8251 10965 8263 10968
rect 8205 10959 8263 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 10778 10996 10784 11008
rect 9640 10968 10784 10996
rect 9640 10956 9646 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11379 10999 11437 11005
rect 11379 10965 11391 10999
rect 11425 10996 11437 10999
rect 12618 10996 12624 11008
rect 11425 10968 12624 10996
rect 11425 10965 11437 10968
rect 11379 10959 11437 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 12860 10968 13277 10996
rect 12860 10956 12866 10968
rect 13265 10965 13277 10968
rect 13311 10965 13323 10999
rect 13265 10959 13323 10965
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 14240 10968 14289 10996
rect 14240 10956 14246 10968
rect 14277 10965 14289 10968
rect 14323 10965 14335 10999
rect 14277 10959 14335 10965
rect 15887 10999 15945 11005
rect 15887 10965 15899 10999
rect 15933 10996 15945 10999
rect 16482 10996 16488 11008
rect 15933 10968 16488 10996
rect 15933 10965 15945 10968
rect 15887 10959 15945 10965
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 17678 10996 17684 11008
rect 17639 10968 17684 10996
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 18046 10996 18052 11008
rect 18007 10968 18052 10996
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 19886 10996 19892 11008
rect 19847 10968 19892 10996
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3326 10792 3332 10804
rect 3287 10764 3332 10792
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 3476 10764 4169 10792
rect 3476 10752 3482 10764
rect 4157 10761 4169 10764
rect 4203 10792 4215 10795
rect 4522 10792 4528 10804
rect 4203 10764 4528 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 5500 10764 6285 10792
rect 5500 10752 5506 10764
rect 6273 10761 6285 10764
rect 6319 10792 6331 10795
rect 7926 10792 7932 10804
rect 6319 10764 7932 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 9824 10764 10609 10792
rect 9824 10752 9830 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 17770 10752 17776 10804
rect 17828 10792 17834 10804
rect 19886 10792 19892 10804
rect 17828 10764 19892 10792
rect 17828 10752 17834 10764
rect 19886 10752 19892 10764
rect 19944 10792 19950 10804
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 19944 10764 20361 10792
rect 19944 10752 19950 10764
rect 20349 10761 20361 10764
rect 20395 10792 20407 10795
rect 20714 10792 20720 10804
rect 20395 10764 20720 10792
rect 20395 10761 20407 10764
rect 20349 10755 20407 10761
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 21140 10764 21557 10792
rect 21140 10752 21146 10764
rect 21545 10761 21557 10764
rect 21591 10761 21603 10795
rect 22554 10792 22560 10804
rect 22515 10764 22560 10792
rect 21545 10755 21603 10761
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 24673 10795 24731 10801
rect 24673 10761 24685 10795
rect 24719 10792 24731 10795
rect 24854 10792 24860 10804
rect 24719 10764 24860 10792
rect 24719 10761 24731 10764
rect 24673 10755 24731 10761
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 2038 10724 2044 10736
rect 1504 10696 2044 10724
rect 1504 10665 1532 10696
rect 2038 10684 2044 10696
rect 2096 10724 2102 10736
rect 17037 10727 17095 10733
rect 2096 10696 3188 10724
rect 2096 10684 2102 10696
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 1489 10619 1547 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 2222 10520 2228 10532
rect 1627 10492 2228 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 3053 10523 3111 10529
rect 3053 10489 3065 10523
rect 3099 10489 3111 10523
rect 3160 10520 3188 10696
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 19518 10724 19524 10736
rect 17083 10696 19524 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 19518 10684 19524 10696
rect 19576 10724 19582 10736
rect 19613 10727 19671 10733
rect 19613 10724 19625 10727
rect 19576 10696 19625 10724
rect 19576 10684 19582 10696
rect 19613 10693 19625 10696
rect 19659 10693 19671 10727
rect 20070 10724 20076 10736
rect 20031 10696 20076 10724
rect 19613 10687 19671 10693
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 22005 10727 22063 10733
rect 22005 10724 22017 10727
rect 21048 10696 22017 10724
rect 21048 10684 21054 10696
rect 22005 10693 22017 10696
rect 22051 10724 22063 10727
rect 22922 10724 22928 10736
rect 22051 10696 22928 10724
rect 22051 10693 22063 10696
rect 22005 10687 22063 10693
rect 22922 10684 22928 10696
rect 22980 10684 22986 10736
rect 5166 10656 5172 10668
rect 5000 10628 5172 10656
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 4430 10588 4436 10600
rect 3292 10560 3337 10588
rect 4391 10560 4436 10588
rect 3292 10548 3298 10560
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 5000 10597 5028 10628
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 7374 10656 7380 10668
rect 6748 10628 7380 10656
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 4856 10560 4997 10588
rect 4856 10548 4862 10560
rect 4985 10557 4997 10560
rect 5031 10557 5043 10591
rect 4985 10551 5043 10557
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5258 10588 5264 10600
rect 5132 10560 5264 10588
rect 5132 10548 5138 10560
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5408 10560 5825 10588
rect 5408 10548 5414 10560
rect 5813 10557 5825 10560
rect 5859 10588 5871 10591
rect 6270 10588 6276 10600
rect 5859 10560 6276 10588
rect 5859 10557 5871 10560
rect 5813 10551 5871 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10588 6607 10591
rect 6748 10588 6776 10628
rect 7374 10616 7380 10628
rect 7432 10656 7438 10668
rect 8938 10656 8944 10668
rect 7432 10628 8944 10656
rect 7432 10616 7438 10628
rect 7098 10588 7104 10600
rect 6595 10560 6776 10588
rect 7059 10560 7104 10588
rect 6595 10557 6607 10560
rect 6549 10551 6607 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7558 10588 7564 10600
rect 7519 10560 7564 10588
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 7926 10588 7932 10600
rect 7887 10560 7932 10588
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8496 10597 8524 10628
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 12526 10656 12532 10668
rect 12487 10628 12532 10656
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 16482 10656 16488 10668
rect 16443 10628 16488 10656
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 16816 10628 17785 10656
rect 16816 10616 16822 10628
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 17773 10619 17831 10625
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19058 10656 19064 10668
rect 18923 10628 19064 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19058 10616 19064 10628
rect 19116 10656 19122 10668
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 19116 10628 22109 10656
rect 19116 10616 19122 10628
rect 22097 10625 22109 10628
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 9398 10588 9404 10600
rect 8619 10560 9404 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 11216 10591 11274 10597
rect 11216 10588 11228 10591
rect 9548 10560 11228 10588
rect 9548 10548 9554 10560
rect 11216 10557 11228 10560
rect 11262 10588 11274 10591
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 11262 10560 11621 10588
rect 11262 10557 11274 10560
rect 11216 10551 11274 10557
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14182 10588 14188 10600
rect 14047 10560 14188 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 14182 10548 14188 10560
rect 14240 10588 14246 10600
rect 15562 10588 15568 10600
rect 14240 10560 15568 10588
rect 14240 10548 14246 10560
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21542 10588 21548 10600
rect 21315 10560 21548 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 22738 10548 22744 10600
rect 22796 10588 22802 10600
rect 23728 10591 23786 10597
rect 23728 10588 23740 10591
rect 22796 10560 23740 10588
rect 22796 10548 22802 10560
rect 23728 10557 23740 10560
rect 23774 10588 23786 10591
rect 24121 10591 24179 10597
rect 24121 10588 24133 10591
rect 23774 10560 24133 10588
rect 23774 10557 23786 10560
rect 23728 10551 23786 10557
rect 24121 10557 24133 10560
rect 24167 10557 24179 10591
rect 24121 10551 24179 10557
rect 9030 10520 9036 10532
rect 3160 10492 9036 10520
rect 3053 10483 3111 10489
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 2004 10424 2421 10452
rect 2004 10412 2010 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2409 10415 2467 10421
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3068 10452 3096 10483
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10520 9367 10523
rect 9722 10523 9780 10529
rect 9722 10520 9734 10523
rect 9355 10492 9734 10520
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 9722 10489 9734 10492
rect 9768 10520 9780 10523
rect 10134 10520 10140 10532
rect 9768 10492 10140 10520
rect 9768 10489 9780 10492
rect 9722 10483 9780 10489
rect 10134 10480 10140 10492
rect 10192 10520 10198 10532
rect 11054 10520 11060 10532
rect 10192 10492 11060 10520
rect 10192 10480 10198 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10520 12679 10523
rect 12802 10520 12808 10532
rect 12667 10492 12808 10520
rect 12667 10489 12679 10492
rect 12621 10483 12679 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 13170 10520 13176 10532
rect 13131 10492 13176 10520
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 14322 10523 14380 10529
rect 14322 10520 14334 10523
rect 13964 10492 14334 10520
rect 13964 10480 13970 10492
rect 14322 10489 14334 10492
rect 14368 10489 14380 10523
rect 14322 10483 14380 10489
rect 14550 10480 14556 10532
rect 14608 10520 14614 10532
rect 15746 10520 15752 10532
rect 14608 10492 15752 10520
rect 14608 10480 14614 10492
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 16301 10523 16359 10529
rect 16301 10489 16313 10523
rect 16347 10520 16359 10523
rect 16577 10523 16635 10529
rect 16577 10520 16589 10523
rect 16347 10492 16589 10520
rect 16347 10489 16359 10492
rect 16301 10483 16359 10489
rect 16577 10489 16589 10492
rect 16623 10520 16635 10523
rect 17678 10520 17684 10532
rect 16623 10492 17684 10520
rect 16623 10489 16635 10492
rect 16577 10483 16635 10489
rect 17678 10480 17684 10492
rect 17736 10480 17742 10532
rect 19058 10520 19064 10532
rect 19019 10492 19064 10520
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 19150 10480 19156 10532
rect 19208 10520 19214 10532
rect 20622 10520 20628 10532
rect 19208 10492 19253 10520
rect 20583 10492 20628 10520
rect 19208 10480 19214 10492
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 20772 10492 20817 10520
rect 20772 10480 20778 10492
rect 3418 10452 3424 10464
rect 3007 10424 3424 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5224 10424 5641 10452
rect 5224 10412 5230 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 8018 10452 8024 10464
rect 6788 10424 8024 10452
rect 6788 10412 6794 10424
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8720 10424 8861 10452
rect 8720 10412 8726 10424
rect 8849 10421 8861 10424
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9640 10424 10333 10452
rect 9640 10412 9646 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11287 10455 11345 10461
rect 11287 10452 11299 10455
rect 11020 10424 11299 10452
rect 11020 10412 11026 10424
rect 11287 10421 11299 10424
rect 11333 10421 11345 10455
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 11287 10415 11345 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 12400 10424 13461 10452
rect 12400 10412 12406 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13449 10415 13507 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14921 10455 14979 10461
rect 13872 10424 13917 10452
rect 13872 10412 13878 10424
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15654 10452 15660 10464
rect 14967 10424 15660 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 16850 10412 16856 10464
rect 16908 10452 16914 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 16908 10424 17417 10452
rect 16908 10412 16914 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 19168 10452 19196 10480
rect 18555 10424 19196 10452
rect 23799 10455 23857 10461
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 23799 10421 23811 10455
rect 23845 10452 23857 10455
rect 24578 10452 24584 10464
rect 23845 10424 24584 10452
rect 23845 10421 23857 10424
rect 23799 10415 23857 10421
rect 24578 10412 24584 10424
rect 24636 10412 24642 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3510 10248 3516 10260
rect 3471 10220 3516 10248
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 7190 10248 7196 10260
rect 6595 10220 7196 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8018 10248 8024 10260
rect 7979 10220 8024 10248
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 9030 10248 9036 10260
rect 8991 10220 9036 10248
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9398 10248 9404 10260
rect 9359 10220 9404 10248
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 10686 10248 10692 10260
rect 9907 10220 10692 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 14090 10248 14096 10260
rect 10933 10220 13492 10248
rect 14003 10220 14096 10248
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 3050 10180 3056 10192
rect 2915 10152 3056 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 3050 10140 3056 10152
rect 3108 10180 3114 10192
rect 4798 10180 4804 10192
rect 3108 10152 4804 10180
rect 3108 10140 3114 10152
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 5813 10183 5871 10189
rect 5813 10149 5825 10183
rect 5859 10180 5871 10183
rect 8662 10180 8668 10192
rect 5859 10152 8668 10180
rect 5859 10149 5871 10152
rect 5813 10143 5871 10149
rect 8662 10140 8668 10152
rect 8720 10140 8726 10192
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 10933 10180 10961 10220
rect 8803 10152 10961 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 11054 10140 11060 10192
rect 11112 10180 11118 10192
rect 11194 10183 11252 10189
rect 11194 10180 11206 10183
rect 11112 10152 11206 10180
rect 11112 10140 11118 10152
rect 11194 10149 11206 10152
rect 11240 10180 11252 10183
rect 11606 10180 11612 10192
rect 11240 10152 11612 10180
rect 11240 10149 11252 10152
rect 11194 10143 11252 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 12802 10180 12808 10192
rect 11808 10152 12808 10180
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2222 10112 2228 10124
rect 2087 10084 2228 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3142 10112 3148 10124
rect 3007 10084 3148 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3752 10084 4077 10112
rect 3752 10072 3758 10084
rect 4065 10081 4077 10084
rect 4111 10112 4123 10115
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4111 10084 4537 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 5258 10112 5264 10124
rect 5219 10084 5264 10112
rect 4525 10075 4583 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 6641 10115 6699 10121
rect 6641 10081 6653 10115
rect 6687 10112 6699 10115
rect 6822 10112 6828 10124
rect 6687 10084 6828 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6932 10044 6960 10075
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 7064 10084 8217 10112
rect 7064 10072 7070 10084
rect 8205 10081 8217 10084
rect 8251 10112 8263 10115
rect 8294 10112 8300 10124
rect 8251 10084 8300 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 9122 10112 9128 10124
rect 8444 10084 9128 10112
rect 8444 10072 8450 10084
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10134 10112 10140 10124
rect 9723 10084 10140 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11808 10121 11836 10152
rect 12802 10140 12808 10152
rect 12860 10140 12866 10192
rect 13354 10180 13360 10192
rect 13315 10152 13360 10180
rect 13354 10140 13360 10152
rect 13412 10140 13418 10192
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10081 11851 10115
rect 12066 10112 12072 10124
rect 12027 10084 12072 10112
rect 11793 10075 11851 10081
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 7374 10044 7380 10056
rect 6144 10016 6960 10044
rect 7335 10016 7380 10044
rect 6144 10004 6150 10016
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 10870 10044 10876 10056
rect 10831 10016 10876 10044
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 12084 10044 12112 10072
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12084 10016 12725 10044
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 13372 10044 13400 10140
rect 13464 10112 13492 10220
rect 14090 10208 14096 10220
rect 14148 10248 14154 10260
rect 15378 10248 15384 10260
rect 14148 10220 15384 10248
rect 14148 10208 14154 10220
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 20993 10251 21051 10257
rect 20993 10248 21005 10251
rect 16776 10220 21005 10248
rect 15470 10180 15476 10192
rect 15431 10152 15476 10180
rect 15470 10140 15476 10152
rect 15528 10140 15534 10192
rect 15562 10140 15568 10192
rect 15620 10180 15626 10192
rect 16776 10180 16804 10220
rect 20993 10217 21005 10220
rect 21039 10217 21051 10251
rect 20993 10211 21051 10217
rect 23658 10208 23664 10260
rect 23716 10257 23722 10260
rect 23716 10251 23765 10257
rect 23716 10217 23719 10251
rect 23753 10217 23765 10251
rect 23716 10211 23765 10217
rect 23716 10208 23722 10211
rect 15620 10152 16804 10180
rect 15620 10140 15626 10152
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17174 10183 17232 10189
rect 17174 10180 17186 10183
rect 17000 10152 17186 10180
rect 17000 10140 17006 10152
rect 17174 10149 17186 10152
rect 17220 10149 17232 10183
rect 17174 10143 17232 10149
rect 17678 10140 17684 10192
rect 17736 10180 17742 10192
rect 18969 10183 19027 10189
rect 18969 10180 18981 10183
rect 17736 10152 18981 10180
rect 17736 10140 17742 10152
rect 18969 10149 18981 10152
rect 19015 10180 19027 10183
rect 19150 10180 19156 10192
rect 19015 10152 19156 10180
rect 19015 10149 19027 10152
rect 18969 10143 19027 10149
rect 19150 10140 19156 10152
rect 19208 10180 19214 10192
rect 21082 10180 21088 10192
rect 19208 10152 21088 10180
rect 19208 10140 19214 10152
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 13630 10112 13636 10124
rect 13464 10084 13636 10112
rect 13630 10072 13636 10084
rect 13688 10112 13694 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13688 10084 14197 10112
rect 13688 10072 13694 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 16206 10072 16212 10124
rect 16264 10112 16270 10124
rect 16853 10115 16911 10121
rect 16853 10112 16865 10115
rect 16264 10084 16865 10112
rect 16264 10072 16270 10084
rect 16853 10081 16865 10084
rect 16899 10112 16911 10115
rect 17310 10112 17316 10124
rect 16899 10084 17316 10112
rect 16899 10081 16911 10084
rect 16853 10075 16911 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 20898 10112 20904 10124
rect 20859 10084 20904 10112
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21358 10112 21364 10124
rect 21319 10084 21364 10112
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 23566 10112 23572 10124
rect 23527 10084 23572 10112
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 24578 10112 24584 10124
rect 24539 10084 24584 10112
rect 24578 10072 24584 10084
rect 24636 10072 24642 10124
rect 13722 10044 13728 10056
rect 13372 10016 13728 10044
rect 12713 10007 12771 10013
rect 13722 10004 13728 10016
rect 13780 10044 13786 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 13780 10016 15393 10044
rect 13780 10004 13786 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 15381 10007 15439 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 18874 10044 18880 10056
rect 18739 10016 18880 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 19334 10044 19340 10056
rect 19295 10016 19340 10044
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 5074 9976 5080 9988
rect 3896 9948 5080 9976
rect 3896 9920 3924 9948
rect 5074 9936 5080 9948
rect 5132 9976 5138 9988
rect 6365 9979 6423 9985
rect 6365 9976 6377 9979
rect 5132 9948 6377 9976
rect 5132 9936 5138 9948
rect 6365 9945 6377 9948
rect 6411 9976 6423 9979
rect 6549 9979 6607 9985
rect 6549 9976 6561 9979
rect 6411 9948 6561 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 6549 9945 6561 9948
rect 6595 9945 6607 9979
rect 6730 9976 6736 9988
rect 6691 9948 6736 9976
rect 6549 9939 6607 9945
rect 6730 9936 6736 9948
rect 6788 9976 6794 9988
rect 7558 9976 7564 9988
rect 6788 9948 7564 9976
rect 6788 9936 6794 9948
rect 7558 9936 7564 9948
rect 7616 9976 7622 9988
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 7616 9948 7665 9976
rect 7616 9936 7622 9948
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 14369 9979 14427 9985
rect 14369 9976 14381 9979
rect 13596 9948 14381 9976
rect 13596 9936 13602 9948
rect 14369 9945 14381 9948
rect 14415 9945 14427 9979
rect 14369 9939 14427 9945
rect 2406 9908 2412 9920
rect 2367 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4890 9908 4896 9920
rect 4120 9880 4896 9908
rect 4120 9868 4126 9880
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5258 9868 5264 9920
rect 5316 9908 5322 9920
rect 9582 9908 9588 9920
rect 5316 9880 9588 9908
rect 5316 9868 5322 9880
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 12434 9908 12440 9920
rect 12395 9880 12440 9908
rect 12434 9868 12440 9880
rect 12492 9908 12498 9920
rect 12894 9908 12900 9920
rect 12492 9880 12900 9908
rect 12492 9868 12498 9880
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14001 9911 14059 9917
rect 14001 9908 14013 9911
rect 13964 9880 14013 9908
rect 13964 9868 13970 9880
rect 14001 9877 14013 9880
rect 14047 9877 14059 9911
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 14001 9871 14059 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 18138 9908 18144 9920
rect 18099 9880 18144 9908
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 19886 9908 19892 9920
rect 19116 9880 19892 9908
rect 19116 9868 19122 9880
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20622 9908 20628 9920
rect 20583 9880 20628 9908
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 24762 9908 24768 9920
rect 24723 9880 24768 9908
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 14 9664 20 9716
rect 72 9704 78 9716
rect 4338 9704 4344 9716
rect 72 9676 4344 9704
rect 72 9664 78 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6086 9704 6092 9716
rect 5951 9676 6092 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 6641 9707 6699 9713
rect 6641 9673 6653 9707
rect 6687 9704 6699 9707
rect 6822 9704 6828 9716
rect 6687 9676 6828 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8352 9676 8953 9704
rect 8352 9664 8358 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 14734 9704 14740 9716
rect 13786 9676 14740 9704
rect 13786 9674 13814 9676
rect 8941 9667 8999 9673
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 4580 9608 6285 9636
rect 4580 9596 4586 9608
rect 6273 9605 6285 9608
rect 6319 9636 6331 9639
rect 7834 9636 7840 9648
rect 6319 9608 7840 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 7834 9596 7840 9608
rect 7892 9636 7898 9648
rect 7892 9608 8248 9636
rect 7892 9596 7898 9608
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3476 9540 4016 9568
rect 3476 9528 3482 9540
rect 3510 9500 3516 9512
rect 3471 9472 3516 9500
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3988 9509 4016 9540
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6788 9540 7328 9568
rect 6788 9528 6794 9540
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 4304 9472 4353 9500
rect 4304 9460 4310 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 5350 9500 5356 9512
rect 4939 9472 5356 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7098 9500 7104 9512
rect 6871 9472 7104 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 1489 9435 1547 9441
rect 1489 9432 1501 9435
rect 1412 9404 1501 9432
rect 1412 9376 1440 9404
rect 1489 9401 1501 9404
rect 1535 9401 1547 9435
rect 1489 9395 1547 9401
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1670 9432 1676 9444
rect 1627 9404 1676 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2556 9404 3648 9432
rect 2556 9392 2562 9404
rect 1394 9324 1400 9376
rect 1452 9324 1458 9376
rect 1688 9364 1716 9392
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 1688 9336 2421 9364
rect 2409 9333 2421 9336
rect 2455 9333 2467 9367
rect 2409 9327 2467 9333
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3142 9364 3148 9376
rect 3099 9336 3148 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3620 9373 3648 9404
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 6840 9432 6868 9463
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7300 9509 7328 9540
rect 8220 9509 8248 9608
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 13740 9646 13814 9674
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 15105 9707 15163 9713
rect 15105 9673 15117 9707
rect 15151 9704 15163 9707
rect 15470 9704 15476 9716
rect 15151 9676 15476 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15712 9676 15761 9704
rect 15712 9664 15718 9676
rect 15749 9673 15761 9676
rect 15795 9673 15807 9707
rect 15749 9667 15807 9673
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 16945 9707 17003 9713
rect 16945 9704 16957 9707
rect 16908 9676 16957 9704
rect 16908 9664 16914 9676
rect 16945 9673 16957 9676
rect 16991 9673 17003 9707
rect 17310 9704 17316 9716
rect 17271 9676 17316 9704
rect 16945 9667 17003 9673
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 17770 9704 17776 9716
rect 17731 9676 17776 9704
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 19150 9704 19156 9716
rect 19111 9676 19156 9704
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 21315 9707 21373 9713
rect 21315 9704 21327 9707
rect 19944 9676 21327 9704
rect 19944 9664 19950 9676
rect 21315 9673 21327 9676
rect 21361 9673 21373 9707
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 21315 9667 21373 9673
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8444 9608 8585 9636
rect 8444 9596 8450 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 13740 9636 13768 9646
rect 8573 9599 8631 9605
rect 11256 9608 13768 9636
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8386 9500 8392 9512
rect 8251 9472 8392 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 5132 9404 6868 9432
rect 5132 9392 5138 9404
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 7852 9432 7880 9463
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8588 9500 8616 9599
rect 9674 9568 9680 9580
rect 9635 9540 9680 9568
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 11146 9568 11152 9580
rect 11107 9540 11152 9568
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 8588 9472 9321 9500
rect 9309 9469 9321 9472
rect 9355 9500 9367 9503
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9355 9472 9965 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 7926 9432 7932 9444
rect 7616 9404 7932 9432
rect 7616 9392 7622 9404
rect 7926 9392 7932 9404
rect 7984 9432 7990 9444
rect 9122 9432 9128 9444
rect 7984 9404 9128 9432
rect 7984 9392 7990 9404
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 10505 9435 10563 9441
rect 10505 9401 10517 9435
rect 10551 9432 10563 9435
rect 10888 9432 10916 9463
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11256 9500 11284 9608
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 16577 9639 16635 9645
rect 16577 9636 16589 9639
rect 16080 9608 16589 9636
rect 16080 9596 16086 9608
rect 16577 9605 16589 9608
rect 16623 9636 16635 9639
rect 23566 9636 23572 9648
rect 16623 9608 23572 9636
rect 16623 9605 16635 9608
rect 16577 9599 16635 9605
rect 23566 9596 23572 9608
rect 23624 9636 23630 9648
rect 23845 9639 23903 9645
rect 23845 9636 23857 9639
rect 23624 9608 23857 9636
rect 23624 9596 23630 9608
rect 23845 9605 23857 9608
rect 23891 9605 23903 9639
rect 23845 9599 23903 9605
rect 11606 9568 11612 9580
rect 11567 9540 11612 9568
rect 11606 9528 11612 9540
rect 11664 9568 11670 9580
rect 13354 9568 13360 9580
rect 11664 9540 13360 9568
rect 11664 9528 11670 9540
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19334 9568 19340 9580
rect 18831 9540 19340 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19484 9540 20116 9568
rect 19484 9528 19490 9540
rect 11112 9472 11284 9500
rect 12713 9503 12771 9509
rect 11112 9460 11118 9472
rect 12713 9469 12725 9503
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 12253 9435 12311 9441
rect 12253 9432 12265 9435
rect 10551 9404 12265 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 12253 9401 12265 9404
rect 12299 9432 12311 9435
rect 12728 9432 12756 9463
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12952 9472 13001 9500
rect 12952 9460 12958 9472
rect 12989 9469 13001 9472
rect 13035 9500 13047 9503
rect 13262 9500 13268 9512
rect 13035 9472 13268 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 13372 9500 13400 9528
rect 14182 9500 14188 9512
rect 13372 9472 13676 9500
rect 14143 9472 14188 9500
rect 13538 9432 13544 9444
rect 12299 9404 13544 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 13648 9432 13676 9472
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9500 19579 9503
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19567 9472 19625 9500
rect 19567 9469 19579 9472
rect 19521 9463 19579 9469
rect 19613 9469 19625 9472
rect 19659 9500 19671 9503
rect 19978 9500 19984 9512
rect 19659 9472 19984 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20088 9509 20116 9540
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 21244 9503 21302 9509
rect 21244 9469 21256 9503
rect 21290 9500 21302 9503
rect 21290 9472 21680 9500
rect 21290 9469 21302 9472
rect 21244 9463 21302 9469
rect 14001 9435 14059 9441
rect 14001 9432 14013 9435
rect 13648 9404 14013 9432
rect 14001 9401 14013 9404
rect 14047 9432 14059 9435
rect 14506 9435 14564 9441
rect 14506 9432 14518 9435
rect 14047 9404 14518 9432
rect 14047 9401 14059 9404
rect 14001 9395 14059 9401
rect 14506 9401 14518 9404
rect 14552 9401 14564 9435
rect 16022 9432 16028 9444
rect 15983 9404 16028 9432
rect 14506 9395 14564 9401
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9401 16175 9435
rect 18138 9432 18144 9444
rect 18099 9404 18144 9432
rect 16117 9395 16175 9401
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9333 3663 9367
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 3605 9327 3663 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 16132 9364 16160 9395
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 19996 9432 20024 9460
rect 20898 9432 20904 9444
rect 19996 9404 20904 9432
rect 18233 9395 18291 9401
rect 15712 9336 16160 9364
rect 15712 9324 15718 9336
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18248 9364 18276 9395
rect 20898 9392 20904 9404
rect 20956 9392 20962 9444
rect 21652 9376 21680 9472
rect 17828 9336 18276 9364
rect 17828 9324 17834 9336
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 19705 9367 19763 9373
rect 19705 9364 19717 9367
rect 19576 9336 19717 9364
rect 19576 9324 19582 9336
rect 19705 9333 19717 9336
rect 19751 9333 19763 9367
rect 21634 9364 21640 9376
rect 21595 9336 21640 9364
rect 19705 9327 19763 9333
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2685 9163 2743 9169
rect 2685 9129 2697 9163
rect 2731 9160 2743 9163
rect 3510 9160 3516 9172
rect 2731 9132 3516 9160
rect 2731 9129 2743 9132
rect 2685 9123 2743 9129
rect 3510 9120 3516 9132
rect 3568 9160 3574 9172
rect 4154 9160 4160 9172
rect 3568 9132 4160 9160
rect 3568 9120 3574 9132
rect 4154 9120 4160 9132
rect 4212 9160 4218 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4212 9132 4629 9160
rect 4212 9120 4218 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 4617 9123 4675 9129
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 4755 9132 6469 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 6457 9129 6469 9132
rect 6503 9160 6515 9163
rect 6730 9160 6736 9172
rect 6503 9132 6736 9160
rect 6503 9129 6515 9132
rect 6457 9123 6515 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7558 9160 7564 9172
rect 7331 9132 7564 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 9122 9160 9128 9172
rect 9083 9132 9128 9160
rect 9122 9120 9128 9132
rect 9180 9120 9186 9172
rect 9858 9160 9864 9172
rect 9819 9132 9864 9160
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 10928 9132 11069 9160
rect 10928 9120 10934 9132
rect 11057 9129 11069 9132
rect 11103 9160 11115 9163
rect 12526 9160 12532 9172
rect 11103 9132 12532 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 16022 9160 16028 9172
rect 13228 9132 16028 9160
rect 13228 9120 13234 9132
rect 16022 9120 16028 9132
rect 16080 9160 16086 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 16080 9132 16313 9160
rect 16080 9120 16086 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 21039 9163 21097 9169
rect 21039 9160 21051 9163
rect 18196 9132 21051 9160
rect 18196 9120 18202 9132
rect 21039 9129 21051 9132
rect 21085 9129 21097 9163
rect 21358 9160 21364 9172
rect 21319 9132 21364 9160
rect 21039 9123 21097 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 1759 9095 1817 9101
rect 1759 9061 1771 9095
rect 1805 9092 1817 9095
rect 1946 9092 1952 9104
rect 1805 9064 1952 9092
rect 1805 9061 1817 9064
rect 1759 9055 1817 9061
rect 1946 9052 1952 9064
rect 2004 9092 2010 9104
rect 2498 9092 2504 9104
rect 2004 9064 2504 9092
rect 2004 9052 2010 9064
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 3234 9052 3240 9104
rect 3292 9092 3298 9104
rect 5534 9092 5540 9104
rect 3292 9064 5540 9092
rect 3292 9052 3298 9064
rect 5534 9052 5540 9064
rect 5592 9092 5598 9104
rect 6748 9092 6776 9120
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 5592 9064 5672 9092
rect 6748 9064 7665 9092
rect 5592 9052 5598 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2406 9024 2412 9036
rect 1443 8996 2412 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 4338 9024 4344 9036
rect 4299 8996 4344 9024
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 9024 4675 9027
rect 5074 9024 5080 9036
rect 4663 8996 5080 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 5132 8996 5181 9024
rect 5132 8984 5138 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5350 9024 5356 9036
rect 5311 8996 5356 9024
rect 5169 8987 5227 8993
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5644 9033 5672 9064
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 11511 9095 11569 9101
rect 11511 9061 11523 9095
rect 11557 9092 11569 9095
rect 11606 9092 11612 9104
rect 11557 9064 11612 9092
rect 11557 9061 11569 9064
rect 11511 9055 11569 9061
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 12860 9064 13093 9092
rect 12860 9052 12866 9064
rect 13081 9061 13093 9064
rect 13127 9092 13139 9095
rect 13446 9092 13452 9104
rect 13127 9064 13452 9092
rect 13127 9061 13139 9064
rect 13081 9055 13139 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13906 9052 13912 9104
rect 13964 9092 13970 9104
rect 14642 9092 14648 9104
rect 13964 9064 14648 9092
rect 13964 9052 13970 9064
rect 14642 9052 14648 9064
rect 14700 9092 14706 9104
rect 15013 9095 15071 9101
rect 15013 9092 15025 9095
rect 14700 9064 15025 9092
rect 14700 9052 14706 9064
rect 15013 9061 15025 9064
rect 15059 9061 15071 9095
rect 15470 9092 15476 9104
rect 15431 9064 15476 9092
rect 15013 9055 15071 9061
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 17589 9095 17647 9101
rect 17589 9061 17601 9095
rect 17635 9092 17647 9095
rect 18046 9092 18052 9104
rect 17635 9064 18052 9092
rect 17635 9061 17647 9064
rect 17589 9055 17647 9061
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 18288 9064 18920 9092
rect 18288 9052 18294 9064
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 8202 9024 8208 9036
rect 8163 8996 8208 9024
rect 5629 8987 5687 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 11146 9024 11152 9036
rect 11107 8996 11152 9024
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 9024 12127 9027
rect 12342 9024 12348 9036
rect 12115 8996 12348 9024
rect 12115 8993 12127 8996
rect 12069 8987 12127 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13688 8996 14197 9024
rect 13688 8984 13694 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16114 9024 16120 9036
rect 16071 8996 16120 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 17126 9024 17132 9036
rect 17087 8996 17132 9024
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 18598 9024 18604 9036
rect 17460 8996 18604 9024
rect 17460 8984 17466 8996
rect 18598 8984 18604 8996
rect 18656 8984 18662 9036
rect 18892 9033 18920 9064
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 20162 9024 20168 9036
rect 18923 8996 20168 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 20530 8984 20536 9036
rect 20588 9024 20594 9036
rect 20936 9027 20994 9033
rect 20936 9024 20948 9027
rect 20588 8996 20948 9024
rect 20588 8984 20594 8996
rect 20936 8993 20948 8996
rect 20982 8993 20994 9027
rect 20936 8987 20994 8993
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 1636 8928 4721 8956
rect 1636 8916 1642 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 4709 8919 4767 8925
rect 5000 8928 5825 8956
rect 1946 8848 1952 8900
rect 2004 8888 2010 8900
rect 5000 8888 5028 8928
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 5813 8919 5871 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8956 10747 8959
rect 11054 8956 11060 8968
rect 10735 8928 11060 8956
rect 10735 8925 10747 8928
rect 10689 8919 10747 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12618 8916 12624 8968
rect 12676 8956 12682 8968
rect 12986 8956 12992 8968
rect 12676 8928 12992 8956
rect 12676 8916 12682 8928
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13906 8956 13912 8968
rect 13780 8928 13912 8956
rect 13780 8916 13786 8928
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 14016 8928 15393 8956
rect 5442 8888 5448 8900
rect 2004 8860 5028 8888
rect 5403 8860 5448 8888
rect 2004 8848 2010 8860
rect 5442 8848 5448 8860
rect 5500 8848 5506 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9858 8888 9864 8900
rect 8536 8860 9864 8888
rect 8536 8848 8542 8860
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 13280 8888 13308 8916
rect 14016 8888 14044 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 18969 8959 19027 8965
rect 18969 8956 18981 8959
rect 16540 8928 18981 8956
rect 16540 8916 16546 8928
rect 18969 8925 18981 8928
rect 19015 8925 19027 8959
rect 18969 8919 19027 8925
rect 19518 8888 19524 8900
rect 13280 8860 14044 8888
rect 16224 8860 19524 8888
rect 1854 8780 1860 8832
rect 1912 8820 1918 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 1912 8792 2329 8820
rect 1912 8780 1918 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2958 8820 2964 8832
rect 2919 8792 2964 8820
rect 2317 8783 2375 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 4062 8820 4068 8832
rect 3651 8792 4068 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 4062 8780 4068 8792
rect 4120 8820 4126 8832
rect 4246 8820 4252 8832
rect 4120 8792 4252 8820
rect 4120 8780 4126 8792
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 6822 8820 6828 8832
rect 6783 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 10134 8820 10140 8832
rect 10095 8792 10140 8820
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 12526 8820 12532 8832
rect 12487 8792 12532 8820
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 14240 8792 14657 8820
rect 14240 8780 14246 8792
rect 14645 8789 14657 8792
rect 14691 8820 14703 8823
rect 16224 8820 16252 8860
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 18138 8820 18144 8832
rect 14691 8792 16252 8820
rect 18099 8792 18144 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19392 8792 19625 8820
rect 19392 8780 19398 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19613 8783 19671 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2774 8616 2780 8628
rect 2372 8588 2780 8616
rect 2372 8576 2378 8588
rect 2774 8576 2780 8588
rect 2832 8616 2838 8628
rect 4338 8616 4344 8628
rect 2832 8588 3096 8616
rect 4299 8588 4344 8616
rect 2832 8576 2838 8588
rect 2038 8548 2044 8560
rect 1999 8520 2044 8548
rect 2038 8508 2044 8520
rect 2096 8508 2102 8560
rect 3068 8557 3096 8588
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 5534 8616 5540 8628
rect 5495 8588 5540 8616
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 7558 8616 7564 8628
rect 6043 8588 7564 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 3053 8551 3111 8557
rect 3053 8517 3065 8551
rect 3099 8548 3111 8551
rect 4154 8548 4160 8560
rect 3099 8520 4160 8548
rect 3099 8517 3111 8520
rect 3053 8511 3111 8517
rect 4154 8508 4160 8520
rect 4212 8508 4218 8560
rect 5350 8508 5356 8560
rect 5408 8548 5414 8560
rect 6012 8548 6040 8579
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11664 8588 11805 8616
rect 11664 8576 11670 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 11793 8579 11851 8585
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 14921 8619 14979 8625
rect 14921 8585 14933 8619
rect 14967 8616 14979 8619
rect 15289 8619 15347 8625
rect 15289 8616 15301 8619
rect 14967 8588 15301 8616
rect 14967 8585 14979 8588
rect 14921 8579 14979 8585
rect 15289 8585 15301 8588
rect 15335 8616 15347 8619
rect 15470 8616 15476 8628
rect 15335 8588 15476 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 17862 8616 17868 8628
rect 17775 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8616 17926 8628
rect 18230 8616 18236 8628
rect 17920 8588 18236 8616
rect 17920 8576 17926 8588
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18656 8588 19073 8616
rect 18656 8576 18662 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 24762 8616 24768 8628
rect 24723 8588 24768 8616
rect 19061 8579 19119 8585
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 5408 8520 6040 8548
rect 5408 8508 5414 8520
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 9490 8548 9496 8560
rect 6144 8520 9496 8548
rect 6144 8508 6150 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 16942 8548 16948 8560
rect 13596 8520 16948 8548
rect 13596 8508 13602 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 18690 8548 18696 8560
rect 17092 8520 18696 8548
rect 17092 8508 17098 8520
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 3694 8480 3700 8492
rect 3655 8452 3700 8480
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 10134 8480 10140 8492
rect 9171 8452 10140 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10367 8452 10885 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 10873 8449 10885 8452
rect 10919 8480 10931 8483
rect 10962 8480 10968 8492
rect 10919 8452 10968 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 13262 8480 13268 8492
rect 11563 8452 13268 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13817 8483 13875 8489
rect 13817 8480 13829 8483
rect 13412 8452 13829 8480
rect 13412 8440 13418 8452
rect 13817 8449 13829 8452
rect 13863 8480 13875 8483
rect 16485 8483 16543 8489
rect 13863 8452 14365 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 2958 8412 2964 8424
rect 2464 8384 2964 8412
rect 2464 8372 2470 8384
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 4295 8384 4537 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 1854 8344 1860 8356
rect 1627 8316 1860 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 2866 8344 2872 8356
rect 2547 8316 2872 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 2866 8304 2872 8316
rect 2924 8344 2930 8356
rect 3252 8344 3280 8375
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4798 8412 4804 8424
rect 4672 8384 4717 8412
rect 4759 8384 4804 8412
rect 4672 8372 4678 8384
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 6822 8412 6828 8424
rect 6783 8384 6828 8412
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7101 8415 7159 8421
rect 6972 8384 7017 8412
rect 6972 8372 6978 8384
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 8386 8412 8392 8424
rect 8347 8384 8392 8412
rect 7101 8375 7159 8381
rect 4816 8344 4844 8372
rect 2924 8316 4844 8344
rect 2924 8304 2930 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 3016 8248 3985 8276
rect 3016 8236 3022 8248
rect 3973 8245 3985 8248
rect 4019 8276 4031 8279
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 4019 8248 4261 8276
rect 4019 8245 4031 8248
rect 3973 8239 4031 8245
rect 4249 8245 4261 8248
rect 4295 8245 4307 8279
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4249 8239 4307 8245
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 6546 8276 6552 8288
rect 6507 8248 6552 8276
rect 6546 8236 6552 8248
rect 6604 8276 6610 8288
rect 7116 8276 7144 8375
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8481 8415 8539 8421
rect 8481 8381 8493 8415
rect 8527 8381 8539 8415
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8481 8375 8539 8381
rect 7282 8276 7288 8288
rect 6604 8248 7144 8276
rect 7243 8248 7288 8276
rect 6604 8236 6610 8248
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 7929 8279 7987 8285
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 8202 8276 8208 8288
rect 7975 8248 8208 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 8202 8236 8208 8248
rect 8260 8276 8266 8288
rect 8496 8276 8524 8375
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12713 8415 12771 8421
rect 12713 8412 12725 8415
rect 12299 8384 12725 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12713 8381 12725 8384
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13446 8412 13452 8424
rect 13035 8384 13452 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 10689 8347 10747 8353
rect 10689 8313 10701 8347
rect 10735 8344 10747 8347
rect 10965 8347 11023 8353
rect 10965 8344 10977 8347
rect 10735 8316 10977 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 10965 8313 10977 8316
rect 11011 8344 11023 8347
rect 12342 8344 12348 8356
rect 11011 8316 12348 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 12342 8304 12348 8316
rect 12400 8304 12406 8356
rect 12728 8344 12756 8375
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14182 8412 14188 8424
rect 14047 8384 14188 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 13538 8344 13544 8356
rect 12728 8316 13544 8344
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 14337 8353 14365 8452
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16758 8480 16764 8492
rect 16531 8452 16764 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 18138 8480 18144 8492
rect 18051 8452 18144 8480
rect 18138 8440 18144 8452
rect 18196 8480 18202 8492
rect 21315 8483 21373 8489
rect 21315 8480 21327 8483
rect 18196 8452 21327 8480
rect 18196 8440 18202 8452
rect 21315 8449 21327 8452
rect 21361 8449 21373 8483
rect 21315 8443 21373 8449
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 15896 8384 16313 8412
rect 15896 8372 15902 8384
rect 16301 8381 16313 8384
rect 16347 8412 16359 8415
rect 17310 8412 17316 8424
rect 16347 8384 17316 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 19613 8415 19671 8421
rect 19613 8381 19625 8415
rect 19659 8381 19671 8415
rect 20070 8412 20076 8424
rect 20031 8384 20076 8412
rect 19613 8375 19671 8381
rect 14322 8347 14380 8353
rect 14322 8313 14334 8347
rect 14368 8313 14380 8347
rect 14322 8307 14380 8313
rect 15657 8347 15715 8353
rect 15657 8313 15669 8347
rect 15703 8344 15715 8347
rect 17402 8344 17408 8356
rect 15703 8316 17408 8344
rect 15703 8313 15715 8316
rect 15657 8307 15715 8313
rect 9766 8276 9772 8288
rect 8260 8248 8524 8276
rect 9727 8248 9772 8276
rect 8260 8236 8266 8248
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 12526 8276 12532 8288
rect 12487 8248 12532 8276
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 14090 8236 14096 8288
rect 14148 8276 14154 8288
rect 15672 8276 15700 8307
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 18230 8344 18236 8356
rect 18191 8316 18236 8344
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19426 8344 19432 8356
rect 19387 8316 19432 8344
rect 19426 8304 19432 8316
rect 19484 8344 19490 8356
rect 19628 8344 19656 8375
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 21212 8415 21270 8421
rect 21212 8412 21224 8415
rect 20312 8384 21224 8412
rect 20312 8372 20318 8384
rect 21212 8381 21224 8384
rect 21258 8412 21270 8415
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 21258 8384 21649 8412
rect 21258 8381 21270 8384
rect 21212 8375 21270 8381
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21637 8375 21695 8381
rect 24210 8372 24216 8424
rect 24268 8412 24274 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 24268 8384 24593 8412
rect 24268 8372 24274 8384
rect 24581 8381 24593 8384
rect 24627 8412 24639 8415
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24627 8384 25145 8412
rect 24627 8381 24639 8384
rect 24581 8375 24639 8381
rect 25133 8381 25145 8384
rect 25179 8381 25191 8415
rect 25133 8375 25191 8381
rect 19484 8316 19656 8344
rect 19484 8304 19490 8316
rect 14148 8248 15700 8276
rect 16945 8279 17003 8285
rect 14148 8236 14154 8248
rect 16945 8245 16957 8279
rect 16991 8276 17003 8279
rect 17218 8276 17224 8288
rect 16991 8248 17224 8276
rect 16991 8245 17003 8248
rect 16945 8239 17003 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 19334 8276 19340 8288
rect 18196 8248 19340 8276
rect 18196 8236 18202 8248
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 19705 8279 19763 8285
rect 19705 8276 19717 8279
rect 19576 8248 19717 8276
rect 19576 8236 19582 8248
rect 19705 8245 19717 8248
rect 19751 8245 19763 8279
rect 19705 8239 19763 8245
rect 20530 8236 20536 8288
rect 20588 8276 20594 8288
rect 20901 8279 20959 8285
rect 20901 8276 20913 8279
rect 20588 8248 20913 8276
rect 20588 8236 20594 8248
rect 20901 8245 20913 8248
rect 20947 8245 20959 8279
rect 20901 8239 20959 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 2866 8072 2872 8084
rect 2827 8044 2872 8072
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4672 8044 5089 8072
rect 4672 8032 4678 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 5077 8035 5135 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9030 8072 9036 8084
rect 8628 8044 9036 8072
rect 8628 8032 8634 8044
rect 9030 8032 9036 8044
rect 9088 8072 9094 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 9088 8044 9137 8072
rect 9088 8032 9094 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 2317 8007 2375 8013
rect 2317 8004 2329 8007
rect 1412 7976 2329 8004
rect 1412 7945 1440 7976
rect 2317 7973 2329 7976
rect 2363 8004 2375 8007
rect 5460 8004 5488 8032
rect 2363 7976 5488 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 9140 8004 9168 8035
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9824 8044 10149 8072
rect 9824 8032 9830 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 11146 8072 11152 8084
rect 11107 8044 11152 8072
rect 10137 8035 10195 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 11701 8075 11759 8081
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 12526 8072 12532 8084
rect 11747 8044 12532 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 6604 7976 7604 8004
rect 9140 7976 9812 8004
rect 6604 7964 6610 7976
rect 7576 7948 7604 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 1397 7899 1455 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 3384 7908 3801 7936
rect 3384 7896 3390 7908
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 4154 7936 4160 7948
rect 4115 7908 4160 7936
rect 3789 7899 3847 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 5534 7936 5540 7948
rect 4396 7908 5540 7936
rect 4396 7896 4402 7908
rect 5534 7896 5540 7908
rect 5592 7936 5598 7948
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 5592 7908 5825 7936
rect 5592 7896 5598 7908
rect 5813 7905 5825 7908
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7248 7908 7297 7936
rect 7248 7896 7254 7908
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7558 7936 7564 7948
rect 7471 7908 7564 7936
rect 7285 7899 7343 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 8444 7908 8493 7936
rect 8444 7896 8450 7908
rect 8481 7905 8493 7908
rect 8527 7936 8539 7939
rect 9674 7936 9680 7948
rect 8527 7908 9680 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9784 7945 9812 7976
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7905 9827 7939
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9769 7899 9827 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 11808 7945 11836 8044
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12986 8072 12992 8084
rect 12947 8044 12992 8072
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14240 8044 14657 8072
rect 14240 8032 14246 8044
rect 14645 8041 14657 8044
rect 14691 8072 14703 8075
rect 14691 8044 18644 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 12155 8007 12213 8013
rect 12155 7973 12167 8007
rect 12201 7973 12213 8007
rect 13725 8007 13783 8013
rect 13725 8004 13737 8007
rect 12155 7967 12213 7973
rect 12728 7976 13737 8004
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3436 7840 4077 7868
rect 3436 7744 3464 7840
rect 4065 7837 4077 7840
rect 4111 7868 4123 7871
rect 4614 7868 4620 7880
rect 4111 7840 4620 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6822 7868 6828 7880
rect 6503 7840 6828 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 7024 7840 7757 7868
rect 5994 7760 6000 7812
rect 6052 7800 6058 7812
rect 7024 7800 7052 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12176 7868 12204 7967
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12728 7945 12756 7976
rect 13725 7973 13737 7976
rect 13771 8004 13783 8007
rect 14090 8004 14096 8016
rect 13771 7976 14096 8004
rect 13771 7973 13783 7976
rect 13725 7967 13783 7973
rect 14090 7964 14096 7976
rect 14148 7964 14154 8016
rect 15838 8004 15844 8016
rect 15799 7976 15844 8004
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 16298 7964 16304 8016
rect 16356 8004 16362 8016
rect 16806 8007 16864 8013
rect 16806 8004 16818 8007
rect 16356 7976 16818 8004
rect 16356 7964 16362 7976
rect 16806 7973 16818 7976
rect 16852 7973 16864 8007
rect 16806 7967 16864 7973
rect 18322 7964 18328 8016
rect 18380 8004 18386 8016
rect 18417 8007 18475 8013
rect 18417 8004 18429 8007
rect 18380 7976 18429 8004
rect 18380 7964 18386 7976
rect 18417 7973 18429 7976
rect 18463 7973 18475 8007
rect 18616 8004 18644 8044
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 19935 8075 19993 8081
rect 19935 8072 19947 8075
rect 18932 8044 19947 8072
rect 18932 8032 18938 8044
rect 19935 8041 19947 8044
rect 19981 8041 19993 8075
rect 19935 8035 19993 8041
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 21085 8075 21143 8081
rect 21085 8072 21097 8075
rect 20220 8044 21097 8072
rect 20220 8032 20226 8044
rect 21085 8041 21097 8044
rect 21131 8041 21143 8075
rect 21085 8035 21143 8041
rect 19518 8004 19524 8016
rect 18616 7976 19524 8004
rect 18417 7967 18475 7973
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12676 7908 12725 7936
rect 12676 7896 12682 7908
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 12713 7899 12771 7905
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 16482 7936 16488 7948
rect 16443 7908 16488 7936
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 19864 7939 19922 7945
rect 19864 7905 19876 7939
rect 19910 7936 19922 7939
rect 20162 7936 20168 7948
rect 19910 7908 20168 7936
rect 19910 7905 19922 7908
rect 19864 7899 19922 7905
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 20898 7936 20904 7948
rect 20859 7908 20904 7936
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 13630 7868 13636 7880
rect 11664 7840 12204 7868
rect 13591 7840 13636 7868
rect 11664 7828 11670 7840
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13786 7840 14289 7868
rect 6052 7772 7052 7800
rect 7377 7803 7435 7809
rect 6052 7760 6058 7772
rect 7377 7769 7389 7803
rect 7423 7800 7435 7803
rect 8202 7800 8208 7812
rect 7423 7772 8208 7800
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2038 7732 2044 7744
rect 1995 7704 2044 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2038 7692 2044 7704
rect 2096 7732 2102 7744
rect 2498 7732 2504 7744
rect 2096 7704 2504 7732
rect 2096 7692 2102 7704
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 6914 7732 6920 7744
rect 6827 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7732 6978 7744
rect 7392 7732 7420 7763
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 13786 7800 13814 7840
rect 14277 7837 14289 7840
rect 14323 7868 14335 7871
rect 16117 7871 16175 7877
rect 16117 7868 16129 7871
rect 14323 7840 16129 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 16117 7837 16129 7840
rect 16163 7837 16175 7871
rect 18138 7868 18144 7880
rect 16117 7831 16175 7837
rect 16868 7840 18144 7868
rect 15930 7800 15936 7812
rect 13320 7772 13814 7800
rect 15396 7772 15936 7800
rect 13320 7760 13326 7772
rect 6972 7704 7420 7732
rect 6972 7692 6978 7704
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 8720 7704 8769 7732
rect 8720 7692 8726 7704
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 8757 7695 8815 7701
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 11330 7732 11336 7744
rect 10919 7704 11336 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 15396 7732 15424 7772
rect 15930 7760 15936 7772
rect 15988 7800 15994 7812
rect 16868 7800 16896 7840
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 18322 7868 18328 7880
rect 18283 7840 18328 7868
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7868 19027 7871
rect 19518 7868 19524 7880
rect 19015 7840 19524 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 19518 7828 19524 7840
rect 19576 7828 19582 7880
rect 15988 7772 16896 7800
rect 15988 7760 15994 7772
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 17000 7772 19625 7800
rect 17000 7760 17006 7772
rect 19613 7769 19625 7772
rect 19659 7800 19671 7803
rect 20070 7800 20076 7812
rect 19659 7772 20076 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 13504 7704 15424 7732
rect 13504 7692 13510 7704
rect 15470 7692 15476 7744
rect 15528 7732 15534 7744
rect 17405 7735 17463 7741
rect 15528 7704 15573 7732
rect 15528 7692 15534 7704
rect 17405 7701 17417 7735
rect 17451 7732 17463 7735
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 17451 7704 18153 7732
rect 17451 7701 17463 7704
rect 17405 7695 17463 7701
rect 18141 7701 18153 7704
rect 18187 7732 18199 7735
rect 18230 7732 18236 7744
rect 18187 7704 18236 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7528 1676 7540
rect 1631 7500 1676 7528
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5442 7528 5448 7540
rect 5307 7500 5448 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5592 7500 5825 7528
rect 5592 7488 5598 7500
rect 5813 7497 5825 7500
rect 5859 7528 5871 7531
rect 7190 7528 7196 7540
rect 5859 7500 7196 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 7616 7500 8769 7528
rect 7616 7488 7622 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 8757 7491 8815 7497
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3418 7460 3424 7472
rect 3099 7432 3424 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2314 7392 2320 7404
rect 1912 7364 2320 7392
rect 1912 7352 1918 7364
rect 2056 7333 2084 7364
rect 2314 7352 2320 7364
rect 2372 7392 2378 7404
rect 3326 7392 3332 7404
rect 2372 7364 3332 7392
rect 2372 7352 2378 7364
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 8772 7392 8800 7491
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 9732 7500 10333 7528
rect 9732 7488 9738 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10321 7491 10379 7497
rect 11606 7488 11612 7540
rect 11664 7528 11670 7540
rect 11882 7528 11888 7540
rect 11664 7500 11888 7528
rect 11664 7488 11670 7500
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13630 7488 13636 7500
rect 13688 7528 13694 7540
rect 19337 7531 19395 7537
rect 19337 7528 19349 7531
rect 13688 7500 19349 7528
rect 13688 7488 13694 7500
rect 19337 7497 19349 7500
rect 19383 7497 19395 7531
rect 19337 7491 19395 7497
rect 20898 7488 20904 7540
rect 20956 7528 20962 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20956 7500 21465 7528
rect 20956 7488 20962 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 9030 7460 9036 7472
rect 8991 7432 9036 7460
rect 9030 7420 9036 7432
rect 9088 7420 9094 7472
rect 14642 7460 14648 7472
rect 14603 7432 14648 7460
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 17034 7460 17040 7472
rect 16995 7432 17040 7460
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 19061 7463 19119 7469
rect 19061 7460 19073 7463
rect 18288 7432 19073 7460
rect 18288 7420 18294 7432
rect 19061 7429 19073 7432
rect 19107 7429 19119 7463
rect 19061 7423 19119 7429
rect 9677 7395 9735 7401
rect 8772 7364 9260 7392
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 2498 7284 2504 7336
rect 2556 7324 2562 7336
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2556 7296 2973 7324
rect 2556 7284 2562 7296
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 3237 7287 3295 7293
rect 4126 7296 4721 7324
rect 3252 7256 3280 7287
rect 2976 7228 3280 7256
rect 2976 7200 3004 7228
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 2869 7191 2927 7197
rect 2869 7188 2881 7191
rect 2547 7160 2881 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 2869 7157 2881 7160
rect 2915 7188 2927 7191
rect 2958 7188 2964 7200
rect 2915 7160 2964 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 4126 7188 4154 7296
rect 4709 7293 4721 7296
rect 4755 7324 4767 7327
rect 4893 7327 4951 7333
rect 4893 7324 4905 7327
rect 4755 7296 4905 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4893 7293 4905 7296
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 7834 7324 7840 7336
rect 7795 7296 7840 7324
rect 7653 7287 7711 7293
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7668 7256 7696 7287
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8938 7324 8944 7336
rect 8899 7296 8944 7324
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9232 7333 9260 7364
rect 9677 7361 9689 7395
rect 9723 7392 9735 7395
rect 11606 7392 11612 7404
rect 9723 7364 11612 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12986 7392 12992 7404
rect 12575 7364 12992 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14918 7392 14924 7404
rect 14139 7364 14924 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15286 7392 15292 7404
rect 15247 7364 15292 7392
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 18414 7392 18420 7404
rect 16531 7364 17540 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9950 7324 9956 7336
rect 9263 7296 9956 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 11054 7324 11060 7336
rect 11015 7296 11060 7324
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 11330 7324 11336 7336
rect 11291 7296 11336 7324
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 17512 7333 17540 7364
rect 17788 7364 18420 7392
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 17586 7324 17592 7336
rect 17543 7296 17592 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 11072 7256 11100 7284
rect 11514 7256 11520 7268
rect 7432 7228 11100 7256
rect 11475 7228 11520 7256
rect 7432 7216 7438 7228
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12676 7228 12721 7256
rect 12676 7216 12682 7228
rect 14182 7216 14188 7268
rect 14240 7256 14246 7268
rect 14240 7228 14285 7256
rect 14240 7216 14246 7228
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 15620 7228 16221 7256
rect 15620 7216 15626 7228
rect 16209 7225 16221 7228
rect 16255 7256 16267 7259
rect 16298 7256 16304 7268
rect 16255 7228 16304 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 17788 7265 17816 7364
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 20763 7395 20821 7401
rect 20763 7392 20775 7395
rect 18656 7364 20775 7392
rect 18656 7352 18662 7364
rect 20763 7361 20775 7364
rect 20809 7361 20821 7395
rect 20763 7355 20821 7361
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7324 19395 7327
rect 19613 7327 19671 7333
rect 19613 7324 19625 7327
rect 19383 7296 19625 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 19613 7293 19625 7296
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 20530 7284 20536 7336
rect 20588 7324 20594 7336
rect 20660 7327 20718 7333
rect 20660 7324 20672 7327
rect 20588 7296 20672 7324
rect 20588 7284 20594 7296
rect 20660 7293 20672 7296
rect 20706 7324 20718 7327
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20706 7296 21097 7324
rect 20706 7293 20718 7296
rect 20660 7287 20718 7293
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 16577 7259 16635 7265
rect 16577 7225 16589 7259
rect 16623 7256 16635 7259
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 16623 7228 17785 7256
rect 16623 7225 16635 7228
rect 16577 7219 16635 7225
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 18138 7256 18144 7268
rect 18099 7228 18144 7256
rect 17773 7219 17831 7225
rect 3476 7160 4154 7188
rect 3476 7148 3482 7160
rect 6178 7148 6184 7200
rect 6236 7188 6242 7200
rect 6546 7188 6552 7200
rect 6236 7160 6552 7188
rect 6236 7148 6242 7160
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 7650 7188 7656 7200
rect 7611 7160 7656 7188
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8260 7160 8401 7188
rect 8260 7148 8266 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8389 7151 8447 7157
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12636 7188 12664 7216
rect 12299 7160 12664 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 15841 7191 15899 7197
rect 15841 7188 15853 7191
rect 15804 7160 15853 7188
rect 15804 7148 15810 7160
rect 15841 7157 15853 7160
rect 15887 7188 15899 7191
rect 16592 7188 16620 7219
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 18233 7219 18291 7225
rect 15887 7160 16620 7188
rect 18248 7188 18276 7219
rect 18322 7216 18328 7268
rect 18380 7256 18386 7268
rect 18782 7256 18788 7268
rect 18380 7228 18644 7256
rect 18743 7228 18788 7256
rect 18380 7216 18386 7228
rect 18414 7188 18420 7200
rect 18248 7160 18420 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 18616 7188 18644 7228
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 18616 7160 19441 7188
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 20162 7188 20168 7200
rect 20123 7160 20168 7188
rect 19429 7151 19487 7157
rect 20162 7148 20168 7160
rect 20220 7148 20226 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 2280 6956 3801 6984
rect 2280 6944 2286 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 5258 6984 5264 6996
rect 5219 6956 5264 6984
rect 3789 6947 3847 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 5408 6956 7297 6984
rect 5408 6944 5414 6956
rect 7285 6953 7297 6956
rect 7331 6984 7343 6987
rect 7374 6984 7380 6996
rect 7331 6956 7380 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9088 6956 9413 6984
rect 9088 6944 9094 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9766 6984 9772 6996
rect 9727 6956 9772 6984
rect 9401 6947 9459 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 11054 6984 11060 6996
rect 10919 6956 11060 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 14090 6984 14096 6996
rect 14051 6956 14096 6984
rect 14090 6944 14096 6956
rect 14148 6984 14154 6996
rect 14461 6987 14519 6993
rect 14461 6984 14473 6987
rect 14148 6956 14473 6984
rect 14148 6944 14154 6956
rect 14461 6953 14473 6956
rect 14507 6953 14519 6987
rect 14461 6947 14519 6953
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 16669 6987 16727 6993
rect 16669 6984 16681 6987
rect 16540 6956 16681 6984
rect 16540 6944 16546 6956
rect 16669 6953 16681 6956
rect 16715 6953 16727 6987
rect 16669 6947 16727 6953
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 19843 6987 19901 6993
rect 19843 6984 19855 6987
rect 18564 6956 19855 6984
rect 18564 6944 18570 6956
rect 19843 6953 19855 6956
rect 19889 6953 19901 6987
rect 19843 6947 19901 6953
rect 2133 6919 2191 6925
rect 2133 6885 2145 6919
rect 2179 6916 2191 6919
rect 2498 6916 2504 6928
rect 2179 6888 2504 6916
rect 2179 6885 2191 6888
rect 2133 6879 2191 6885
rect 2498 6876 2504 6888
rect 2556 6916 2562 6928
rect 2777 6919 2835 6925
rect 2777 6916 2789 6919
rect 2556 6888 2789 6916
rect 2556 6876 2562 6888
rect 2777 6885 2789 6888
rect 2823 6916 2835 6919
rect 3421 6919 3479 6925
rect 3421 6916 3433 6919
rect 2823 6888 3433 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 3421 6885 3433 6888
rect 3467 6885 3479 6919
rect 5994 6916 6000 6928
rect 3421 6879 3479 6885
rect 4816 6888 6000 6916
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2996 6851 3054 6857
rect 2996 6848 3008 6851
rect 2740 6820 3008 6848
rect 2740 6808 2746 6820
rect 2996 6817 3008 6820
rect 3042 6848 3054 6851
rect 3694 6848 3700 6860
rect 3042 6820 3700 6848
rect 3042 6817 3054 6820
rect 2996 6811 3054 6817
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 4816 6857 4844 6888
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 6549 6919 6607 6925
rect 6549 6885 6561 6919
rect 6595 6916 6607 6919
rect 8294 6916 8300 6928
rect 6595 6888 8300 6916
rect 6595 6885 6607 6888
rect 6549 6879 6607 6885
rect 8294 6876 8300 6888
rect 8352 6916 8358 6928
rect 8662 6916 8668 6928
rect 8352 6888 8668 6916
rect 8352 6876 8358 6888
rect 8662 6876 8668 6888
rect 8720 6876 8726 6928
rect 11698 6916 11704 6928
rect 10152 6888 11704 6916
rect 10152 6860 10180 6888
rect 11698 6876 11704 6888
rect 11756 6916 11762 6928
rect 11756 6888 12020 6916
rect 11756 6876 11762 6888
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6817 4859 6851
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 4801 6811 4859 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7374 6848 7380 6860
rect 6840 6820 7380 6848
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 1544 6752 4261 6780
rect 1544 6740 1550 6752
rect 4249 6749 4261 6752
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 6840 6780 6868 6820
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7834 6848 7840 6860
rect 7747 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9548 6820 9965 6848
rect 9548 6808 9554 6820
rect 9953 6817 9965 6820
rect 9999 6817 10011 6851
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 9953 6811 10011 6817
rect 5132 6752 6868 6780
rect 7101 6783 7159 6789
rect 5132 6740 5138 6752
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7852 6780 7880 6808
rect 8110 6780 8116 6792
rect 7147 6752 7880 6780
rect 8023 6752 8116 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 8110 6740 8116 6752
rect 8168 6780 8174 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8168 6752 8401 6780
rect 8168 6740 8174 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 9968 6780 9996 6811
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 11790 6848 11796 6860
rect 11751 6820 11796 6848
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 11992 6857 12020 6888
rect 12912 6888 13584 6916
rect 12912 6860 12940 6888
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12023 6820 12541 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12529 6817 12541 6820
rect 12575 6848 12587 6851
rect 12894 6848 12900 6860
rect 12575 6820 12900 6848
rect 12575 6817 12587 6820
rect 12529 6811 12587 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13446 6848 13452 6860
rect 13403 6820 13452 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 13556 6857 13584 6888
rect 15562 6876 15568 6928
rect 15620 6916 15626 6928
rect 15794 6919 15852 6925
rect 15794 6916 15806 6919
rect 15620 6888 15806 6916
rect 15620 6876 15626 6888
rect 15794 6885 15806 6888
rect 15840 6885 15852 6919
rect 15794 6879 15852 6885
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 18325 6919 18383 6925
rect 18325 6916 18337 6919
rect 18288 6888 18337 6916
rect 18288 6876 18294 6888
rect 18325 6885 18337 6888
rect 18371 6885 18383 6919
rect 18325 6879 18383 6885
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 17862 6848 17868 6860
rect 14884 6820 17868 6848
rect 14884 6808 14890 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 19610 6808 19616 6860
rect 19668 6848 19674 6860
rect 19740 6851 19798 6857
rect 19740 6848 19752 6851
rect 19668 6820 19752 6848
rect 19668 6808 19674 6820
rect 19740 6817 19752 6820
rect 19786 6817 19798 6851
rect 19740 6811 19798 6817
rect 24581 6851 24639 6857
rect 24581 6817 24593 6851
rect 24627 6848 24639 6851
rect 24670 6848 24676 6860
rect 24627 6820 24676 6848
rect 24627 6817 24639 6820
rect 24581 6811 24639 6817
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 10686 6780 10692 6792
rect 9968 6752 10692 6780
rect 8389 6743 8447 6749
rect 10686 6740 10692 6752
rect 10744 6740 10750 6792
rect 12066 6780 12072 6792
rect 12027 6752 12072 6780
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 13630 6780 13636 6792
rect 13591 6752 13636 6780
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 15470 6780 15476 6792
rect 13786 6752 15476 6780
rect 3099 6715 3157 6721
rect 3099 6681 3111 6715
rect 3145 6712 3157 6715
rect 9030 6712 9036 6724
rect 3145 6684 9036 6712
rect 3145 6681 3157 6684
rect 3099 6675 3157 6681
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 13786 6712 13814 6752
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 19242 6780 19248 6792
rect 18279 6752 19248 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 14918 6712 14924 6724
rect 11572 6684 13814 6712
rect 14831 6684 14924 6712
rect 11572 6672 11578 6684
rect 14918 6672 14924 6684
rect 14976 6712 14982 6724
rect 18049 6715 18107 6721
rect 14976 6684 17448 6712
rect 14976 6672 14982 6684
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 4985 6647 5043 6653
rect 4985 6644 4997 6647
rect 2648 6616 4997 6644
rect 2648 6604 2654 6616
rect 4985 6613 4997 6616
rect 5031 6644 5043 6647
rect 5350 6644 5356 6656
rect 5031 6616 5356 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6604 6616 6837 6644
rect 6604 6604 6610 6616
rect 6825 6613 6837 6616
rect 6871 6644 6883 6647
rect 7101 6647 7159 6653
rect 7101 6644 7113 6647
rect 6871 6616 7113 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7101 6613 7113 6616
rect 7147 6613 7159 6647
rect 7101 6607 7159 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8938 6644 8944 6656
rect 7984 6616 8944 6644
rect 7984 6604 7990 6616
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 12986 6644 12992 6656
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 15804 6616 16405 6644
rect 15804 6604 15810 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 17420 6644 17448 6684
rect 18049 6681 18061 6715
rect 18095 6712 18107 6715
rect 18138 6712 18144 6724
rect 18095 6684 18144 6712
rect 18095 6681 18107 6684
rect 18049 6675 18107 6681
rect 18138 6672 18144 6684
rect 18196 6712 18202 6724
rect 18598 6712 18604 6724
rect 18196 6684 18604 6712
rect 18196 6672 18202 6684
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 18782 6712 18788 6724
rect 18743 6684 18788 6712
rect 18782 6672 18788 6684
rect 18840 6672 18846 6724
rect 24719 6647 24777 6653
rect 24719 6644 24731 6647
rect 17420 6616 24731 6644
rect 16393 6607 16451 6613
rect 24719 6613 24731 6616
rect 24765 6613 24777 6647
rect 24719 6607 24777 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 4065 6443 4123 6449
rect 4065 6440 4077 6443
rect 1452 6412 4077 6440
rect 1452 6400 1458 6412
rect 4065 6409 4077 6412
rect 4111 6409 4123 6443
rect 4065 6403 4123 6409
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 5132 6412 5365 6440
rect 5132 6400 5138 6412
rect 5353 6409 5365 6412
rect 5399 6409 5411 6443
rect 5353 6403 5411 6409
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5994 6440 6000 6452
rect 5675 6412 6000 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 7282 6440 7288 6452
rect 6687 6412 7288 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 6546 6372 6552 6384
rect 1903 6344 6552 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 3142 6304 3148 6316
rect 2639 6276 3004 6304
rect 3103 6276 3148 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 2976 6248 3004 6276
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3694 6304 3700 6316
rect 3655 6276 3700 6304
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 4614 6304 4620 6316
rect 4527 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6304 4678 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4672 6276 5273 6304
rect 4672 6264 4678 6276
rect 5261 6273 5273 6276
rect 5307 6304 5319 6307
rect 6086 6304 6092 6316
rect 5307 6276 6092 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1946 6236 1952 6248
rect 1719 6208 1952 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2498 6196 2504 6248
rect 2556 6236 2562 6248
rect 2685 6239 2743 6245
rect 2685 6236 2697 6239
rect 2556 6208 2697 6236
rect 2556 6196 2562 6208
rect 2685 6205 2697 6208
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 2958 6236 2964 6248
rect 2832 6208 2877 6236
rect 2919 6208 2964 6236
rect 2832 6196 2838 6208
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6656 6236 6684 6403
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 7892 6412 9045 6440
rect 7892 6400 7898 6412
rect 9033 6409 9045 6412
rect 9079 6440 9091 6443
rect 10134 6440 10140 6452
rect 9079 6412 10140 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 10134 6400 10140 6412
rect 10192 6440 10198 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10192 6412 10609 6440
rect 10192 6400 10198 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 15528 6412 17141 6440
rect 15528 6400 15534 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 19242 6440 19248 6452
rect 19203 6412 19248 6440
rect 17129 6403 17187 6409
rect 19242 6400 19248 6412
rect 19300 6440 19306 6452
rect 19935 6443 19993 6449
rect 19935 6440 19947 6443
rect 19300 6412 19947 6440
rect 19300 6400 19306 6412
rect 19935 6409 19947 6412
rect 19981 6409 19993 6443
rect 19935 6403 19993 6409
rect 20162 6400 20168 6452
rect 20220 6440 20226 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 20220 6412 20361 6440
rect 20220 6400 20226 6412
rect 20349 6409 20361 6412
rect 20395 6440 20407 6443
rect 27614 6440 27620 6452
rect 20395 6412 27620 6440
rect 20395 6409 20407 6412
rect 20349 6403 20407 6409
rect 27614 6400 27620 6412
rect 27672 6400 27678 6452
rect 7009 6375 7067 6381
rect 7009 6341 7021 6375
rect 7055 6372 7067 6375
rect 7926 6372 7932 6384
rect 7055 6344 7932 6372
rect 7055 6341 7067 6344
rect 7009 6335 7067 6341
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 9490 6372 9496 6384
rect 9451 6344 9496 6372
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 11333 6375 11391 6381
rect 11333 6341 11345 6375
rect 11379 6372 11391 6375
rect 13446 6372 13452 6384
rect 11379 6344 13452 6372
rect 11379 6341 11391 6344
rect 11333 6335 11391 6341
rect 13446 6332 13452 6344
rect 13504 6332 13510 6384
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8110 6304 8116 6316
rect 7883 6276 8116 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9088 6276 9689 6304
rect 9088 6264 9094 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 10134 6304 10140 6316
rect 10095 6276 10140 6304
rect 9677 6267 9735 6273
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11790 6304 11796 6316
rect 11747 6276 11796 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11790 6264 11796 6276
rect 11848 6304 11854 6316
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 11848 6276 14197 6304
rect 11848 6264 11854 6276
rect 14185 6273 14197 6276
rect 14231 6304 14243 6307
rect 15378 6304 15384 6316
rect 14231 6276 15384 6304
rect 14231 6273 14243 6276
rect 14185 6267 14243 6273
rect 6822 6236 6828 6248
rect 5767 6208 6684 6236
rect 6735 6208 6828 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 6822 6196 6828 6208
rect 6880 6236 6886 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 6880 6208 7297 6236
rect 6880 6196 6886 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 7285 6199 7343 6205
rect 10980 6208 11161 6236
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 6178 6168 6184 6180
rect 5500 6140 6184 6168
rect 5500 6128 5506 6140
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 8158 6171 8216 6177
rect 8158 6137 8170 6171
rect 8204 6137 8216 6171
rect 9769 6171 9827 6177
rect 8158 6131 8216 6137
rect 8956 6140 9628 6168
rect 1026 6060 1032 6112
rect 1084 6100 1090 6112
rect 1578 6100 1584 6112
rect 1084 6072 1584 6100
rect 1084 6060 1090 6072
rect 1578 6060 1584 6072
rect 1636 6100 1642 6112
rect 2133 6103 2191 6109
rect 2133 6100 2145 6103
rect 1636 6072 2145 6100
rect 1636 6060 1642 6072
rect 2133 6069 2145 6072
rect 2179 6069 2191 6103
rect 2133 6063 2191 6069
rect 4847 6103 4905 6109
rect 4847 6069 4859 6103
rect 4893 6100 4905 6103
rect 5074 6100 5080 6112
rect 4893 6072 5080 6100
rect 4893 6069 4905 6072
rect 4847 6063 4905 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6100 5411 6103
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 5399 6072 5917 6100
rect 5399 6069 5411 6072
rect 5353 6063 5411 6069
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 7742 6100 7748 6112
rect 7703 6072 7748 6100
rect 5905 6063 5963 6069
rect 7742 6060 7748 6072
rect 7800 6100 7806 6112
rect 8173 6100 8201 6131
rect 8956 6112 8984 6140
rect 7800 6072 8201 6100
rect 8757 6103 8815 6109
rect 7800 6060 7806 6072
rect 8757 6069 8769 6103
rect 8803 6100 8815 6103
rect 8938 6100 8944 6112
rect 8803 6072 8944 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9600 6100 9628 6140
rect 9769 6137 9781 6171
rect 9815 6137 9827 6171
rect 9769 6131 9827 6137
rect 9784 6100 9812 6131
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10980 6177 11008 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12299 6208 12725 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12894 6236 12900 6248
rect 12855 6208 12900 6236
rect 12713 6199 12771 6205
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 10100 6140 10977 6168
rect 10100 6128 10106 6140
rect 10965 6137 10977 6140
rect 11011 6137 11023 6171
rect 12728 6168 12756 6199
rect 12894 6196 12900 6208
rect 12952 6236 12958 6248
rect 14384 6245 14412 6276
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18196 6276 18613 6304
rect 18196 6264 18202 6276
rect 18601 6273 18613 6276
rect 18647 6304 18659 6307
rect 18782 6304 18788 6316
rect 18647 6276 18788 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19610 6304 19616 6316
rect 19571 6276 19616 6304
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 12952 6208 13829 6236
rect 12952 6196 12958 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14826 6236 14832 6248
rect 14787 6208 14832 6236
rect 14369 6199 14427 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6236 15163 6239
rect 15930 6236 15936 6248
rect 15151 6208 15936 6236
rect 15151 6205 15163 6208
rect 15105 6199 15163 6205
rect 15930 6196 15936 6208
rect 15988 6196 15994 6248
rect 19864 6239 19922 6245
rect 19864 6205 19876 6239
rect 19910 6236 19922 6239
rect 20162 6236 20168 6248
rect 19910 6208 20168 6236
rect 19910 6205 19922 6208
rect 19864 6199 19922 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 13078 6168 13084 6180
rect 12728 6140 13084 6168
rect 10965 6131 11023 6137
rect 13078 6128 13084 6140
rect 13136 6168 13142 6180
rect 15654 6168 15660 6180
rect 13136 6140 15660 6168
rect 13136 6128 13142 6140
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 16254 6171 16312 6177
rect 16254 6137 16266 6171
rect 16300 6137 16312 6171
rect 16254 6131 16312 6137
rect 17865 6171 17923 6177
rect 17865 6137 17877 6171
rect 17911 6168 17923 6171
rect 18322 6168 18328 6180
rect 17911 6140 18328 6168
rect 17911 6137 17923 6140
rect 17865 6131 17923 6137
rect 9600 6072 9812 6100
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 12308 6072 12541 6100
rect 12308 6060 12314 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 12529 6063 12587 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 15470 6060 15476 6072
rect 15528 6100 15534 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15528 6072 15761 6100
rect 15528 6060 15534 6072
rect 15749 6069 15761 6072
rect 15795 6100 15807 6103
rect 16269 6100 16297 6131
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 18417 6171 18475 6177
rect 18417 6137 18429 6171
rect 18463 6168 18475 6171
rect 18598 6168 18604 6180
rect 18463 6140 18604 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 15795 6072 16297 6100
rect 16853 6103 16911 6109
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 17770 6100 17776 6112
rect 16899 6072 17776 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 24670 6100 24676 6112
rect 24583 6072 24676 6100
rect 24670 6060 24676 6072
rect 24728 6100 24734 6112
rect 26878 6100 26884 6112
rect 24728 6072 26884 6100
rect 24728 6060 24734 6072
rect 26878 6060 26884 6072
rect 26936 6060 26942 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1673 5899 1731 5905
rect 1673 5896 1685 5899
rect 1544 5868 1685 5896
rect 1544 5856 1550 5868
rect 1673 5865 1685 5868
rect 1719 5865 1731 5899
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1673 5859 1731 5865
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2774 5896 2780 5908
rect 2735 5868 2780 5896
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 3108 5868 3157 5896
rect 3108 5856 3114 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 3145 5859 3203 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4948 5868 5089 5896
rect 4948 5856 4954 5868
rect 5077 5865 5089 5868
rect 5123 5896 5135 5899
rect 6454 5896 6460 5908
rect 5123 5868 6460 5896
rect 5123 5865 5135 5868
rect 5077 5859 5135 5865
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 7374 5896 7380 5908
rect 7335 5868 7380 5896
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 11609 5899 11667 5905
rect 8803 5868 9904 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9876 5840 9904 5868
rect 11609 5865 11621 5899
rect 11655 5896 11667 5899
rect 11698 5896 11704 5908
rect 11655 5868 11704 5896
rect 11655 5865 11667 5868
rect 11609 5859 11667 5865
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13955 5899 14013 5905
rect 13955 5896 13967 5899
rect 13044 5868 13967 5896
rect 13044 5856 13050 5868
rect 13955 5865 13967 5868
rect 14001 5865 14013 5899
rect 13955 5859 14013 5865
rect 14461 5899 14519 5905
rect 14461 5865 14473 5899
rect 14507 5896 14519 5899
rect 14826 5896 14832 5908
rect 14507 5868 14832 5896
rect 14507 5865 14519 5868
rect 14461 5859 14519 5865
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5490 5831 5548 5837
rect 5490 5828 5502 5831
rect 5316 5800 5502 5828
rect 5316 5788 5322 5800
rect 5490 5797 5502 5800
rect 5536 5797 5548 5831
rect 5490 5791 5548 5797
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 8158 5831 8216 5837
rect 8158 5828 8170 5831
rect 7800 5800 8170 5828
rect 7800 5788 7806 5800
rect 8158 5797 8170 5800
rect 8204 5797 8216 5831
rect 8158 5791 8216 5797
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 9214 5828 9220 5840
rect 8996 5800 9220 5828
rect 8996 5788 9002 5800
rect 9214 5788 9220 5800
rect 9272 5828 9278 5840
rect 9401 5831 9459 5837
rect 9401 5828 9413 5831
rect 9272 5800 9413 5828
rect 9272 5788 9278 5800
rect 9401 5797 9413 5800
rect 9447 5797 9459 5831
rect 9858 5828 9864 5840
rect 9771 5800 9864 5828
rect 9401 5791 9459 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 12390 5831 12448 5837
rect 12390 5828 12402 5831
rect 11940 5800 12402 5828
rect 11940 5788 11946 5800
rect 12390 5797 12402 5800
rect 12436 5797 12448 5831
rect 12390 5791 12448 5797
rect 1464 5763 1522 5769
rect 1464 5729 1476 5763
rect 1510 5760 1522 5763
rect 1762 5760 1768 5772
rect 1510 5732 1768 5760
rect 1510 5729 1522 5732
rect 1464 5723 1522 5729
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3418 5760 3424 5772
rect 3007 5732 3424 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4338 5760 4344 5772
rect 4111 5732 4344 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4338 5720 4344 5732
rect 4396 5760 4402 5772
rect 4982 5760 4988 5772
rect 4396 5732 4988 5760
rect 4396 5720 4402 5732
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5166 5760 5172 5772
rect 5127 5732 5172 5760
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 7650 5720 7656 5772
rect 7708 5760 7714 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7708 5732 7849 5760
rect 7708 5720 7714 5732
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 7837 5723 7895 5729
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 12066 5760 12072 5772
rect 12027 5732 12072 5760
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 13872 5732 13917 5760
rect 13872 5720 13878 5732
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 5132 5664 9781 5692
rect 5132 5652 5138 5664
rect 9769 5661 9781 5664
rect 9815 5692 9827 5695
rect 9950 5692 9956 5704
rect 9815 5664 9956 5692
rect 9815 5661 9827 5664
rect 9769 5655 9827 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 14476 5692 14504 5859
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 15930 5856 15936 5908
rect 15988 5896 15994 5908
rect 16485 5899 16543 5905
rect 16485 5896 16497 5899
rect 15988 5868 16497 5896
rect 15988 5856 15994 5868
rect 16485 5865 16497 5868
rect 16531 5865 16543 5899
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 16485 5859 16543 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 18340 5868 19564 5896
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 15657 5831 15715 5837
rect 15657 5828 15669 5831
rect 15436 5800 15669 5828
rect 15436 5788 15442 5800
rect 15657 5797 15669 5800
rect 15703 5828 15715 5831
rect 15746 5828 15752 5840
rect 15703 5800 15752 5828
rect 15703 5797 15715 5800
rect 15657 5791 15715 5797
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 17358 5831 17416 5837
rect 17358 5828 17370 5831
rect 17184 5800 17370 5828
rect 17184 5788 17190 5800
rect 17358 5797 17370 5800
rect 17404 5797 17416 5831
rect 17358 5791 17416 5797
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5760 16267 5763
rect 16482 5760 16488 5772
rect 16255 5732 16488 5760
rect 16255 5729 16267 5732
rect 16209 5723 16267 5729
rect 16482 5720 16488 5732
rect 16540 5760 16546 5772
rect 18340 5760 18368 5868
rect 19536 5840 19564 5868
rect 18598 5788 18604 5840
rect 18656 5828 18662 5840
rect 18969 5831 19027 5837
rect 18969 5828 18981 5831
rect 18656 5800 18981 5828
rect 18656 5788 18662 5800
rect 18969 5797 18981 5800
rect 19015 5797 19027 5831
rect 19518 5828 19524 5840
rect 19479 5800 19524 5828
rect 18969 5791 19027 5797
rect 19518 5788 19524 5800
rect 19576 5788 19582 5840
rect 16540 5732 18368 5760
rect 16540 5720 16546 5732
rect 15562 5692 15568 5704
rect 11388 5664 14504 5692
rect 15523 5664 15568 5692
rect 11388 5652 11394 5664
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17586 5692 17592 5704
rect 17083 5664 17592 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5692 18935 5695
rect 19794 5692 19800 5704
rect 18923 5664 19800 5692
rect 18923 5661 18935 5664
rect 18877 5655 18935 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 12989 5627 13047 5633
rect 12989 5593 13001 5627
rect 13035 5624 13047 5627
rect 14182 5624 14188 5636
rect 13035 5596 14188 5624
rect 13035 5593 13047 5596
rect 12989 5587 13047 5593
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 17957 5627 18015 5633
rect 17957 5593 17969 5627
rect 18003 5624 18015 5627
rect 18003 5596 18644 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 18616 5568 18644 5596
rect 6086 5556 6092 5568
rect 6047 5528 6092 5556
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 18598 5556 18604 5568
rect 18559 5528 18604 5556
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1535 5355 1593 5361
rect 1535 5352 1547 5355
rect 1452 5324 1547 5352
rect 1452 5312 1458 5324
rect 1535 5321 1547 5324
rect 1581 5321 1593 5355
rect 1535 5315 1593 5321
rect 1762 5312 1768 5364
rect 1820 5352 1826 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 1820 5324 2237 5352
rect 1820 5312 1826 5324
rect 2225 5321 2237 5324
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3660 5324 3801 5352
rect 3660 5312 3666 5324
rect 3789 5321 3801 5324
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7708 5324 8217 5352
rect 7708 5312 7714 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10008 5324 10885 5352
rect 10008 5312 10014 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 11425 5355 11483 5361
rect 11425 5321 11437 5355
rect 11471 5352 11483 5355
rect 12066 5352 12072 5364
rect 11471 5324 12072 5352
rect 11471 5321 11483 5324
rect 11425 5315 11483 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 15378 5352 15384 5364
rect 13872 5324 13917 5352
rect 15339 5324 15384 5352
rect 13872 5312 13878 5324
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 19794 5352 19800 5364
rect 19755 5324 19800 5352
rect 19794 5312 19800 5324
rect 19852 5352 19858 5364
rect 20119 5355 20177 5361
rect 20119 5352 20131 5355
rect 19852 5324 20131 5352
rect 19852 5312 19858 5324
rect 20119 5321 20131 5324
rect 20165 5321 20177 5355
rect 20119 5315 20177 5321
rect 3145 5287 3203 5293
rect 3145 5253 3157 5287
rect 3191 5284 3203 5287
rect 3878 5284 3884 5296
rect 3191 5256 3884 5284
rect 3191 5253 3203 5256
rect 3145 5247 3203 5253
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4709 5287 4767 5293
rect 4023 5256 4154 5284
rect 1118 5108 1124 5160
rect 1176 5148 1182 5160
rect 1432 5151 1490 5157
rect 1432 5148 1444 5151
rect 1176 5120 1444 5148
rect 1176 5108 1182 5120
rect 1432 5117 1444 5120
rect 1478 5148 1490 5151
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1478 5120 1869 5148
rect 1478 5117 1490 5120
rect 1432 5111 1490 5117
rect 1857 5117 1869 5120
rect 1903 5148 1915 5151
rect 1946 5148 1952 5160
rect 1903 5120 1952 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3602 5148 3608 5160
rect 3007 5120 3608 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 4023 5157 4051 5256
rect 4126 5216 4154 5256
rect 4709 5253 4721 5287
rect 4755 5284 4767 5287
rect 5258 5284 5264 5296
rect 4755 5256 5264 5284
rect 4755 5253 4767 5256
rect 4709 5247 4767 5253
rect 5258 5244 5264 5256
rect 5316 5284 5322 5296
rect 6181 5287 6239 5293
rect 6181 5284 6193 5287
rect 5316 5256 6193 5284
rect 5316 5244 5322 5256
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4126 5188 4537 5216
rect 4525 5185 4537 5188
rect 4571 5216 4583 5219
rect 5534 5216 5540 5228
rect 4571 5188 5540 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 4008 5151 4066 5157
rect 4008 5117 4020 5151
rect 4054 5117 4066 5151
rect 4008 5111 4066 5117
rect 4890 5108 4896 5160
rect 4948 5148 4954 5160
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4948 5120 4997 5148
rect 4948 5108 4954 5120
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 2038 5040 2044 5092
rect 2096 5080 2102 5092
rect 4709 5083 4767 5089
rect 4709 5080 4721 5083
rect 2096 5052 4721 5080
rect 2096 5040 2102 5052
rect 4709 5049 4721 5052
rect 4755 5080 4767 5083
rect 4801 5083 4859 5089
rect 4801 5080 4813 5083
rect 4755 5052 4813 5080
rect 4755 5049 4767 5052
rect 4709 5043 4767 5049
rect 4801 5049 4813 5052
rect 4847 5049 4859 5083
rect 4801 5043 4859 5049
rect 5326 5083 5384 5089
rect 5326 5049 5338 5083
rect 5372 5080 5384 5083
rect 5644 5080 5672 5256
rect 6181 5253 6193 5256
rect 6227 5284 6239 5287
rect 7742 5284 7748 5296
rect 6227 5256 7748 5284
rect 6227 5253 6239 5256
rect 6181 5247 6239 5253
rect 7742 5244 7748 5256
rect 7800 5284 7806 5296
rect 7837 5287 7895 5293
rect 7837 5284 7849 5287
rect 7800 5256 7849 5284
rect 7800 5244 7806 5256
rect 7837 5253 7849 5256
rect 7883 5284 7895 5287
rect 9493 5287 9551 5293
rect 9493 5284 9505 5287
rect 7883 5256 9505 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 9493 5253 9505 5256
rect 9539 5284 9551 5287
rect 11882 5284 11888 5296
rect 9539 5256 11888 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 6914 5216 6920 5228
rect 6827 5188 6920 5216
rect 6914 5176 6920 5188
rect 6972 5216 6978 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 6972 5188 8677 5216
rect 6972 5176 6978 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8456 5151 8514 5157
rect 8456 5117 8468 5151
rect 8502 5148 8514 5151
rect 8502 5120 8984 5148
rect 8502 5117 8514 5120
rect 8456 5111 8514 5117
rect 6086 5080 6092 5092
rect 5372 5052 5672 5080
rect 5736 5052 6092 5080
rect 5372 5049 5384 5052
rect 5326 5043 5384 5049
rect 3418 5012 3424 5024
rect 3379 4984 3424 5012
rect 3418 4972 3424 4984
rect 3476 4972 3482 5024
rect 4111 5015 4169 5021
rect 4111 4981 4123 5015
rect 4157 5012 4169 5015
rect 4522 5012 4528 5024
rect 4157 4984 4528 5012
rect 4157 4981 4169 4984
rect 4111 4975 4169 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5736 5012 5764 5052
rect 6086 5040 6092 5052
rect 6144 5080 6150 5092
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 6144 5052 6561 5080
rect 6144 5040 6150 5052
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 7002 5083 7060 5089
rect 7002 5049 7014 5083
rect 7048 5049 7060 5083
rect 7558 5080 7564 5092
rect 7519 5052 7564 5080
rect 7002 5043 7060 5049
rect 4948 4984 5764 5012
rect 5905 5015 5963 5021
rect 4948 4972 4954 4984
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 5994 5012 6000 5024
rect 5951 4984 6000 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6564 5012 6592 5043
rect 7024 5012 7052 5043
rect 7558 5040 7564 5052
rect 7616 5040 7622 5092
rect 8956 5024 8984 5120
rect 9600 5080 9628 5256
rect 11882 5244 11888 5256
rect 11940 5284 11946 5296
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 11940 5256 12173 5284
rect 11940 5244 11946 5256
rect 12161 5253 12173 5256
rect 12207 5284 12219 5287
rect 12618 5284 12624 5296
rect 12207 5256 12624 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 12618 5244 12624 5256
rect 12676 5244 12682 5296
rect 20533 5287 20591 5293
rect 20533 5253 20545 5287
rect 20579 5284 20591 5287
rect 21634 5284 21640 5296
rect 20579 5256 21640 5284
rect 20579 5253 20591 5256
rect 20533 5247 20591 5253
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 9766 5216 9772 5228
rect 9723 5188 9772 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 10192 5188 12817 5216
rect 10192 5176 10198 5188
rect 12805 5185 12817 5188
rect 12851 5216 12863 5219
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 12851 5188 14105 5216
rect 12851 5185 12863 5188
rect 12805 5179 12863 5185
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 14734 5216 14740 5228
rect 14139 5188 14740 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18748 5188 18797 5216
rect 18748 5176 18754 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 10686 5148 10692 5160
rect 10643 5120 10692 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 10744 5120 12265 5148
rect 10744 5108 10750 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 15105 5151 15163 5157
rect 15105 5117 15117 5151
rect 15151 5148 15163 5151
rect 15286 5148 15292 5160
rect 15151 5120 15292 5148
rect 15151 5117 15163 5120
rect 15105 5111 15163 5117
rect 15286 5108 15292 5120
rect 15344 5148 15350 5160
rect 15933 5151 15991 5157
rect 15933 5148 15945 5151
rect 15344 5120 15945 5148
rect 15344 5108 15350 5120
rect 15933 5117 15945 5120
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 20048 5151 20106 5157
rect 20048 5117 20060 5151
rect 20094 5148 20106 5151
rect 20548 5148 20576 5247
rect 21634 5244 21640 5256
rect 21692 5284 21698 5296
rect 27614 5284 27620 5296
rect 21692 5256 27620 5284
rect 21692 5244 21698 5256
rect 27614 5244 27620 5256
rect 27672 5244 27678 5296
rect 20094 5120 20576 5148
rect 20094 5117 20106 5120
rect 20048 5111 20106 5117
rect 9998 5083 10056 5089
rect 9998 5080 10010 5083
rect 9600 5052 10010 5080
rect 9998 5049 10010 5052
rect 10044 5049 10056 5083
rect 12529 5083 12587 5089
rect 12529 5080 12541 5083
rect 9998 5043 10056 5049
rect 11716 5052 12541 5080
rect 8938 5012 8944 5024
rect 6564 4984 7052 5012
rect 8899 4984 8944 5012
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11716 5021 11744 5052
rect 12529 5049 12541 5052
rect 12575 5049 12587 5083
rect 12529 5043 12587 5049
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5080 12679 5083
rect 13449 5083 13507 5089
rect 13449 5080 13461 5083
rect 12667 5052 13461 5080
rect 12667 5049 12679 5052
rect 12621 5043 12679 5049
rect 13449 5049 13461 5052
rect 13495 5049 13507 5083
rect 14182 5080 14188 5092
rect 14143 5052 14188 5080
rect 13449 5043 13507 5049
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11572 4984 11713 5012
rect 11572 4972 11578 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12636 5012 12664 5043
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 14734 5080 14740 5092
rect 14695 5052 14740 5080
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 16254 5083 16312 5089
rect 16254 5080 16266 5083
rect 15764 5052 16266 5080
rect 12299 4984 12664 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 15764 5021 15792 5052
rect 16254 5049 16266 5052
rect 16300 5080 16312 5083
rect 17126 5080 17132 5092
rect 16300 5052 17132 5080
rect 16300 5049 16312 5052
rect 16254 5043 16312 5049
rect 17126 5040 17132 5052
rect 17184 5040 17190 5092
rect 18506 5080 18512 5092
rect 18467 5052 18512 5080
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 18598 5040 18604 5092
rect 18656 5080 18662 5092
rect 18656 5052 18749 5080
rect 18656 5040 18662 5052
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15528 4984 15761 5012
rect 15528 4972 15534 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 16850 5012 16856 5024
rect 16811 4984 16856 5012
rect 15749 4975 15807 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18325 5015 18383 5021
rect 18325 4981 18337 5015
rect 18371 5012 18383 5015
rect 18616 5012 18644 5040
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 18371 4984 19441 5012
rect 18371 4981 18383 4984
rect 18325 4975 18383 4981
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 19429 4975 19487 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 1535 4811 1593 4817
rect 1535 4808 1547 4811
rect 1360 4780 1547 4808
rect 1360 4768 1366 4780
rect 1535 4777 1547 4780
rect 1581 4777 1593 4811
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 1535 4771 1593 4777
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5224 4780 5825 4808
rect 5224 4768 5230 4780
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 7469 4811 7527 4817
rect 7469 4808 7481 4811
rect 5813 4771 5871 4777
rect 7116 4780 7481 4808
rect 5537 4743 5595 4749
rect 5537 4709 5549 4743
rect 5583 4740 5595 4743
rect 6454 4740 6460 4752
rect 5583 4712 6460 4740
rect 5583 4709 5595 4712
rect 5537 4703 5595 4709
rect 6454 4700 6460 4712
rect 6512 4740 6518 4752
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 6512 4712 6561 4740
rect 6512 4700 6518 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 7116 4749 7144 4780
rect 7469 4777 7481 4780
rect 7515 4808 7527 4811
rect 7558 4808 7564 4820
rect 7515 4780 7564 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 9824 4780 10241 4808
rect 9824 4768 9830 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 12250 4808 12256 4820
rect 12207 4780 12256 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12618 4808 12624 4820
rect 12579 4780 12624 4808
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14461 4811 14519 4817
rect 14461 4808 14473 4811
rect 14240 4780 14473 4808
rect 14240 4768 14246 4780
rect 14461 4777 14473 4780
rect 14507 4777 14519 4811
rect 14461 4771 14519 4777
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 15562 4808 15568 4820
rect 15151 4780 15568 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 18506 4808 18512 4820
rect 18467 4780 18512 4808
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 7101 4743 7159 4749
rect 7101 4740 7113 4743
rect 6972 4712 7113 4740
rect 6972 4700 6978 4712
rect 7101 4709 7113 4712
rect 7147 4709 7159 4743
rect 9858 4740 9864 4752
rect 9819 4712 9864 4740
rect 7101 4703 7159 4709
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 10597 4743 10655 4749
rect 10597 4709 10609 4743
rect 10643 4740 10655 4743
rect 10686 4740 10692 4752
rect 10643 4712 10692 4740
rect 10643 4709 10655 4712
rect 10597 4703 10655 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1670 4672 1676 4684
rect 1510 4644 1676 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1670 4632 1676 4644
rect 1728 4672 1734 4684
rect 2130 4672 2136 4684
rect 1728 4644 2136 4672
rect 1728 4632 1734 4644
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7984 4644 8033 4672
rect 7984 4632 7990 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8021 4635 8079 4641
rect 8294 4632 8300 4644
rect 8352 4672 8358 4684
rect 8570 4672 8576 4684
rect 8352 4644 8576 4672
rect 8352 4632 8358 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 10042 4672 10048 4684
rect 8803 4644 10048 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 12268 4681 12296 4768
rect 15470 4700 15476 4752
rect 15528 4740 15534 4752
rect 15702 4743 15760 4749
rect 15702 4740 15714 4743
rect 15528 4712 15714 4740
rect 15528 4700 15534 4712
rect 15702 4709 15714 4712
rect 15748 4709 15760 4743
rect 15702 4703 15760 4709
rect 16850 4700 16856 4752
rect 16908 4740 16914 4752
rect 17402 4740 17408 4752
rect 16908 4712 17408 4740
rect 16908 4700 16914 4712
rect 17402 4700 17408 4712
rect 17460 4740 17466 4752
rect 17497 4743 17555 4749
rect 17497 4740 17509 4743
rect 17460 4712 17509 4740
rect 17460 4700 17466 4712
rect 17497 4709 17509 4712
rect 17543 4709 17555 4743
rect 17497 4703 17555 4709
rect 18322 4700 18328 4752
rect 18380 4740 18386 4752
rect 18877 4743 18935 4749
rect 18877 4740 18889 4743
rect 18380 4712 18889 4740
rect 18380 4700 18386 4712
rect 18877 4709 18889 4712
rect 18923 4709 18935 4743
rect 18877 4703 18935 4709
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4641 12311 4675
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 12253 4635 12311 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6328 4576 6469 4604
rect 6328 4564 6334 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 6457 4567 6515 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10778 4604 10784 4616
rect 10739 4576 10784 4604
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 15378 4604 15384 4616
rect 15339 4576 15384 4604
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17678 4604 17684 4616
rect 17639 4576 17684 4604
rect 17405 4567 17463 4573
rect 8110 4536 8116 4548
rect 8071 4508 8116 4536
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 13173 4539 13231 4545
rect 13173 4505 13185 4539
rect 13219 4536 13231 4539
rect 14366 4536 14372 4548
rect 13219 4508 14372 4536
rect 13219 4505 13231 4508
rect 13173 4499 13231 4505
rect 14366 4496 14372 4508
rect 14424 4496 14430 4548
rect 17420 4536 17448 4567
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 17954 4536 17960 4548
rect 17420 4508 17960 4536
rect 17954 4496 17960 4508
rect 18012 4536 18018 4548
rect 18690 4536 18696 4548
rect 18012 4508 18696 4536
rect 18012 4496 18018 4508
rect 18690 4496 18696 4508
rect 18748 4496 18754 4548
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 14139 4471 14197 4477
rect 14139 4468 14151 4471
rect 11940 4440 14151 4468
rect 11940 4428 11946 4440
rect 14139 4437 14151 4440
rect 14185 4437 14197 4471
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 14139 4431 14197 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 6454 4264 6460 4276
rect 6415 4236 6460 4264
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 9214 4264 9220 4276
rect 8404 4236 8984 4264
rect 9175 4236 9220 4264
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 8404 4196 8432 4236
rect 5684 4168 8432 4196
rect 5684 4156 5690 4168
rect 8570 4156 8576 4208
rect 8628 4196 8634 4208
rect 8757 4199 8815 4205
rect 8757 4196 8769 4199
rect 8628 4168 8769 4196
rect 8628 4156 8634 4168
rect 8757 4165 8769 4168
rect 8803 4165 8815 4199
rect 8956 4196 8984 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 10502 4264 10508 4276
rect 9324 4236 10508 4264
rect 9324 4196 9352 4236
rect 10502 4224 10508 4236
rect 10560 4264 10566 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10560 4236 10793 4264
rect 10560 4224 10566 4236
rect 10781 4233 10793 4236
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12618 4264 12624 4276
rect 12299 4236 12624 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 13630 4264 13636 4276
rect 13591 4236 13636 4264
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 16298 4264 16304 4276
rect 16259 4236 16304 4264
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 17770 4264 17776 4276
rect 17731 4236 17776 4264
rect 17770 4224 17776 4236
rect 17828 4264 17834 4276
rect 18230 4264 18236 4276
rect 17828 4236 18236 4264
rect 17828 4224 17834 4236
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 8956 4168 9352 4196
rect 8757 4159 8815 4165
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7190 4128 7196 4140
rect 7151 4100 7196 4128
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 7984 4100 8401 4128
rect 7984 4088 7990 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9582 4128 9588 4140
rect 9447 4100 9588 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9582 4088 9588 4100
rect 9640 4128 9646 4140
rect 11882 4128 11888 4140
rect 9640 4100 11888 4128
rect 9640 4088 9646 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 13648 4128 13676 4224
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 15749 4199 15807 4205
rect 15749 4196 15761 4199
rect 15436 4168 15761 4196
rect 15436 4156 15442 4168
rect 15749 4165 15761 4168
rect 15795 4165 15807 4199
rect 15749 4159 15807 4165
rect 16482 4128 16488 4140
rect 12483 4100 13676 4128
rect 16443 4100 16488 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17678 4128 17684 4140
rect 17175 4100 17684 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17678 4088 17684 4100
rect 17736 4128 17742 4140
rect 18414 4128 18420 4140
rect 17736 4100 18420 4128
rect 17736 4088 17742 4100
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 24026 4088 24032 4140
rect 24084 4128 24090 4140
rect 24719 4131 24777 4137
rect 24719 4128 24731 4131
rect 24084 4100 24731 4128
rect 24084 4088 24090 4100
rect 24719 4097 24731 4100
rect 24765 4097 24777 4131
rect 24719 4091 24777 4097
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5316 4032 5825 4060
rect 5316 4020 5322 4032
rect 5813 4029 5825 4032
rect 5859 4060 5871 4063
rect 11400 4063 11458 4069
rect 5859 4032 6040 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6012 4004 6040 4032
rect 11400 4029 11412 4063
rect 11446 4060 11458 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11446 4032 11805 4060
rect 11446 4029 11458 4032
rect 11400 4023 11458 4029
rect 11793 4029 11805 4032
rect 11839 4060 11851 4063
rect 13630 4060 13636 4072
rect 11839 4032 13636 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 24632 4063 24690 4069
rect 24632 4029 24644 4063
rect 24678 4060 24690 4063
rect 24678 4032 25176 4060
rect 24678 4029 24690 4032
rect 24632 4023 24690 4029
rect 5902 3992 5908 4004
rect 5863 3964 5908 3992
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 5994 3952 6000 4004
rect 6052 3992 6058 4004
rect 7009 3995 7067 4001
rect 7009 3992 7021 3995
rect 6052 3964 7021 3992
rect 6052 3952 6058 3964
rect 7009 3961 7021 3964
rect 7055 3992 7067 3995
rect 7374 3992 7380 4004
rect 7055 3964 7380 3992
rect 7055 3961 7067 3964
rect 7009 3955 7067 3961
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3961 9551 3995
rect 10042 3992 10048 4004
rect 10003 3964 10048 3992
rect 9493 3955 9551 3961
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9508 3924 9536 3955
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 11609 3995 11667 4001
rect 11609 3992 11621 3995
rect 10192 3964 11621 3992
rect 10192 3952 10198 3964
rect 11609 3961 11621 3964
rect 11655 3961 11667 3995
rect 11609 3955 11667 3961
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 12758 3995 12816 4001
rect 12758 3992 12770 3995
rect 12676 3964 12770 3992
rect 12676 3952 12682 3964
rect 12758 3961 12770 3964
rect 12804 3961 12816 3995
rect 12758 3955 12816 3961
rect 12894 3952 12900 4004
rect 12952 3992 12958 4004
rect 14274 3992 14280 4004
rect 12952 3964 14280 3992
rect 12952 3952 12958 3964
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 14424 3964 14469 3992
rect 14424 3952 14430 3964
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14792 3964 14933 3992
rect 14792 3952 14798 3964
rect 14921 3961 14933 3964
rect 14967 3992 14979 3995
rect 16206 3992 16212 4004
rect 14967 3964 16212 3992
rect 14967 3961 14979 3964
rect 14921 3955 14979 3961
rect 16206 3952 16212 3964
rect 16264 3952 16270 4004
rect 16298 3952 16304 4004
rect 16356 3992 16362 4004
rect 16577 3995 16635 4001
rect 16577 3992 16589 3995
rect 16356 3964 16589 3992
rect 16356 3952 16362 3964
rect 16577 3961 16589 3964
rect 16623 3961 16635 3995
rect 18138 3992 18144 4004
rect 18099 3964 18144 3992
rect 16577 3955 16635 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 18288 3952 18294 3964
rect 9272 3896 9536 3924
rect 10505 3927 10563 3933
rect 9272 3884 9278 3896
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10686 3924 10692 3936
rect 10551 3896 10692 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10686 3884 10692 3896
rect 10744 3924 10750 3936
rect 11330 3924 11336 3936
rect 10744 3896 11336 3924
rect 10744 3884 10750 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 13354 3924 13360 3936
rect 13315 3896 13360 3924
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13998 3924 14004 3936
rect 13959 3896 14004 3924
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14182 3884 14188 3936
rect 14240 3924 14246 3936
rect 15381 3927 15439 3933
rect 15381 3924 15393 3927
rect 14240 3896 15393 3924
rect 14240 3884 14246 3896
rect 15381 3893 15393 3896
rect 15427 3924 15439 3927
rect 15470 3924 15476 3936
rect 15427 3896 15476 3924
rect 15427 3893 15439 3896
rect 15381 3887 15439 3893
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 25148 3933 25176 4032
rect 25133 3927 25191 3933
rect 25133 3893 25145 3927
rect 25179 3924 25191 3927
rect 27614 3924 27620 3936
rect 25179 3896 27620 3924
rect 25179 3893 25191 3896
rect 25133 3887 25191 3893
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 5491 3723 5549 3729
rect 5491 3689 5503 3723
rect 5537 3720 5549 3723
rect 5626 3720 5632 3732
rect 5537 3692 5632 3720
rect 5537 3689 5549 3692
rect 5491 3683 5549 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 5994 3720 6000 3732
rect 5859 3692 6000 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 5994 3680 6000 3692
rect 6052 3720 6058 3732
rect 7374 3720 7380 3732
rect 6052 3692 7144 3720
rect 7335 3692 7380 3720
rect 6052 3680 6058 3692
rect 5902 3612 5908 3664
rect 5960 3652 5966 3664
rect 6454 3652 6460 3664
rect 5960 3624 6460 3652
rect 5960 3612 5966 3624
rect 6454 3612 6460 3624
rect 6512 3652 6518 3664
rect 7116 3661 7144 3692
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 9401 3723 9459 3729
rect 9401 3689 9413 3723
rect 9447 3720 9459 3723
rect 9582 3720 9588 3732
rect 9447 3692 9588 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 12529 3723 12587 3729
rect 10428 3692 12020 3720
rect 6549 3655 6607 3661
rect 6549 3652 6561 3655
rect 6512 3624 6561 3652
rect 6512 3612 6518 3624
rect 6549 3621 6561 3624
rect 6595 3621 6607 3655
rect 6549 3615 6607 3621
rect 7101 3655 7159 3661
rect 7101 3621 7113 3655
rect 7147 3652 7159 3655
rect 7190 3652 7196 3664
rect 7147 3624 7196 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 8205 3655 8263 3661
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 9214 3652 9220 3664
rect 8251 3624 9220 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 9766 3652 9772 3664
rect 9324 3624 9772 3652
rect 1464 3587 1522 3593
rect 1464 3553 1476 3587
rect 1510 3584 1522 3587
rect 1762 3584 1768 3596
rect 1510 3556 1768 3584
rect 1510 3553 1522 3556
rect 1464 3547 1522 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 5350 3584 5356 3596
rect 5311 3556 5356 3584
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 8812 3556 8857 3584
rect 8812 3544 8818 3556
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 4387 3488 6469 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 6457 3485 6469 3488
rect 6503 3516 6515 3519
rect 6914 3516 6920 3528
rect 6503 3488 6920 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7248 3488 8125 3516
rect 7248 3476 7254 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 9324 3516 9352 3624
rect 9766 3612 9772 3624
rect 9824 3652 9830 3664
rect 9861 3655 9919 3661
rect 9861 3652 9873 3655
rect 9824 3624 9873 3652
rect 9824 3612 9830 3624
rect 9861 3621 9873 3624
rect 9907 3621 9919 3655
rect 9861 3615 9919 3621
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10428 3661 10456 3692
rect 10413 3655 10471 3661
rect 10413 3652 10425 3655
rect 10100 3624 10425 3652
rect 10100 3612 10106 3624
rect 10413 3621 10425 3624
rect 10459 3621 10471 3655
rect 11422 3652 11428 3664
rect 11383 3624 11428 3652
rect 10413 3615 10471 3621
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 11992 3661 12020 3692
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 12618 3720 12624 3732
rect 12575 3692 12624 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 14182 3720 14188 3732
rect 12676 3692 14188 3720
rect 12676 3680 12682 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14277 3723 14335 3729
rect 14277 3689 14289 3723
rect 14323 3720 14335 3723
rect 14366 3720 14372 3732
rect 14323 3692 14372 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14884 3692 15025 3720
rect 14884 3680 14890 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 15378 3720 15384 3732
rect 15339 3692 15384 3720
rect 15013 3683 15071 3689
rect 11977 3655 12035 3661
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 12894 3652 12900 3664
rect 12023 3624 12900 3652
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 12989 3655 13047 3661
rect 12989 3621 13001 3655
rect 13035 3652 13047 3655
rect 13354 3652 13360 3664
rect 13035 3624 13360 3652
rect 13035 3621 13047 3624
rect 12989 3615 13047 3621
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 13541 3655 13599 3661
rect 13541 3621 13553 3655
rect 13587 3652 13599 3655
rect 14734 3652 14740 3664
rect 13587 3624 14740 3652
rect 13587 3621 13599 3624
rect 13541 3615 13599 3621
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 15028 3652 15056 3683
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 16482 3720 16488 3732
rect 16443 3692 16488 3720
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 17954 3720 17960 3732
rect 17915 3692 17960 3720
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 18196 3692 18245 3720
rect 18196 3680 18202 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 15470 3652 15476 3664
rect 15028 3624 15476 3652
rect 15470 3612 15476 3624
rect 15528 3652 15534 3664
rect 17586 3652 17592 3664
rect 15528 3624 17356 3652
rect 17547 3624 17592 3652
rect 15528 3612 15534 3624
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14332 3556 14565 3584
rect 14332 3544 14338 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 15562 3584 15568 3596
rect 15523 3556 15568 3584
rect 14553 3547 14611 3553
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 15764 3593 15792 3624
rect 15749 3587 15807 3593
rect 15749 3553 15761 3587
rect 15795 3553 15807 3587
rect 17126 3584 17132 3596
rect 17087 3556 17132 3584
rect 15749 3547 15807 3553
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 17328 3593 17356 3624
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 17313 3587 17371 3593
rect 17313 3553 17325 3587
rect 17359 3584 17371 3587
rect 17402 3584 17408 3596
rect 17359 3556 17408 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18414 3584 18420 3596
rect 18375 3556 18420 3584
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 8352 3488 9352 3516
rect 9769 3519 9827 3525
rect 8352 3476 8358 3488
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 10686 3516 10692 3528
rect 9815 3488 10692 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11698 3516 11704 3528
rect 11379 3488 11704 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 1535 3451 1593 3457
rect 1535 3417 1547 3451
rect 1581 3448 1593 3451
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 1581 3420 7757 3448
rect 1581 3417 1593 3420
rect 1535 3411 1593 3417
rect 7745 3417 7757 3420
rect 7791 3448 7803 3451
rect 7834 3448 7840 3460
rect 7791 3420 7840 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 10134 3448 10140 3460
rect 9508 3420 10140 3448
rect 6270 3380 6276 3392
rect 6183 3352 6276 3380
rect 6270 3340 6276 3352
rect 6328 3380 6334 3392
rect 9508 3380 9536 3420
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 18138 3448 18144 3460
rect 12768 3420 18144 3448
rect 12768 3408 12774 3420
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 6328 3352 9536 3380
rect 6328 3340 6334 3352
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 9916 3352 10701 3380
rect 9916 3340 9922 3352
rect 10689 3349 10701 3352
rect 10735 3349 10747 3383
rect 10689 3343 10747 3349
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 18555 3383 18613 3389
rect 18555 3380 18567 3383
rect 17552 3352 18567 3380
rect 17552 3340 17558 3352
rect 18555 3349 18567 3352
rect 18601 3349 18613 3383
rect 18555 3343 18613 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1820 3148 1869 3176
rect 1820 3136 1826 3148
rect 1857 3145 1869 3148
rect 1903 3145 1915 3179
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 1857 3139 1915 3145
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 6454 3176 6460 3188
rect 6415 3148 6460 3176
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6972 3148 7021 3176
rect 6972 3136 6978 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9214 3176 9220 3188
rect 8895 3148 9220 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 9824 3148 10333 3176
rect 9824 3136 9830 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10321 3139 10379 3145
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 11664 3148 12173 3176
rect 11664 3136 11670 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 13081 3179 13139 3185
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13354 3176 13360 3188
rect 13127 3148 13360 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 4847 3111 4905 3117
rect 4847 3077 4859 3111
rect 4893 3108 4905 3111
rect 9858 3108 9864 3120
rect 4893 3080 9864 3108
rect 4893 3077 4905 3080
rect 4847 3071 4905 3077
rect 1535 3043 1593 3049
rect 1535 3009 1547 3043
rect 1581 3040 1593 3043
rect 7558 3040 7564 3052
rect 1581 3012 7564 3040
rect 1581 3009 1593 3012
rect 1535 3003 1593 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 7834 3040 7840 3052
rect 7795 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 8754 3040 8760 3052
rect 8527 3012 8760 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9416 3049 9444 3080
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 9953 3111 10011 3117
rect 9953 3077 9965 3111
rect 9999 3108 10011 3111
rect 10134 3108 10140 3120
rect 9999 3080 10140 3108
rect 9999 3077 10011 3080
rect 9953 3071 10011 3077
rect 10134 3068 10140 3080
rect 10192 3108 10198 3120
rect 10962 3108 10968 3120
rect 10192 3080 10968 3108
rect 10192 3068 10198 3080
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3040 10931 3043
rect 11514 3040 11520 3052
rect 10919 3012 11520 3040
rect 10919 3009 10931 3012
rect 10873 3003 10931 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11698 3040 11704 3052
rect 11659 3012 11704 3040
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 106 2932 112 2984
rect 164 2972 170 2984
rect 1432 2975 1490 2981
rect 1432 2972 1444 2975
rect 164 2944 1444 2972
rect 164 2932 170 2944
rect 1432 2941 1444 2944
rect 1478 2972 1490 2975
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 1478 2944 2237 2972
rect 1478 2941 1490 2944
rect 1432 2935 1490 2941
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4744 2975 4802 2981
rect 4744 2972 4756 2975
rect 4663 2944 4756 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 4744 2941 4756 2944
rect 4790 2972 4802 2975
rect 5626 2972 5632 2984
rect 4790 2944 5632 2972
rect 4790 2941 4802 2944
rect 4744 2935 4802 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 5788 2975 5846 2981
rect 5788 2941 5800 2975
rect 5834 2972 5846 2975
rect 5994 2972 6000 2984
rect 5834 2944 6000 2972
rect 5834 2941 5846 2944
rect 5788 2935 5846 2941
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 12176 2972 12204 3139
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 14829 3179 14887 3185
rect 14829 3176 14841 3179
rect 13504 3148 14841 3176
rect 13504 3136 13510 3148
rect 14829 3145 14841 3148
rect 14875 3145 14887 3179
rect 14829 3139 14887 3145
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3108 12679 3111
rect 13722 3108 13728 3120
rect 12667 3080 13728 3108
rect 12667 3077 12679 3080
rect 12621 3071 12679 3077
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 12952 3012 13369 3040
rect 12952 3000 12958 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12176 2944 12449 2972
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 14550 2972 14556 2984
rect 13955 2944 14556 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 14844 2972 14872 3139
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16025 3179 16083 3185
rect 16025 3176 16037 3179
rect 15620 3148 16037 3176
rect 15620 3136 15626 3148
rect 16025 3145 16037 3148
rect 16071 3145 16083 3179
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 16025 3139 16083 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17460 3148 17509 3176
rect 17460 3136 17466 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 17497 3139 17555 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14844 2944 15025 2972
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 15013 2935 15071 2941
rect 15470 2932 15476 2944
rect 15528 2972 15534 2984
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 15528 2944 16405 2972
rect 15528 2932 15534 2944
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16393 2935 16451 2941
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2972 16635 2975
rect 17494 2972 17500 2984
rect 16623 2944 17500 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 17494 2932 17500 2944
rect 17552 2932 17558 2984
rect 3835 2907 3893 2913
rect 3835 2873 3847 2907
rect 3881 2904 3893 2907
rect 7653 2907 7711 2913
rect 3881 2876 7604 2904
rect 3881 2873 3893 2876
rect 3835 2867 3893 2873
rect 3605 2839 3663 2845
rect 3605 2805 3617 2839
rect 3651 2836 3663 2839
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 3651 2808 4261 2836
rect 3651 2805 3663 2808
rect 3605 2799 3663 2805
rect 4249 2805 4261 2808
rect 4295 2836 4307 2839
rect 4430 2836 4436 2848
rect 4295 2808 4436 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 5859 2839 5917 2845
rect 5859 2836 5871 2839
rect 5776 2808 5871 2836
rect 5776 2796 5782 2808
rect 5859 2805 5871 2808
rect 5905 2805 5917 2839
rect 7576 2836 7604 2876
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 7929 2907 7987 2913
rect 7929 2904 7941 2907
rect 7699 2876 7941 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 7929 2873 7941 2876
rect 7975 2904 7987 2907
rect 8294 2904 8300 2916
rect 7975 2876 8300 2904
rect 7975 2873 7987 2876
rect 7929 2867 7987 2873
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 9493 2907 9551 2913
rect 9493 2873 9505 2907
rect 9539 2904 9551 2907
rect 11514 2904 11520 2916
rect 9539 2876 11520 2904
rect 9539 2873 9551 2876
rect 9493 2867 9551 2873
rect 8570 2836 8576 2848
rect 7576 2808 8576 2836
rect 5859 2799 5917 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9217 2839 9275 2845
rect 9217 2836 9229 2839
rect 8812 2808 9229 2836
rect 8812 2796 8818 2808
rect 9217 2805 9229 2808
rect 9263 2836 9275 2839
rect 9508 2836 9536 2867
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 15378 2904 15384 2916
rect 14200 2876 15384 2904
rect 9263 2808 9536 2836
rect 14093 2839 14151 2845
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 14200 2836 14228 2876
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 14550 2836 14556 2848
rect 14139 2808 14228 2836
rect 14511 2808 14556 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 15286 2836 15292 2848
rect 15247 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 16758 2836 16764 2848
rect 16719 2808 16764 2836
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 7156 2604 7297 2632
rect 7156 2592 7162 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 7742 2632 7748 2644
rect 7703 2604 7748 2632
rect 7285 2595 7343 2601
rect 4709 2567 4767 2573
rect 4709 2533 4721 2567
rect 4755 2564 4767 2567
rect 7190 2564 7196 2576
rect 4755 2536 7196 2564
rect 4755 2533 4767 2536
rect 4709 2527 4767 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2496 3086 2499
rect 3510 2496 3516 2508
rect 3074 2468 3516 2496
rect 3074 2465 3086 2468
rect 3028 2459 3086 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4500 2499 4558 2505
rect 4500 2465 4512 2499
rect 4546 2496 4558 2499
rect 4890 2496 4896 2508
rect 4546 2468 4896 2496
rect 4546 2465 4558 2468
rect 4500 2459 4558 2465
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5718 2496 5724 2508
rect 5679 2468 5724 2496
rect 5718 2456 5724 2468
rect 5776 2496 5782 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5776 2468 6285 2496
rect 5776 2456 5782 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 7208 2428 7236 2524
rect 7300 2496 7328 2595
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8754 2632 8760 2644
rect 8715 2604 8760 2632
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 11471 2635 11529 2641
rect 11471 2632 11483 2635
rect 10744 2604 11483 2632
rect 10744 2592 10750 2604
rect 11471 2601 11483 2604
rect 11517 2601 11529 2635
rect 11471 2595 11529 2601
rect 15657 2635 15715 2641
rect 15657 2601 15669 2635
rect 15703 2632 15715 2635
rect 17678 2632 17684 2644
rect 15703 2604 17684 2632
rect 15703 2601 15715 2604
rect 15657 2595 15715 2601
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18463 2635 18521 2641
rect 18463 2632 18475 2635
rect 18196 2604 18475 2632
rect 18196 2592 18202 2604
rect 18463 2601 18475 2604
rect 18509 2601 18521 2635
rect 18463 2595 18521 2601
rect 20211 2635 20269 2641
rect 20211 2601 20223 2635
rect 20257 2632 20269 2635
rect 20622 2632 20628 2644
rect 20257 2604 20628 2632
rect 20257 2601 20269 2604
rect 20211 2595 20269 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 7760 2564 7788 2592
rect 8158 2567 8216 2573
rect 8158 2564 8170 2567
rect 7760 2536 8170 2564
rect 8158 2533 8170 2536
rect 8204 2533 8216 2567
rect 8158 2527 8216 2533
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 9953 2567 10011 2573
rect 9953 2564 9965 2567
rect 9631 2536 9965 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 9953 2533 9965 2536
rect 9999 2564 10011 2567
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 9999 2536 12633 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 12621 2533 12633 2536
rect 12667 2533 12679 2567
rect 17494 2564 17500 2576
rect 17455 2536 17500 2564
rect 12621 2527 12679 2533
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 19116 2536 23121 2564
rect 19116 2524 19122 2536
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 7300 2468 7849 2496
rect 7837 2465 7849 2468
rect 7883 2465 7895 2499
rect 7837 2459 7895 2465
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 11400 2499 11458 2505
rect 8628 2468 9536 2496
rect 8628 2456 8634 2468
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 7208 2400 9045 2428
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9508 2428 9536 2468
rect 11400 2465 11412 2499
rect 11446 2465 11458 2499
rect 11400 2459 11458 2465
rect 9858 2428 9864 2440
rect 9508 2400 9864 2428
rect 9033 2391 9091 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11415 2428 11443 2459
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 12437 2499 12495 2505
rect 12437 2496 12449 2499
rect 11572 2468 12449 2496
rect 11572 2456 11578 2468
rect 12437 2465 12449 2468
rect 12483 2496 12495 2499
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12483 2468 12725 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13688 2468 14197 2496
rect 13688 2456 13694 2468
rect 14185 2465 14197 2468
rect 14231 2496 14243 2499
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14231 2468 14749 2496
rect 14231 2465 14243 2468
rect 14185 2459 14243 2465
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 15519 2468 16160 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 11790 2428 11796 2440
rect 11415 2400 11796 2428
rect 11790 2388 11796 2400
rect 11848 2428 11854 2440
rect 14550 2428 14556 2440
rect 11848 2400 14556 2428
rect 11848 2388 11854 2400
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 3099 2363 3157 2369
rect 3099 2329 3111 2363
rect 3145 2360 3157 2363
rect 5905 2363 5963 2369
rect 3145 2332 5764 2360
rect 3145 2329 3157 2332
rect 3099 2323 3157 2329
rect 3510 2292 3516 2304
rect 3471 2264 3516 2292
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 4890 2292 4896 2304
rect 4851 2264 4896 2292
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 5736 2292 5764 2332
rect 5905 2329 5917 2363
rect 5951 2360 5963 2363
rect 10042 2360 10048 2372
rect 5951 2332 10048 2360
rect 5951 2329 5963 2332
rect 5905 2323 5963 2329
rect 10042 2320 10048 2332
rect 10100 2320 10106 2372
rect 16132 2369 16160 2468
rect 16206 2456 16212 2508
rect 16264 2496 16270 2508
rect 22572 2505 22600 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 23109 2527 23167 2533
rect 16644 2499 16702 2505
rect 16644 2496 16656 2499
rect 16264 2468 16656 2496
rect 16264 2456 16270 2468
rect 16644 2465 16656 2468
rect 16690 2496 16702 2499
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 16690 2468 17049 2496
rect 16690 2465 16702 2468
rect 16644 2459 16702 2465
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 18392 2499 18450 2505
rect 18392 2465 18404 2499
rect 18438 2465 18450 2499
rect 18392 2459 18450 2465
rect 20140 2499 20198 2505
rect 20140 2465 20152 2499
rect 20186 2465 20198 2499
rect 20140 2459 20198 2465
rect 22557 2499 22615 2505
rect 22557 2465 22569 2499
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 18407 2428 18435 2459
rect 18874 2428 18880 2440
rect 18407 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 20155 2428 20183 2459
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20155 2400 20637 2428
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 23198 2428 23204 2440
rect 20671 2400 23204 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 16117 2363 16175 2369
rect 16117 2329 16129 2363
rect 16163 2360 16175 2363
rect 16715 2363 16773 2369
rect 16715 2360 16727 2363
rect 16163 2332 16727 2360
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 16715 2329 16727 2332
rect 16761 2329 16773 2363
rect 16715 2323 16773 2329
rect 22741 2363 22799 2369
rect 22741 2329 22753 2363
rect 22787 2360 22799 2363
rect 24670 2360 24676 2372
rect 22787 2332 24676 2360
rect 22787 2329 22799 2332
rect 22741 2323 22799 2329
rect 24670 2320 24676 2332
rect 24728 2320 24734 2372
rect 9306 2292 9312 2304
rect 5736 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 9916 2264 10793 2292
rect 9916 2252 9922 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 14366 2292 14372 2304
rect 14327 2264 14372 2292
rect 10781 2255 10839 2261
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 26050 2292 26056 2304
rect 23256 2264 26056 2292
rect 23256 2252 23262 2264
rect 26050 2252 26056 2264
rect 26108 2252 26114 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 20254 2088 20260 2100
rect 14608 2060 20260 2088
rect 14608 2048 14614 2060
rect 20254 2048 20260 2060
rect 20312 2048 20318 2100
rect 14366 76 14372 128
rect 14424 116 14430 128
rect 23290 116 23296 128
rect 14424 88 23296 116
rect 14424 76 14430 88
rect 23290 76 23296 88
rect 23348 76 23354 128
<< via1 >>
rect 3056 27480 3108 27532
rect 3884 27480 3936 27532
rect 13912 27480 13964 27532
rect 14556 27480 14608 27532
rect 24860 27480 24912 27532
rect 25964 27480 26016 27532
rect 6920 26596 6972 26648
rect 8116 26596 8168 26648
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1860 24216 1912 24268
rect 6000 24216 6052 24268
rect 8760 24216 8812 24268
rect 2688 24012 2740 24064
rect 9220 24012 9272 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1860 23851 1912 23860
rect 1860 23817 1869 23851
rect 1869 23817 1903 23851
rect 1903 23817 1912 23851
rect 1860 23808 1912 23817
rect 8760 23851 8812 23860
rect 8760 23817 8769 23851
rect 8769 23817 8803 23851
rect 8803 23817 8812 23851
rect 8760 23808 8812 23817
rect 10692 23808 10744 23860
rect 15752 23808 15804 23860
rect 20904 23808 20956 23860
rect 23388 23808 23440 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 4344 23672 4396 23724
rect 1308 23604 1360 23656
rect 7196 23604 7248 23656
rect 9864 23647 9916 23656
rect 9864 23613 9873 23647
rect 9873 23613 9907 23647
rect 9907 23613 9916 23647
rect 9864 23604 9916 23613
rect 1400 23468 1452 23520
rect 7104 23468 7156 23520
rect 8668 23468 8720 23520
rect 17408 23604 17460 23656
rect 17500 23604 17552 23656
rect 19432 23536 19484 23588
rect 25136 23604 25188 23656
rect 15292 23468 15344 23520
rect 16488 23468 16540 23520
rect 17408 23511 17460 23520
rect 17408 23477 17417 23511
rect 17417 23477 17451 23511
rect 17451 23477 17460 23511
rect 17408 23468 17460 23477
rect 22928 23468 22980 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 9864 23264 9916 23316
rect 1584 23128 1636 23180
rect 10140 23128 10192 23180
rect 3792 22924 3844 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 9404 22720 9456 22772
rect 11980 22720 12032 22772
rect 24768 22763 24820 22772
rect 24768 22729 24777 22763
rect 24777 22729 24811 22763
rect 24811 22729 24820 22763
rect 24768 22720 24820 22729
rect 23664 22516 23716 22568
rect 9496 22423 9548 22432
rect 9496 22389 9505 22423
rect 9505 22389 9539 22423
rect 9539 22389 9548 22423
rect 9496 22380 9548 22389
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 10140 22380 10192 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 9496 22176 9548 22228
rect 8760 22040 8812 22092
rect 9864 22083 9916 22092
rect 9864 22049 9873 22083
rect 9873 22049 9907 22083
rect 9907 22049 9916 22083
rect 9864 22040 9916 22049
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 7840 21836 7892 21888
rect 9956 21879 10008 21888
rect 9956 21845 9965 21879
rect 9965 21845 9999 21879
rect 9999 21845 10008 21879
rect 9956 21836 10008 21845
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 9772 21632 9824 21684
rect 8760 21539 8812 21548
rect 8760 21505 8769 21539
rect 8769 21505 8803 21539
rect 8803 21505 8812 21539
rect 8760 21496 8812 21505
rect 10692 21496 10744 21548
rect 10876 21539 10928 21548
rect 10876 21505 10885 21539
rect 10885 21505 10919 21539
rect 10919 21505 10928 21539
rect 10876 21496 10928 21505
rect 8300 21471 8352 21480
rect 8300 21437 8309 21471
rect 8309 21437 8343 21471
rect 8343 21437 8352 21471
rect 8300 21428 8352 21437
rect 8208 21292 8260 21344
rect 8852 21292 8904 21344
rect 9680 21360 9732 21412
rect 11704 21360 11756 21412
rect 9772 21335 9824 21344
rect 9772 21301 9781 21335
rect 9781 21301 9815 21335
rect 9815 21301 9824 21335
rect 9772 21292 9824 21301
rect 10692 21292 10744 21344
rect 11244 21292 11296 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 10048 21131 10100 21140
rect 10048 21097 10057 21131
rect 10057 21097 10091 21131
rect 10091 21097 10100 21131
rect 10048 21088 10100 21097
rect 7840 21063 7892 21072
rect 7840 21029 7849 21063
rect 7849 21029 7883 21063
rect 7883 21029 7892 21063
rect 7840 21020 7892 21029
rect 7932 21063 7984 21072
rect 7932 21029 7941 21063
rect 7941 21029 7975 21063
rect 7975 21029 7984 21063
rect 10324 21063 10376 21072
rect 7932 21020 7984 21029
rect 10324 21029 10333 21063
rect 10333 21029 10367 21063
rect 10367 21029 10376 21063
rect 10324 21020 10376 21029
rect 10876 21063 10928 21072
rect 10876 21029 10885 21063
rect 10885 21029 10919 21063
rect 10919 21029 10928 21063
rect 10876 21020 10928 21029
rect 1952 20952 2004 21004
rect 6644 20952 6696 21004
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 22836 20995 22888 21004
rect 22836 20961 22854 20995
rect 22854 20961 22888 20995
rect 22836 20952 22888 20961
rect 24676 20952 24728 21004
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 10324 20884 10376 20936
rect 11060 20884 11112 20936
rect 6828 20748 6880 20800
rect 8760 20791 8812 20800
rect 8760 20757 8769 20791
rect 8769 20757 8803 20791
rect 8803 20757 8812 20791
rect 8760 20748 8812 20757
rect 18328 20748 18380 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 9956 20544 10008 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 8760 20408 8812 20460
rect 10048 20451 10100 20460
rect 10048 20417 10057 20451
rect 10057 20417 10091 20451
rect 10091 20417 10100 20451
rect 10048 20408 10100 20417
rect 10232 20408 10284 20460
rect 14280 20544 14332 20596
rect 17500 20544 17552 20596
rect 22836 20587 22888 20596
rect 22836 20553 22845 20587
rect 22845 20553 22879 20587
rect 22879 20553 22888 20587
rect 22836 20544 22888 20553
rect 8208 20315 8260 20324
rect 8208 20281 8217 20315
rect 8217 20281 8251 20315
rect 8251 20281 8260 20315
rect 8208 20272 8260 20281
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 10692 20315 10744 20324
rect 1952 20204 2004 20256
rect 3700 20204 3752 20256
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 6000 20204 6052 20256
rect 6276 20247 6328 20256
rect 6276 20213 6285 20247
rect 6285 20213 6319 20247
rect 6319 20213 6328 20247
rect 6276 20204 6328 20213
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 7196 20204 7248 20256
rect 7932 20204 7984 20256
rect 9956 20204 10008 20256
rect 10692 20281 10701 20315
rect 10701 20281 10735 20315
rect 10735 20281 10744 20315
rect 10692 20272 10744 20281
rect 13084 20204 13136 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 11704 20000 11756 20052
rect 7196 19975 7248 19984
rect 7196 19941 7205 19975
rect 7205 19941 7239 19975
rect 7239 19941 7248 19975
rect 7196 19932 7248 19941
rect 8116 19975 8168 19984
rect 8116 19941 8125 19975
rect 8125 19941 8159 19975
rect 8159 19941 8168 19975
rect 8116 19932 8168 19941
rect 8208 19975 8260 19984
rect 8208 19941 8217 19975
rect 8217 19941 8251 19975
rect 8251 19941 8260 19975
rect 8760 19975 8812 19984
rect 8208 19932 8260 19941
rect 8760 19941 8769 19975
rect 8769 19941 8803 19975
rect 8803 19941 8812 19975
rect 8760 19932 8812 19941
rect 9772 19932 9824 19984
rect 10692 19932 10744 19984
rect 11612 19975 11664 19984
rect 11612 19941 11621 19975
rect 11621 19941 11655 19975
rect 11655 19941 11664 19975
rect 11612 19932 11664 19941
rect 13084 19975 13136 19984
rect 13084 19941 13093 19975
rect 13093 19941 13127 19975
rect 13127 19941 13136 19975
rect 13084 19932 13136 19941
rect 13268 19932 13320 19984
rect 4988 19907 5040 19916
rect 4988 19873 4997 19907
rect 4997 19873 5031 19907
rect 5031 19873 5040 19907
rect 4988 19864 5040 19873
rect 6552 19907 6604 19916
rect 6552 19873 6561 19907
rect 6561 19873 6595 19907
rect 6595 19873 6604 19907
rect 6552 19864 6604 19873
rect 3976 19796 4028 19848
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 11428 19728 11480 19780
rect 11704 19796 11756 19848
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 13728 19660 13780 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 4068 19456 4120 19508
rect 4988 19499 5040 19508
rect 4988 19465 4997 19499
rect 4997 19465 5031 19499
rect 5031 19465 5040 19499
rect 4988 19456 5040 19465
rect 6552 19499 6604 19508
rect 6552 19465 6561 19499
rect 6561 19465 6595 19499
rect 6595 19465 6604 19499
rect 6552 19456 6604 19465
rect 7748 19456 7800 19508
rect 10140 19499 10192 19508
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 7196 19388 7248 19440
rect 9496 19388 9548 19440
rect 4344 19363 4396 19372
rect 4344 19329 4353 19363
rect 4353 19329 4387 19363
rect 4387 19329 4396 19363
rect 4344 19320 4396 19329
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 9956 19320 10008 19372
rect 13360 19320 13412 19372
rect 1124 19252 1176 19304
rect 5264 19252 5316 19304
rect 2044 19116 2096 19168
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 4160 19227 4212 19236
rect 4160 19193 4169 19227
rect 4169 19193 4203 19227
rect 4203 19193 4212 19227
rect 4160 19184 4212 19193
rect 8576 19252 8628 19304
rect 7656 19227 7708 19236
rect 7656 19193 7665 19227
rect 7665 19193 7699 19227
rect 7699 19193 7708 19227
rect 7656 19184 7708 19193
rect 7748 19227 7800 19236
rect 7748 19193 7757 19227
rect 7757 19193 7791 19227
rect 7791 19193 7800 19227
rect 7748 19184 7800 19193
rect 9956 19184 10008 19236
rect 3424 19116 3476 19125
rect 6736 19116 6788 19168
rect 7840 19116 7892 19168
rect 8208 19116 8260 19168
rect 9128 19116 9180 19168
rect 10140 19116 10192 19168
rect 10876 19116 10928 19168
rect 11612 19184 11664 19236
rect 11428 19159 11480 19168
rect 11428 19125 11437 19159
rect 11437 19125 11471 19159
rect 11471 19125 11480 19159
rect 11428 19116 11480 19125
rect 12256 19116 12308 19168
rect 13360 19116 13412 19168
rect 14004 19184 14056 19236
rect 14372 19227 14424 19236
rect 14372 19193 14381 19227
rect 14381 19193 14415 19227
rect 14415 19193 14424 19227
rect 14372 19184 14424 19193
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 3424 18912 3476 18964
rect 6920 18912 6972 18964
rect 5080 18887 5132 18896
rect 5080 18853 5089 18887
rect 5089 18853 5123 18887
rect 5123 18853 5132 18887
rect 5080 18844 5132 18853
rect 7104 18887 7156 18896
rect 7104 18853 7107 18887
rect 7107 18853 7141 18887
rect 7141 18853 7156 18887
rect 7104 18844 7156 18853
rect 7748 18912 7800 18964
rect 8116 18912 8168 18964
rect 13084 18955 13136 18964
rect 13084 18921 13093 18955
rect 13093 18921 13127 18955
rect 13127 18921 13136 18955
rect 13084 18912 13136 18921
rect 13728 18912 13780 18964
rect 14004 18912 14056 18964
rect 9496 18844 9548 18896
rect 10876 18887 10928 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 8484 18819 8536 18828
rect 8484 18785 8493 18819
rect 8493 18785 8527 18819
rect 8527 18785 8536 18819
rect 8484 18776 8536 18785
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 13820 18887 13872 18896
rect 13820 18853 13829 18887
rect 13829 18853 13863 18887
rect 13863 18853 13872 18887
rect 14372 18887 14424 18896
rect 13820 18844 13872 18853
rect 14372 18853 14381 18887
rect 14381 18853 14415 18887
rect 14415 18853 14424 18887
rect 16488 18887 16540 18896
rect 14372 18844 14424 18853
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 15476 18776 15528 18828
rect 2964 18751 3016 18760
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 2964 18708 3016 18717
rect 5356 18708 5408 18760
rect 6920 18708 6972 18760
rect 11152 18708 11204 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 13452 18708 13504 18760
rect 5540 18683 5592 18692
rect 5540 18649 5549 18683
rect 5549 18649 5583 18683
rect 5583 18649 5592 18683
rect 5540 18640 5592 18649
rect 9312 18640 9364 18692
rect 9956 18640 10008 18692
rect 16028 18708 16080 18760
rect 16488 18853 16497 18887
rect 16497 18853 16531 18887
rect 16531 18853 16540 18887
rect 16488 18844 16540 18853
rect 16580 18887 16632 18896
rect 16580 18853 16589 18887
rect 16589 18853 16623 18887
rect 16623 18853 16632 18887
rect 16580 18844 16632 18853
rect 17684 18708 17736 18760
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 7932 18572 7984 18581
rect 8208 18572 8260 18624
rect 8760 18572 8812 18624
rect 9772 18572 9824 18624
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13728 18572 13780 18624
rect 14648 18572 14700 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1400 18368 1452 18420
rect 4804 18368 4856 18420
rect 2964 18232 3016 18284
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 4344 18232 4396 18284
rect 3976 18096 4028 18148
rect 5080 18368 5132 18420
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 7656 18368 7708 18420
rect 9680 18368 9732 18420
rect 11796 18368 11848 18420
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 12624 18368 12676 18420
rect 14832 18368 14884 18420
rect 15476 18411 15528 18420
rect 15476 18377 15485 18411
rect 15485 18377 15519 18411
rect 15519 18377 15528 18411
rect 15476 18368 15528 18377
rect 19432 18368 19484 18420
rect 25136 18411 25188 18420
rect 25136 18377 25145 18411
rect 25145 18377 25179 18411
rect 25179 18377 25188 18411
rect 25136 18368 25188 18377
rect 8484 18300 8536 18352
rect 8852 18300 8904 18352
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 6276 18232 6328 18284
rect 9220 18232 9272 18284
rect 5724 18164 5776 18216
rect 112 18028 164 18080
rect 4160 18028 4212 18080
rect 5264 18096 5316 18148
rect 7932 18164 7984 18216
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 13636 18300 13688 18352
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 11796 18164 11848 18216
rect 25136 18164 25188 18216
rect 7104 18028 7156 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 10692 18096 10744 18148
rect 14464 18139 14516 18148
rect 14464 18105 14473 18139
rect 14473 18105 14507 18139
rect 14507 18105 14516 18139
rect 14464 18096 14516 18105
rect 14556 18139 14608 18148
rect 14556 18105 14565 18139
rect 14565 18105 14599 18139
rect 14599 18105 14608 18139
rect 14556 18096 14608 18105
rect 7748 18028 7800 18037
rect 10784 18028 10836 18080
rect 10876 18028 10928 18080
rect 11060 18028 11112 18080
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 13544 18028 13596 18080
rect 13820 18028 13872 18080
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 15752 18028 15804 18037
rect 16580 18028 16632 18080
rect 18604 18028 18656 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 2044 17867 2096 17876
rect 2044 17833 2053 17867
rect 2053 17833 2087 17867
rect 2087 17833 2096 17867
rect 2044 17824 2096 17833
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 7840 17867 7892 17876
rect 7840 17833 7849 17867
rect 7849 17833 7883 17867
rect 7883 17833 7892 17867
rect 7840 17824 7892 17833
rect 9220 17824 9272 17876
rect 11060 17824 11112 17876
rect 11152 17867 11204 17876
rect 11152 17833 11161 17867
rect 11161 17833 11195 17867
rect 11195 17833 11204 17867
rect 11152 17824 11204 17833
rect 13544 17867 13596 17876
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 4712 17799 4764 17808
rect 4712 17765 4721 17799
rect 4721 17765 4755 17799
rect 4755 17765 4764 17799
rect 4712 17756 4764 17765
rect 7104 17756 7156 17808
rect 7748 17756 7800 17808
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 10784 17756 10836 17808
rect 11796 17756 11848 17808
rect 13728 17799 13780 17808
rect 13728 17765 13737 17799
rect 13737 17765 13771 17799
rect 13771 17765 13780 17799
rect 13728 17756 13780 17765
rect 14004 17756 14056 17808
rect 14464 17756 14516 17808
rect 1584 17688 1636 17740
rect 2504 17731 2556 17740
rect 2504 17697 2513 17731
rect 2513 17697 2547 17731
rect 2547 17697 2556 17731
rect 2504 17688 2556 17697
rect 5356 17688 5408 17740
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 15568 17688 15620 17740
rect 3424 17620 3476 17672
rect 3056 17552 3108 17604
rect 6184 17620 6236 17672
rect 8668 17620 8720 17672
rect 9588 17620 9640 17672
rect 10692 17620 10744 17672
rect 11244 17620 11296 17672
rect 12256 17620 12308 17672
rect 5172 17552 5224 17604
rect 11980 17595 12032 17604
rect 11980 17561 11989 17595
rect 11989 17561 12023 17595
rect 12023 17561 12032 17595
rect 11980 17552 12032 17561
rect 13636 17552 13688 17604
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 2320 17527 2372 17536
rect 2320 17493 2329 17527
rect 2329 17493 2363 17527
rect 2363 17493 2372 17527
rect 2320 17484 2372 17493
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 6920 17484 6972 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 4712 17280 4764 17332
rect 8760 17323 8812 17332
rect 8760 17289 8769 17323
rect 8769 17289 8803 17323
rect 8803 17289 8812 17323
rect 8760 17280 8812 17289
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 9864 17280 9916 17332
rect 5540 17212 5592 17264
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 2044 17076 2096 17128
rect 8116 17144 8168 17196
rect 8760 17144 8812 17196
rect 5356 17008 5408 17060
rect 6368 17008 6420 17060
rect 7748 17051 7800 17060
rect 7748 17017 7757 17051
rect 7757 17017 7791 17051
rect 7791 17017 7800 17051
rect 7748 17008 7800 17017
rect 8668 17008 8720 17060
rect 11060 17144 11112 17196
rect 11980 17144 12032 17196
rect 14556 17280 14608 17332
rect 14004 17212 14056 17264
rect 14372 17212 14424 17264
rect 24768 17255 24820 17264
rect 24768 17221 24777 17255
rect 24777 17221 24811 17255
rect 24811 17221 24820 17255
rect 24768 17212 24820 17221
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 13176 17076 13228 17128
rect 10692 17008 10744 17060
rect 12256 17051 12308 17060
rect 12256 17017 12265 17051
rect 12265 17017 12299 17051
rect 12299 17017 12308 17051
rect 12256 17008 12308 17017
rect 13636 17008 13688 17060
rect 112 16940 164 16992
rect 1676 16940 1728 16992
rect 2044 16940 2096 16992
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 7104 16940 7156 16992
rect 11428 16940 11480 16992
rect 11796 16983 11848 16992
rect 11796 16949 11805 16983
rect 11805 16949 11839 16983
rect 11839 16949 11848 16983
rect 11796 16940 11848 16949
rect 12900 16940 12952 16992
rect 13360 16983 13412 16992
rect 13360 16949 13369 16983
rect 13369 16949 13403 16983
rect 13403 16949 13412 16983
rect 14004 17076 14056 17128
rect 15292 17076 15344 17128
rect 24216 17076 24268 17128
rect 16396 17051 16448 17060
rect 16396 17017 16405 17051
rect 16405 17017 16439 17051
rect 16439 17017 16448 17051
rect 16948 17051 17000 17060
rect 16396 17008 16448 17017
rect 16948 17017 16957 17051
rect 16957 17017 16991 17051
rect 16991 17017 17000 17051
rect 16948 17008 17000 17017
rect 15384 16983 15436 16992
rect 13360 16940 13412 16949
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 15568 16940 15620 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1768 16736 1820 16788
rect 2320 16736 2372 16788
rect 5264 16736 5316 16788
rect 5540 16736 5592 16788
rect 9956 16736 10008 16788
rect 11796 16736 11848 16788
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 4804 16711 4856 16720
rect 4804 16677 4807 16711
rect 4807 16677 4841 16711
rect 4841 16677 4856 16711
rect 4804 16668 4856 16677
rect 6368 16668 6420 16720
rect 9404 16668 9456 16720
rect 12256 16711 12308 16720
rect 1860 16600 1912 16652
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 2872 16600 2924 16652
rect 6092 16600 6144 16652
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 8300 16643 8352 16652
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 5540 16532 5592 16584
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 12256 16677 12265 16711
rect 12265 16677 12299 16711
rect 12299 16677 12308 16711
rect 12256 16668 12308 16677
rect 12900 16668 12952 16720
rect 13728 16711 13780 16720
rect 13728 16677 13737 16711
rect 13737 16677 13771 16711
rect 13771 16677 13780 16711
rect 13728 16668 13780 16677
rect 14188 16668 14240 16720
rect 7656 16532 7708 16584
rect 9496 16532 9548 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 14740 16668 14792 16720
rect 15660 16668 15712 16720
rect 17776 16711 17828 16720
rect 17776 16677 17785 16711
rect 17785 16677 17819 16711
rect 17819 16677 17828 16711
rect 17776 16668 17828 16677
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 24124 16600 24176 16652
rect 16304 16532 16356 16584
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 4436 16396 4488 16448
rect 8116 16396 8168 16448
rect 10784 16396 10836 16448
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 14188 16396 14240 16448
rect 15752 16396 15804 16448
rect 16948 16396 17000 16448
rect 18512 16396 18564 16448
rect 27620 16396 27672 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 3884 16192 3936 16201
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 6092 16235 6144 16244
rect 6092 16201 6101 16235
rect 6101 16201 6135 16235
rect 6135 16201 6144 16235
rect 6092 16192 6144 16201
rect 10692 16192 10744 16244
rect 12164 16192 12216 16244
rect 13728 16192 13780 16244
rect 15936 16192 15988 16244
rect 17776 16192 17828 16244
rect 24124 16192 24176 16244
rect 4620 16124 4672 16176
rect 9956 16124 10008 16176
rect 13360 16124 13412 16176
rect 18052 16124 18104 16176
rect 3148 16056 3200 16108
rect 9036 16056 9088 16108
rect 2320 15988 2372 16040
rect 3332 15988 3384 16040
rect 3884 15988 3936 16040
rect 4436 16031 4488 16040
rect 4436 15997 4445 16031
rect 4445 15997 4479 16031
rect 4479 15997 4488 16031
rect 4436 15988 4488 15997
rect 7656 16031 7708 16040
rect 5080 15920 5132 15972
rect 6460 15963 6512 15972
rect 6460 15929 6469 15963
rect 6469 15929 6503 15963
rect 6503 15929 6512 15963
rect 6460 15920 6512 15929
rect 7656 15997 7665 16031
rect 7665 15997 7699 16031
rect 7699 15997 7708 16031
rect 7656 15988 7708 15997
rect 10968 16056 11020 16108
rect 11704 16056 11756 16108
rect 12256 16056 12308 16108
rect 13452 16099 13504 16108
rect 12348 15988 12400 16040
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 13636 16056 13688 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 14372 16031 14424 16040
rect 8944 15920 8996 15972
rect 10784 15963 10836 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 5540 15852 5592 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 10784 15929 10793 15963
rect 10793 15929 10827 15963
rect 10827 15929 10836 15963
rect 10784 15920 10836 15929
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 15108 15988 15160 16040
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 9956 15895 10008 15904
rect 8668 15852 8720 15861
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10692 15852 10744 15904
rect 13360 15920 13412 15972
rect 14096 15920 14148 15972
rect 14188 15920 14240 15972
rect 14740 15920 14792 15972
rect 16304 15963 16356 15972
rect 16304 15929 16313 15963
rect 16313 15929 16347 15963
rect 16347 15929 16356 15963
rect 16304 15920 16356 15929
rect 15660 15852 15712 15904
rect 18788 15920 18840 15972
rect 16580 15852 16632 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 4436 15648 4488 15700
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 9036 15691 9088 15700
rect 9036 15657 9045 15691
rect 9045 15657 9079 15691
rect 9079 15657 9088 15691
rect 9036 15648 9088 15657
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 9956 15648 10008 15700
rect 1676 15623 1728 15632
rect 1676 15589 1685 15623
rect 1685 15589 1719 15623
rect 1719 15589 1728 15623
rect 1676 15580 1728 15589
rect 2412 15580 2464 15632
rect 3792 15580 3844 15632
rect 4804 15580 4856 15632
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 4620 15512 4672 15521
rect 5172 15512 5224 15564
rect 7656 15580 7708 15632
rect 5356 15512 5408 15564
rect 3424 15444 3476 15496
rect 4988 15376 5040 15428
rect 6828 15512 6880 15564
rect 7380 15555 7432 15564
rect 7380 15521 7389 15555
rect 7389 15521 7423 15555
rect 7423 15521 7432 15555
rect 7380 15512 7432 15521
rect 7564 15512 7616 15564
rect 9128 15580 9180 15632
rect 10968 15648 11020 15700
rect 11796 15580 11848 15632
rect 8944 15512 8996 15564
rect 9864 15512 9916 15564
rect 13176 15648 13228 15700
rect 15844 15691 15896 15700
rect 15844 15657 15853 15691
rect 15853 15657 15887 15691
rect 15887 15657 15896 15691
rect 15844 15648 15896 15657
rect 17776 15648 17828 15700
rect 18052 15691 18104 15700
rect 18052 15657 18061 15691
rect 18061 15657 18095 15691
rect 18095 15657 18104 15691
rect 18052 15648 18104 15657
rect 15660 15580 15712 15632
rect 17684 15623 17736 15632
rect 17684 15589 17693 15623
rect 17693 15589 17727 15623
rect 17727 15589 17736 15623
rect 17684 15580 17736 15589
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 17960 15512 18012 15521
rect 7104 15444 7156 15496
rect 11612 15444 11664 15496
rect 10140 15376 10192 15428
rect 11704 15376 11756 15428
rect 16856 15444 16908 15496
rect 17868 15444 17920 15496
rect 13452 15376 13504 15428
rect 2596 15351 2648 15360
rect 2596 15317 2605 15351
rect 2605 15317 2639 15351
rect 2639 15317 2648 15351
rect 2596 15308 2648 15317
rect 2688 15308 2740 15360
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1492 15104 1544 15156
rect 1676 15104 1728 15156
rect 4620 15104 4672 15156
rect 10784 15104 10836 15156
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 13268 15104 13320 15156
rect 14096 15104 14148 15156
rect 15660 15104 15712 15156
rect 16396 15104 16448 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 17960 15104 18012 15156
rect 22100 15104 22152 15156
rect 3148 15079 3200 15088
rect 3148 15045 3157 15079
rect 3157 15045 3191 15079
rect 3191 15045 3200 15079
rect 3148 15036 3200 15045
rect 5540 15036 5592 15088
rect 7932 15036 7984 15088
rect 9956 15036 10008 15088
rect 11888 15036 11940 15088
rect 2412 14968 2464 15020
rect 8024 14968 8076 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 4620 14943 4672 14952
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 4620 14900 4672 14909
rect 5172 14943 5224 14952
rect 5172 14909 5181 14943
rect 5181 14909 5215 14943
rect 5215 14909 5224 14943
rect 5172 14900 5224 14909
rect 5264 14943 5316 14952
rect 5264 14909 5273 14943
rect 5273 14909 5307 14943
rect 5307 14909 5316 14943
rect 5816 14943 5868 14952
rect 5264 14900 5316 14909
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7380 14943 7432 14952
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 7564 14900 7616 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 12348 14968 12400 15020
rect 12716 14968 12768 15020
rect 13728 14968 13780 15020
rect 2688 14875 2740 14884
rect 2688 14841 2697 14875
rect 2697 14841 2731 14875
rect 2731 14841 2740 14875
rect 2688 14832 2740 14841
rect 4344 14832 4396 14884
rect 7472 14832 7524 14884
rect 10140 14900 10192 14952
rect 15568 14968 15620 15020
rect 2320 14807 2372 14816
rect 2320 14773 2329 14807
rect 2329 14773 2363 14807
rect 2363 14773 2372 14807
rect 2320 14764 2372 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4804 14764 4856 14816
rect 7564 14764 7616 14816
rect 9956 14764 10008 14816
rect 10876 14832 10928 14884
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 13636 14764 13688 14816
rect 15936 14968 15988 15020
rect 16488 14900 16540 14952
rect 19432 14968 19484 15020
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 15752 14832 15804 14884
rect 17868 14832 17920 14884
rect 18144 14807 18196 14816
rect 18144 14773 18153 14807
rect 18153 14773 18187 14807
rect 18187 14773 18196 14807
rect 18144 14764 18196 14773
rect 20904 14764 20956 14816
rect 21364 14764 21416 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 7656 14560 7708 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 9956 14560 10008 14612
rect 2780 14492 2832 14544
rect 3148 14535 3200 14544
rect 3148 14501 3157 14535
rect 3157 14501 3191 14535
rect 3191 14501 3200 14535
rect 3148 14492 3200 14501
rect 6000 14492 6052 14544
rect 11336 14560 11388 14612
rect 8208 14492 8260 14544
rect 4620 14424 4672 14476
rect 6092 14424 6144 14476
rect 6828 14467 6880 14476
rect 6828 14433 6837 14467
rect 6837 14433 6871 14467
rect 6871 14433 6880 14467
rect 6828 14424 6880 14433
rect 7104 14424 7156 14476
rect 10140 14492 10192 14544
rect 10232 14492 10284 14544
rect 11612 14535 11664 14544
rect 11612 14501 11621 14535
rect 11621 14501 11655 14535
rect 11655 14501 11664 14535
rect 11612 14492 11664 14501
rect 11980 14535 12032 14544
rect 11980 14501 11989 14535
rect 11989 14501 12023 14535
rect 12023 14501 12032 14535
rect 11980 14492 12032 14501
rect 13452 14535 13504 14544
rect 13452 14501 13461 14535
rect 13461 14501 13495 14535
rect 13495 14501 13504 14535
rect 13452 14492 13504 14501
rect 13820 14492 13872 14544
rect 17592 14560 17644 14612
rect 19340 14560 19392 14612
rect 20260 14560 20312 14612
rect 15752 14492 15804 14544
rect 16856 14535 16908 14544
rect 16856 14501 16865 14535
rect 16865 14501 16899 14535
rect 16899 14501 16908 14535
rect 16856 14492 16908 14501
rect 18512 14492 18564 14544
rect 16580 14467 16632 14476
rect 5448 14356 5500 14408
rect 6736 14356 6788 14408
rect 16580 14433 16589 14467
rect 16589 14433 16623 14467
rect 16623 14433 16632 14467
rect 16580 14424 16632 14433
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 8668 14356 8720 14408
rect 9772 14356 9824 14408
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 3608 14288 3660 14340
rect 5264 14288 5316 14340
rect 5816 14288 5868 14340
rect 6368 14288 6420 14340
rect 8116 14288 8168 14340
rect 11704 14288 11756 14340
rect 13636 14288 13688 14340
rect 19800 14424 19852 14476
rect 21088 14467 21140 14476
rect 21088 14433 21097 14467
rect 21097 14433 21131 14467
rect 21131 14433 21140 14467
rect 21088 14424 21140 14433
rect 21824 14356 21876 14408
rect 19340 14288 19392 14340
rect 2228 14220 2280 14272
rect 3700 14220 3752 14272
rect 4160 14220 4212 14272
rect 6552 14263 6604 14272
rect 6552 14229 6561 14263
rect 6561 14229 6595 14263
rect 6595 14229 6604 14263
rect 6552 14220 6604 14229
rect 11152 14220 11204 14272
rect 12624 14220 12676 14272
rect 13728 14220 13780 14272
rect 16120 14220 16172 14272
rect 18512 14220 18564 14272
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 20076 14220 20128 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 7104 14016 7156 14068
rect 11980 14016 12032 14068
rect 13820 14016 13872 14068
rect 15568 14016 15620 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 19800 14059 19852 14068
rect 19800 14025 19809 14059
rect 19809 14025 19843 14059
rect 19843 14025 19852 14059
rect 19800 14016 19852 14025
rect 19984 14016 20036 14068
rect 21088 14016 21140 14068
rect 25136 14059 25188 14068
rect 25136 14025 25145 14059
rect 25145 14025 25179 14059
rect 25179 14025 25188 14059
rect 25136 14016 25188 14025
rect 3148 13948 3200 14000
rect 3884 13948 3936 14000
rect 4160 13948 4212 14000
rect 2596 13880 2648 13932
rect 3516 13880 3568 13932
rect 3884 13855 3936 13864
rect 1952 13744 2004 13796
rect 2136 13676 2188 13728
rect 2320 13676 2372 13728
rect 2780 13719 2832 13728
rect 2780 13685 2789 13719
rect 2789 13685 2823 13719
rect 2823 13685 2832 13719
rect 2780 13676 2832 13685
rect 3516 13719 3568 13728
rect 3516 13685 3525 13719
rect 3525 13685 3559 13719
rect 3559 13685 3568 13719
rect 3516 13676 3568 13685
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 4252 13855 4304 13864
rect 4252 13821 4261 13855
rect 4261 13821 4295 13855
rect 4295 13821 4304 13855
rect 4252 13812 4304 13821
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 9128 13880 9180 13932
rect 9496 13880 9548 13932
rect 10692 13880 10744 13932
rect 11888 13880 11940 13932
rect 13176 13880 13228 13932
rect 15660 13991 15712 14000
rect 15660 13957 15669 13991
rect 15669 13957 15703 13991
rect 15703 13957 15712 13991
rect 15660 13948 15712 13957
rect 6368 13812 6420 13864
rect 6736 13812 6788 13864
rect 6092 13744 6144 13796
rect 6552 13744 6604 13796
rect 5264 13676 5316 13728
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 7196 13676 7248 13728
rect 7932 13812 7984 13864
rect 8852 13812 8904 13864
rect 9036 13744 9088 13796
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 12808 13744 12860 13796
rect 11612 13676 11664 13728
rect 13728 13744 13780 13796
rect 15936 13812 15988 13864
rect 16856 13880 16908 13932
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 21364 13880 21416 13932
rect 16488 13855 16540 13864
rect 16488 13821 16497 13855
rect 16497 13821 16531 13855
rect 16531 13821 16540 13855
rect 16488 13812 16540 13821
rect 17868 13812 17920 13864
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 25136 13812 25188 13864
rect 18512 13787 18564 13796
rect 18512 13753 18521 13787
rect 18521 13753 18555 13787
rect 18555 13753 18564 13787
rect 18512 13744 18564 13753
rect 21272 13787 21324 13796
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 21272 13753 21281 13787
rect 21281 13753 21315 13787
rect 21315 13753 21324 13787
rect 21272 13744 21324 13753
rect 22008 13744 22060 13796
rect 18236 13676 18288 13685
rect 19340 13676 19392 13728
rect 21180 13676 21232 13728
rect 21732 13676 21784 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2688 13472 2740 13524
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 5448 13472 5500 13524
rect 6184 13515 6236 13524
rect 1952 13404 2004 13456
rect 2780 13404 2832 13456
rect 2044 13336 2096 13388
rect 2320 13336 2372 13388
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 8208 13515 8260 13524
rect 8208 13481 8217 13515
rect 8217 13481 8251 13515
rect 8251 13481 8260 13515
rect 8208 13472 8260 13481
rect 7564 13404 7616 13456
rect 9036 13472 9088 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13452 13472 13504 13524
rect 16488 13472 16540 13524
rect 18236 13472 18288 13524
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 11152 13447 11204 13456
rect 11152 13413 11161 13447
rect 11161 13413 11195 13447
rect 11195 13413 11204 13447
rect 11152 13404 11204 13413
rect 11796 13404 11848 13456
rect 13176 13447 13228 13456
rect 13176 13413 13185 13447
rect 13185 13413 13219 13447
rect 13219 13413 13228 13447
rect 13176 13404 13228 13413
rect 13728 13447 13780 13456
rect 13728 13413 13737 13447
rect 13737 13413 13771 13447
rect 13771 13413 13780 13447
rect 13728 13404 13780 13413
rect 17316 13404 17368 13456
rect 19156 13447 19208 13456
rect 19156 13413 19165 13447
rect 19165 13413 19199 13447
rect 19199 13413 19208 13447
rect 19156 13404 19208 13413
rect 21088 13472 21140 13524
rect 21364 13472 21416 13524
rect 21548 13404 21600 13456
rect 21824 13447 21876 13456
rect 21824 13413 21833 13447
rect 21833 13413 21867 13447
rect 21867 13413 21876 13447
rect 21824 13404 21876 13413
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 7196 13336 7248 13388
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 9496 13336 9548 13388
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 15568 13336 15620 13345
rect 15844 13336 15896 13388
rect 16120 13336 16172 13388
rect 22376 13336 22428 13388
rect 23388 13336 23440 13388
rect 3240 13268 3292 13320
rect 3700 13268 3752 13320
rect 11244 13268 11296 13320
rect 11520 13268 11572 13320
rect 13084 13311 13136 13320
rect 13084 13277 13093 13311
rect 13093 13277 13127 13311
rect 13127 13277 13136 13311
rect 13084 13268 13136 13277
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 18144 13268 18196 13320
rect 19524 13268 19576 13320
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 1952 13200 2004 13252
rect 9956 13200 10008 13252
rect 11704 13200 11756 13252
rect 2044 13175 2096 13184
rect 2044 13141 2053 13175
rect 2053 13141 2087 13175
rect 2087 13141 2096 13175
rect 2044 13132 2096 13141
rect 5172 13175 5224 13184
rect 5172 13141 5181 13175
rect 5181 13141 5215 13175
rect 5215 13141 5224 13175
rect 5172 13132 5224 13141
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 11428 13132 11480 13184
rect 19432 13132 19484 13184
rect 24216 13132 24268 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 11612 12928 11664 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 13176 12928 13228 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 16396 12928 16448 12980
rect 18144 12928 18196 12980
rect 21824 12928 21876 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 1768 12792 1820 12844
rect 2412 12792 2464 12844
rect 3516 12792 3568 12844
rect 4436 12860 4488 12912
rect 9496 12792 9548 12844
rect 15660 12860 15712 12912
rect 13728 12792 13780 12844
rect 3148 12724 3200 12776
rect 3424 12724 3476 12776
rect 4252 12767 4304 12776
rect 4252 12733 4261 12767
rect 4261 12733 4295 12767
rect 4295 12733 4304 12767
rect 4252 12724 4304 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4988 12767 5040 12776
rect 4436 12724 4488 12733
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 7104 12724 7156 12776
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 8944 12724 8996 12776
rect 12164 12724 12216 12776
rect 15844 12724 15896 12776
rect 2136 12656 2188 12708
rect 5172 12656 5224 12708
rect 7380 12656 7432 12708
rect 1952 12588 2004 12640
rect 3148 12588 3200 12640
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 5264 12588 5316 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 8668 12588 8720 12640
rect 9772 12588 9824 12640
rect 10140 12588 10192 12640
rect 12900 12656 12952 12708
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 14372 12656 14424 12708
rect 19892 12860 19944 12912
rect 16212 12835 16264 12844
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 17592 12792 17644 12844
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 20076 12835 20128 12844
rect 18880 12792 18932 12801
rect 20076 12801 20085 12835
rect 20085 12801 20119 12835
rect 20119 12801 20128 12835
rect 20076 12792 20128 12801
rect 21548 12792 21600 12844
rect 23756 12767 23808 12776
rect 23756 12733 23774 12767
rect 23774 12733 23808 12767
rect 23756 12724 23808 12733
rect 16764 12656 16816 12708
rect 17316 12656 17368 12708
rect 18236 12699 18288 12708
rect 18236 12665 18245 12699
rect 18245 12665 18279 12699
rect 18279 12665 18288 12699
rect 18236 12656 18288 12665
rect 18328 12699 18380 12708
rect 18328 12665 18337 12699
rect 18337 12665 18371 12699
rect 18371 12665 18380 12699
rect 18328 12656 18380 12665
rect 19432 12656 19484 12708
rect 19892 12699 19944 12708
rect 19892 12665 19901 12699
rect 19901 12665 19935 12699
rect 19935 12665 19944 12699
rect 19892 12656 19944 12665
rect 20076 12656 20128 12708
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 19156 12631 19208 12640
rect 19156 12597 19165 12631
rect 19165 12597 19199 12631
rect 19199 12597 19208 12631
rect 19156 12588 19208 12597
rect 19524 12631 19576 12640
rect 19524 12597 19533 12631
rect 19533 12597 19567 12631
rect 19567 12597 19576 12631
rect 19524 12588 19576 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 4252 12384 4304 12436
rect 7288 12384 7340 12436
rect 8852 12384 8904 12436
rect 9956 12384 10008 12436
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 16212 12427 16264 12436
rect 16212 12393 16221 12427
rect 16221 12393 16255 12427
rect 16255 12393 16264 12427
rect 16212 12384 16264 12393
rect 18328 12384 18380 12436
rect 19156 12384 19208 12436
rect 19984 12384 20036 12436
rect 21732 12427 21784 12436
rect 21732 12393 21741 12427
rect 21741 12393 21775 12427
rect 21775 12393 21784 12427
rect 21732 12384 21784 12393
rect 3884 12316 3936 12368
rect 4896 12316 4948 12368
rect 10324 12316 10376 12368
rect 1308 12248 1360 12300
rect 4436 12248 4488 12300
rect 5172 12248 5224 12300
rect 5540 12248 5592 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 7104 12248 7156 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 8576 12248 8628 12300
rect 8944 12248 8996 12300
rect 10140 12248 10192 12300
rect 13820 12359 13872 12368
rect 13820 12325 13829 12359
rect 13829 12325 13863 12359
rect 13863 12325 13872 12359
rect 13820 12316 13872 12325
rect 16856 12316 16908 12368
rect 21824 12316 21876 12368
rect 12900 12248 12952 12300
rect 14832 12248 14884 12300
rect 15292 12291 15344 12300
rect 15292 12257 15336 12291
rect 15336 12257 15344 12291
rect 15292 12248 15344 12257
rect 16304 12248 16356 12300
rect 16948 12248 17000 12300
rect 18236 12248 18288 12300
rect 19340 12248 19392 12300
rect 20904 12248 20956 12300
rect 24952 12248 25004 12300
rect 1492 12180 1544 12232
rect 6644 12180 6696 12232
rect 10876 12180 10928 12232
rect 14372 12180 14424 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 22744 12180 22796 12232
rect 22836 12180 22888 12232
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 4528 12087 4580 12096
rect 4528 12053 4537 12087
rect 4537 12053 4571 12087
rect 4571 12053 4580 12087
rect 4528 12044 4580 12053
rect 4988 12044 5040 12096
rect 5540 12044 5592 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 9680 12044 9732 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 19800 12087 19852 12096
rect 19800 12053 19809 12087
rect 19809 12053 19843 12087
rect 19843 12053 19852 12087
rect 19800 12044 19852 12053
rect 20352 12044 20404 12096
rect 24860 12044 24912 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 7012 11840 7064 11892
rect 7748 11840 7800 11892
rect 8300 11840 8352 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 12900 11840 12952 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14372 11840 14424 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 16764 11883 16816 11892
rect 16764 11849 16773 11883
rect 16773 11849 16807 11883
rect 16807 11849 16816 11883
rect 16764 11840 16816 11849
rect 16948 11840 17000 11892
rect 19800 11840 19852 11892
rect 21824 11840 21876 11892
rect 22008 11840 22060 11892
rect 3424 11772 3476 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 3332 11636 3384 11688
rect 4252 11704 4304 11756
rect 4528 11704 4580 11756
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 4436 11679 4488 11688
rect 2136 11611 2188 11620
rect 2136 11577 2145 11611
rect 2145 11577 2179 11611
rect 2179 11577 2188 11611
rect 2136 11568 2188 11577
rect 3608 11568 3660 11620
rect 4436 11645 4445 11679
rect 4445 11645 4479 11679
rect 4479 11645 4488 11679
rect 4436 11636 4488 11645
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 8208 11636 8260 11688
rect 12348 11772 12400 11824
rect 13544 11704 13596 11756
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 15568 11636 15620 11688
rect 17408 11704 17460 11756
rect 15844 11636 15896 11688
rect 9128 11568 9180 11620
rect 9588 11611 9640 11620
rect 9588 11577 9597 11611
rect 9597 11577 9631 11611
rect 9631 11577 9640 11611
rect 9588 11568 9640 11577
rect 9680 11611 9732 11620
rect 9680 11577 9689 11611
rect 9689 11577 9723 11611
rect 9723 11577 9732 11611
rect 9680 11568 9732 11577
rect 1860 11500 1912 11552
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 9036 11500 9088 11552
rect 10140 11500 10192 11552
rect 11704 11500 11756 11552
rect 12440 11500 12492 11552
rect 13360 11568 13412 11620
rect 16212 11611 16264 11620
rect 16212 11577 16221 11611
rect 16221 11577 16255 11611
rect 16255 11577 16264 11611
rect 16212 11568 16264 11577
rect 18880 11772 18932 11824
rect 20904 11815 20956 11824
rect 20904 11781 20913 11815
rect 20913 11781 20947 11815
rect 20947 11781 20956 11815
rect 20904 11772 20956 11781
rect 20352 11704 20404 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22836 11704 22888 11756
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 24768 11840 24820 11892
rect 19156 11568 19208 11620
rect 19984 11611 20036 11620
rect 19984 11577 19993 11611
rect 19993 11577 20027 11611
rect 20027 11577 20036 11611
rect 19984 11568 20036 11577
rect 15844 11500 15896 11552
rect 18972 11543 19024 11552
rect 18972 11509 18981 11543
rect 18981 11509 19015 11543
rect 19015 11509 19024 11543
rect 18972 11500 19024 11509
rect 19524 11500 19576 11552
rect 22192 11611 22244 11620
rect 22192 11577 22201 11611
rect 22201 11577 22235 11611
rect 22235 11577 22244 11611
rect 22744 11611 22796 11620
rect 22192 11568 22244 11577
rect 22744 11577 22753 11611
rect 22753 11577 22787 11611
rect 22787 11577 22796 11611
rect 22744 11568 22796 11577
rect 22284 11500 22336 11552
rect 24952 11543 25004 11552
rect 24952 11509 24961 11543
rect 24961 11509 24995 11543
rect 24995 11509 25004 11543
rect 24952 11500 25004 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3240 11296 3292 11348
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 1952 11228 2004 11280
rect 4436 11296 4488 11348
rect 6276 11296 6328 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 5172 11228 5224 11280
rect 8668 11296 8720 11348
rect 2228 11160 2280 11212
rect 4160 11203 4212 11212
rect 4160 11169 4169 11203
rect 4169 11169 4203 11203
rect 4203 11169 4212 11203
rect 4528 11203 4580 11212
rect 4160 11160 4212 11169
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6736 11160 6788 11212
rect 6920 11228 6972 11280
rect 9772 11271 9824 11280
rect 9772 11237 9781 11271
rect 9781 11237 9815 11271
rect 9815 11237 9824 11271
rect 9772 11228 9824 11237
rect 11704 11296 11756 11348
rect 14740 11296 14792 11348
rect 15568 11339 15620 11348
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 12440 11271 12492 11280
rect 12440 11237 12449 11271
rect 12449 11237 12483 11271
rect 12483 11237 12492 11271
rect 12440 11228 12492 11237
rect 16856 11228 16908 11280
rect 18972 11228 19024 11280
rect 19156 11228 19208 11280
rect 20076 11228 20128 11280
rect 21088 11271 21140 11280
rect 21088 11237 21097 11271
rect 21097 11237 21131 11271
rect 21131 11237 21140 11271
rect 21088 11228 21140 11237
rect 22192 11228 22244 11280
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 11980 11160 12032 11212
rect 13820 11203 13872 11212
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 15752 11160 15804 11212
rect 21824 11160 21876 11212
rect 22560 11203 22612 11212
rect 22560 11169 22569 11203
rect 22569 11169 22603 11203
rect 22603 11169 22612 11203
rect 22560 11160 22612 11169
rect 24860 11160 24912 11212
rect 1308 11024 1360 11076
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 12532 11092 12584 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 19064 11092 19116 11144
rect 19340 11135 19392 11144
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 19340 11092 19392 11101
rect 20996 11135 21048 11144
rect 20996 11101 21005 11135
rect 21005 11101 21039 11135
rect 21039 11101 21048 11135
rect 20996 11092 21048 11101
rect 7564 11024 7616 11076
rect 2044 10956 2096 11008
rect 2228 10956 2280 11008
rect 7104 10956 7156 11008
rect 9036 11024 9088 11076
rect 13176 11024 13228 11076
rect 21548 11067 21600 11076
rect 21548 11033 21557 11067
rect 21557 11033 21591 11067
rect 21591 11033 21600 11067
rect 21548 11024 21600 11033
rect 24768 11067 24820 11076
rect 24768 11033 24777 11067
rect 24777 11033 24811 11067
rect 24811 11033 24820 11067
rect 24768 11024 24820 11033
rect 8116 10956 8168 11008
rect 8484 10956 8536 11008
rect 9588 10956 9640 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 12624 10956 12676 11008
rect 12808 10956 12860 11008
rect 14188 10956 14240 11008
rect 16488 10956 16540 11008
rect 17684 10999 17736 11008
rect 17684 10965 17693 10999
rect 17693 10965 17727 10999
rect 17727 10965 17736 10999
rect 17684 10956 17736 10965
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 19892 10999 19944 11008
rect 19892 10965 19901 10999
rect 19901 10965 19935 10999
rect 19935 10965 19944 10999
rect 19892 10956 19944 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 3424 10752 3476 10804
rect 4528 10752 4580 10804
rect 5448 10752 5500 10804
rect 7932 10752 7984 10804
rect 9772 10752 9824 10804
rect 17776 10752 17828 10804
rect 19892 10752 19944 10804
rect 20720 10752 20772 10804
rect 21088 10752 21140 10804
rect 22560 10795 22612 10804
rect 22560 10761 22569 10795
rect 22569 10761 22603 10795
rect 22603 10761 22612 10795
rect 22560 10752 22612 10761
rect 24860 10752 24912 10804
rect 2044 10684 2096 10736
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 2228 10480 2280 10532
rect 19524 10684 19576 10736
rect 20076 10727 20128 10736
rect 20076 10693 20085 10727
rect 20085 10693 20119 10727
rect 20119 10693 20128 10727
rect 20076 10684 20128 10693
rect 20996 10684 21048 10736
rect 22928 10684 22980 10736
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 4436 10591 4488 10600
rect 3240 10548 3292 10557
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 4804 10548 4856 10600
rect 5172 10616 5224 10668
rect 5080 10548 5132 10600
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 5356 10548 5408 10600
rect 6276 10548 6328 10600
rect 7380 10616 7432 10668
rect 7104 10591 7156 10600
rect 7104 10557 7113 10591
rect 7113 10557 7147 10591
rect 7147 10557 7156 10591
rect 7104 10548 7156 10557
rect 7564 10591 7616 10600
rect 7564 10557 7573 10591
rect 7573 10557 7607 10591
rect 7607 10557 7616 10591
rect 7564 10548 7616 10557
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 8944 10616 8996 10668
rect 12532 10659 12584 10668
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 16488 10659 16540 10668
rect 16488 10625 16497 10659
rect 16497 10625 16531 10659
rect 16531 10625 16540 10659
rect 16488 10616 16540 10625
rect 16764 10616 16816 10668
rect 19064 10616 19116 10668
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9496 10548 9548 10600
rect 14188 10548 14240 10600
rect 15568 10548 15620 10600
rect 21548 10548 21600 10600
rect 22744 10548 22796 10600
rect 1952 10412 2004 10464
rect 9036 10480 9088 10532
rect 10140 10480 10192 10532
rect 11060 10480 11112 10532
rect 12808 10480 12860 10532
rect 13176 10523 13228 10532
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 13912 10480 13964 10532
rect 14556 10480 14608 10532
rect 15752 10523 15804 10532
rect 15752 10489 15761 10523
rect 15761 10489 15795 10523
rect 15795 10489 15804 10523
rect 15752 10480 15804 10489
rect 17684 10480 17736 10532
rect 19064 10523 19116 10532
rect 19064 10489 19073 10523
rect 19073 10489 19107 10523
rect 19107 10489 19116 10523
rect 19064 10480 19116 10489
rect 19156 10523 19208 10532
rect 19156 10489 19165 10523
rect 19165 10489 19199 10523
rect 19199 10489 19208 10523
rect 20628 10523 20680 10532
rect 19156 10480 19208 10489
rect 20628 10489 20637 10523
rect 20637 10489 20671 10523
rect 20671 10489 20680 10523
rect 20628 10480 20680 10489
rect 20720 10523 20772 10532
rect 20720 10489 20729 10523
rect 20729 10489 20763 10523
rect 20763 10489 20772 10523
rect 20720 10480 20772 10489
rect 3424 10412 3476 10464
rect 5172 10412 5224 10464
rect 6736 10412 6788 10464
rect 8024 10412 8076 10464
rect 8668 10412 8720 10464
rect 9588 10412 9640 10464
rect 10968 10412 11020 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12348 10412 12400 10464
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 15660 10412 15712 10464
rect 16856 10412 16908 10464
rect 24584 10412 24636 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 7196 10208 7248 10260
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 10692 10208 10744 10260
rect 3056 10140 3108 10192
rect 4804 10140 4856 10192
rect 8668 10140 8720 10192
rect 11060 10140 11112 10192
rect 11612 10140 11664 10192
rect 12808 10183 12860 10192
rect 2228 10072 2280 10124
rect 3148 10072 3200 10124
rect 3700 10072 3752 10124
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 6828 10072 6880 10124
rect 6092 10004 6144 10056
rect 7012 10072 7064 10124
rect 8300 10072 8352 10124
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 9128 10072 9180 10124
rect 10140 10072 10192 10124
rect 12808 10149 12817 10183
rect 12817 10149 12851 10183
rect 12851 10149 12860 10183
rect 12808 10140 12860 10149
rect 13360 10183 13412 10192
rect 13360 10149 13369 10183
rect 13369 10149 13403 10183
rect 13403 10149 13412 10183
rect 13360 10140 13412 10149
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 14096 10208 14148 10260
rect 15384 10208 15436 10260
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 15476 10183 15528 10192
rect 15476 10149 15485 10183
rect 15485 10149 15519 10183
rect 15519 10149 15528 10183
rect 15476 10140 15528 10149
rect 15568 10140 15620 10192
rect 23664 10208 23716 10260
rect 16948 10140 17000 10192
rect 17684 10140 17736 10192
rect 19156 10140 19208 10192
rect 21088 10140 21140 10192
rect 13636 10072 13688 10124
rect 16212 10072 16264 10124
rect 17316 10072 17368 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 23572 10115 23624 10124
rect 23572 10081 23581 10115
rect 23581 10081 23615 10115
rect 23615 10081 23624 10115
rect 23572 10072 23624 10081
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 13728 10004 13780 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 18880 10047 18932 10056
rect 18880 10013 18889 10047
rect 18889 10013 18923 10047
rect 18923 10013 18932 10047
rect 18880 10004 18932 10013
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 5080 9936 5132 9988
rect 6736 9979 6788 9988
rect 6736 9945 6745 9979
rect 6745 9945 6779 9979
rect 6779 9945 6788 9979
rect 6736 9936 6788 9945
rect 7564 9936 7616 9988
rect 13544 9936 13596 9988
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 4068 9868 4120 9920
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 5264 9868 5316 9920
rect 9588 9868 9640 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 12900 9868 12952 9920
rect 13912 9868 13964 9920
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 19064 9868 19116 9920
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 20628 9911 20680 9920
rect 20628 9877 20637 9911
rect 20637 9877 20671 9911
rect 20671 9877 20680 9911
rect 20628 9868 20680 9877
rect 24768 9911 24820 9920
rect 24768 9877 24777 9911
rect 24777 9877 24811 9911
rect 24811 9877 24820 9911
rect 24768 9868 24820 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 20 9664 72 9716
rect 4344 9664 4396 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 6092 9664 6144 9716
rect 6828 9664 6880 9716
rect 8300 9664 8352 9716
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 4528 9596 4580 9648
rect 7840 9596 7892 9648
rect 3424 9528 3476 9580
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 6736 9528 6788 9580
rect 4252 9460 4304 9512
rect 5356 9460 5408 9512
rect 1676 9392 1728 9444
rect 2504 9392 2556 9444
rect 1400 9324 1452 9376
rect 3148 9324 3200 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 5080 9392 5132 9444
rect 7104 9460 7156 9512
rect 8392 9596 8444 9648
rect 14740 9664 14792 9716
rect 15476 9707 15528 9716
rect 15476 9673 15485 9707
rect 15485 9673 15519 9707
rect 15519 9673 15528 9707
rect 15476 9664 15528 9673
rect 15660 9664 15712 9716
rect 16856 9664 16908 9716
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 19892 9664 19944 9716
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 7564 9392 7616 9444
rect 8392 9460 8444 9512
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 7932 9392 7984 9444
rect 9128 9435 9180 9444
rect 9128 9401 9137 9435
rect 9137 9401 9171 9435
rect 9171 9401 9180 9435
rect 9128 9392 9180 9401
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 16028 9596 16080 9648
rect 23572 9596 23624 9648
rect 11612 9571 11664 9580
rect 11612 9537 11621 9571
rect 11621 9537 11655 9571
rect 11655 9537 11664 9571
rect 11612 9528 11664 9537
rect 13360 9528 13412 9580
rect 19340 9528 19392 9580
rect 19432 9528 19484 9580
rect 11060 9460 11112 9469
rect 12900 9460 12952 9512
rect 13268 9460 13320 9512
rect 14188 9503 14240 9512
rect 13544 9392 13596 9444
rect 14188 9469 14197 9503
rect 14197 9469 14231 9503
rect 14231 9469 14240 9503
rect 14188 9460 14240 9469
rect 19984 9460 20036 9512
rect 16028 9435 16080 9444
rect 16028 9401 16037 9435
rect 16037 9401 16071 9435
rect 16071 9401 16080 9435
rect 16028 9392 16080 9401
rect 18144 9435 18196 9444
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 15660 9324 15712 9376
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 20904 9435 20956 9444
rect 17776 9324 17828 9376
rect 20904 9401 20913 9435
rect 20913 9401 20947 9435
rect 20947 9401 20956 9435
rect 20904 9392 20956 9401
rect 19524 9324 19576 9376
rect 21640 9367 21692 9376
rect 21640 9333 21649 9367
rect 21649 9333 21683 9367
rect 21683 9333 21692 9367
rect 21640 9324 21692 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 3516 9120 3568 9172
rect 4160 9120 4212 9172
rect 6736 9120 6788 9172
rect 7564 9120 7616 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 9864 9163 9916 9172
rect 9864 9129 9873 9163
rect 9873 9129 9907 9163
rect 9907 9129 9916 9163
rect 9864 9120 9916 9129
rect 10876 9120 10928 9172
rect 12532 9120 12584 9172
rect 13176 9120 13228 9172
rect 16028 9120 16080 9172
rect 18144 9120 18196 9172
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 1952 9052 2004 9104
rect 2504 9052 2556 9104
rect 3240 9052 3292 9104
rect 5540 9052 5592 9104
rect 2412 8984 2464 9036
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 5080 8984 5132 9036
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 11612 9052 11664 9104
rect 12808 9052 12860 9104
rect 13452 9052 13504 9104
rect 13912 9052 13964 9104
rect 14648 9052 14700 9104
rect 15476 9095 15528 9104
rect 15476 9061 15485 9095
rect 15485 9061 15519 9095
rect 15519 9061 15528 9095
rect 15476 9052 15528 9061
rect 18052 9052 18104 9104
rect 18236 9052 18288 9104
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 9772 8984 9824 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 12348 8984 12400 9036
rect 13636 8984 13688 9036
rect 16120 8984 16172 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17408 8984 17460 9036
rect 18604 9027 18656 9036
rect 18604 8993 18613 9027
rect 18613 8993 18647 9027
rect 18647 8993 18656 9027
rect 18604 8984 18656 8993
rect 20168 8984 20220 9036
rect 20536 8984 20588 9036
rect 1584 8916 1636 8968
rect 1952 8848 2004 8900
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 11060 8916 11112 8968
rect 12624 8916 12676 8968
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13728 8916 13780 8968
rect 13912 8916 13964 8968
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 5448 8848 5500 8857
rect 8484 8848 8536 8900
rect 9864 8848 9916 8900
rect 16488 8916 16540 8968
rect 1860 8780 1912 8832
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 4068 8780 4120 8832
rect 4252 8780 4304 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 10140 8823 10192 8832
rect 10140 8789 10149 8823
rect 10149 8789 10183 8823
rect 10183 8789 10192 8823
rect 10140 8780 10192 8789
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 14188 8780 14240 8832
rect 19524 8848 19576 8900
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 19340 8780 19392 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2320 8576 2372 8628
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 4344 8619 4396 8628
rect 2780 8576 2832 8585
rect 2044 8551 2096 8560
rect 2044 8517 2053 8551
rect 2053 8517 2087 8551
rect 2087 8517 2096 8551
rect 2044 8508 2096 8517
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 4160 8508 4212 8560
rect 5356 8508 5408 8560
rect 7564 8576 7616 8628
rect 11612 8576 11664 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 15476 8576 15528 8628
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18236 8576 18288 8628
rect 18604 8576 18656 8628
rect 24768 8619 24820 8628
rect 24768 8585 24777 8619
rect 24777 8585 24811 8619
rect 24811 8585 24820 8619
rect 24768 8576 24820 8585
rect 6092 8508 6144 8560
rect 9496 8508 9548 8560
rect 13544 8508 13596 8560
rect 16948 8508 17000 8560
rect 17040 8508 17092 8560
rect 18696 8551 18748 8560
rect 18696 8517 18705 8551
rect 18705 8517 18739 8551
rect 18739 8517 18748 8551
rect 18696 8508 18748 8517
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 10140 8440 10192 8492
rect 10968 8440 11020 8492
rect 13268 8440 13320 8492
rect 13360 8440 13412 8492
rect 2412 8372 2464 8424
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1860 8304 1912 8356
rect 2872 8304 2924 8356
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4804 8415 4856 8424
rect 4620 8372 4672 8381
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 8392 8415 8444 8424
rect 2964 8236 3016 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 8668 8415 8720 8424
rect 7288 8279 7340 8288
rect 6552 8236 6604 8245
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 12348 8304 12400 8356
rect 13452 8372 13504 8424
rect 14188 8372 14240 8424
rect 13544 8304 13596 8356
rect 16764 8440 16816 8492
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 15844 8372 15896 8424
rect 17316 8372 17368 8424
rect 20076 8415 20128 8424
rect 9772 8279 9824 8288
rect 8208 8236 8260 8245
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 12532 8279 12584 8288
rect 12532 8245 12541 8279
rect 12541 8245 12575 8279
rect 12575 8245 12584 8279
rect 12532 8236 12584 8245
rect 14096 8236 14148 8288
rect 17408 8304 17460 8356
rect 18236 8347 18288 8356
rect 18236 8313 18245 8347
rect 18245 8313 18279 8347
rect 18279 8313 18288 8347
rect 18236 8304 18288 8313
rect 19432 8347 19484 8356
rect 19432 8313 19441 8347
rect 19441 8313 19475 8347
rect 19475 8313 19484 8347
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 20260 8372 20312 8424
rect 24216 8372 24268 8424
rect 19432 8304 19484 8313
rect 17224 8236 17276 8288
rect 18144 8236 18196 8288
rect 19340 8236 19392 8288
rect 19524 8236 19576 8288
rect 20536 8236 20588 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 4620 8032 4672 8084
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 8576 8032 8628 8084
rect 9036 8032 9088 8084
rect 6552 7964 6604 8016
rect 9772 8032 9824 8084
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3332 7896 3384 7948
rect 4160 7939 4212 7948
rect 4160 7905 4169 7939
rect 4169 7905 4203 7939
rect 4203 7905 4212 7939
rect 4160 7896 4212 7905
rect 4344 7896 4396 7948
rect 5540 7896 5592 7948
rect 7196 7896 7248 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 8392 7896 8444 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 12532 8032 12584 8084
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 14188 8032 14240 8084
rect 4620 7828 4672 7880
rect 6828 7828 6880 7880
rect 6000 7760 6052 7812
rect 11612 7828 11664 7880
rect 12624 7896 12676 7948
rect 14096 7964 14148 8016
rect 15844 8007 15896 8016
rect 15844 7973 15853 8007
rect 15853 7973 15887 8007
rect 15887 7973 15896 8007
rect 15844 7964 15896 7973
rect 16304 7964 16356 8016
rect 18328 7964 18380 8016
rect 18880 8032 18932 8084
rect 20168 8032 20220 8084
rect 19524 7964 19576 8016
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 20168 7896 20220 7948
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 2044 7692 2096 7744
rect 2504 7692 2556 7744
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 8208 7760 8260 7812
rect 13268 7760 13320 7812
rect 6920 7692 6972 7701
rect 8668 7692 8720 7744
rect 11336 7692 11388 7744
rect 13452 7692 13504 7744
rect 15936 7760 15988 7812
rect 18144 7828 18196 7880
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 19524 7828 19576 7880
rect 16948 7760 17000 7812
rect 20076 7760 20128 7812
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 18236 7692 18288 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 5448 7488 5500 7540
rect 5540 7488 5592 7540
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 7564 7488 7616 7540
rect 3424 7420 3476 7472
rect 1860 7352 1912 7404
rect 2320 7352 2372 7404
rect 3332 7352 3384 7404
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 9680 7488 9732 7540
rect 11612 7488 11664 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 20904 7488 20956 7540
rect 9036 7463 9088 7472
rect 9036 7429 9045 7463
rect 9045 7429 9079 7463
rect 9079 7429 9088 7463
rect 9036 7420 9088 7429
rect 14648 7463 14700 7472
rect 14648 7429 14657 7463
rect 14657 7429 14691 7463
rect 14691 7429 14700 7463
rect 14648 7420 14700 7429
rect 17040 7463 17092 7472
rect 17040 7429 17049 7463
rect 17049 7429 17083 7463
rect 17083 7429 17092 7463
rect 17040 7420 17092 7429
rect 18236 7420 18288 7472
rect 2504 7284 2556 7336
rect 2964 7148 3016 7200
rect 3424 7148 3476 7200
rect 7840 7327 7892 7336
rect 7380 7216 7432 7268
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 8944 7327 8996 7336
rect 8944 7293 8953 7327
rect 8953 7293 8987 7327
rect 8987 7293 8996 7327
rect 8944 7284 8996 7293
rect 11612 7352 11664 7404
rect 12992 7352 13044 7404
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 14924 7352 14976 7404
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 17592 7284 17644 7336
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 12624 7259 12676 7268
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 14188 7259 14240 7268
rect 14188 7225 14197 7259
rect 14197 7225 14231 7259
rect 14231 7225 14240 7259
rect 14188 7216 14240 7225
rect 15568 7216 15620 7268
rect 16304 7216 16356 7268
rect 18420 7352 18472 7404
rect 18604 7352 18656 7404
rect 20536 7284 20588 7336
rect 18144 7259 18196 7268
rect 6184 7148 6236 7200
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 6552 7148 6604 7157
rect 7656 7191 7708 7200
rect 7656 7157 7665 7191
rect 7665 7157 7699 7191
rect 7699 7157 7708 7191
rect 7656 7148 7708 7157
rect 8208 7148 8260 7200
rect 15752 7148 15804 7200
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 18328 7216 18380 7268
rect 18788 7259 18840 7268
rect 18420 7148 18472 7200
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2228 6944 2280 6996
rect 5264 6987 5316 6996
rect 5264 6953 5273 6987
rect 5273 6953 5307 6987
rect 5307 6953 5316 6987
rect 5264 6944 5316 6953
rect 5356 6944 5408 6996
rect 7380 6944 7432 6996
rect 9036 6944 9088 6996
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 11060 6944 11112 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 16488 6944 16540 6996
rect 18512 6944 18564 6996
rect 2504 6876 2556 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 2688 6808 2740 6860
rect 3700 6808 3752 6860
rect 6000 6876 6052 6928
rect 8300 6876 8352 6928
rect 8668 6876 8720 6928
rect 11704 6876 11756 6928
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 7380 6851 7432 6860
rect 1492 6740 1544 6792
rect 5080 6740 5132 6792
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 9496 6808 9548 6860
rect 10140 6851 10192 6860
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 11796 6851 11848 6860
rect 11796 6817 11805 6851
rect 11805 6817 11839 6851
rect 11839 6817 11848 6851
rect 11796 6808 11848 6817
rect 12900 6808 12952 6860
rect 13452 6808 13504 6860
rect 15568 6876 15620 6928
rect 18236 6876 18288 6928
rect 14832 6808 14884 6860
rect 17868 6808 17920 6860
rect 19616 6808 19668 6860
rect 24676 6808 24728 6860
rect 10692 6740 10744 6792
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 15476 6783 15528 6792
rect 9036 6672 9088 6724
rect 11520 6672 11572 6724
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 19248 6740 19300 6792
rect 14924 6715 14976 6724
rect 14924 6681 14933 6715
rect 14933 6681 14967 6715
rect 14967 6681 14976 6715
rect 14924 6672 14976 6681
rect 2596 6604 2648 6656
rect 5356 6604 5408 6656
rect 6552 6604 6604 6656
rect 7932 6604 7984 6656
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 15752 6604 15804 6656
rect 18144 6672 18196 6724
rect 18604 6672 18656 6724
rect 18788 6715 18840 6724
rect 18788 6681 18797 6715
rect 18797 6681 18831 6715
rect 18831 6681 18840 6715
rect 18788 6672 18840 6681
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1400 6400 1452 6452
rect 5080 6400 5132 6452
rect 6000 6400 6052 6452
rect 6552 6332 6604 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 6092 6264 6144 6316
rect 1952 6196 2004 6248
rect 2504 6196 2556 6248
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2964 6239 3016 6248
rect 2780 6196 2832 6205
rect 2964 6205 2973 6239
rect 2973 6205 3007 6239
rect 3007 6205 3016 6239
rect 2964 6196 3016 6205
rect 7288 6400 7340 6452
rect 7840 6400 7892 6452
rect 10140 6400 10192 6452
rect 15476 6400 15528 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 20168 6400 20220 6452
rect 27620 6400 27672 6452
rect 7932 6332 7984 6384
rect 9496 6375 9548 6384
rect 9496 6341 9505 6375
rect 9505 6341 9539 6375
rect 9539 6341 9548 6375
rect 9496 6332 9548 6341
rect 13452 6332 13504 6384
rect 8116 6264 8168 6316
rect 9036 6264 9088 6316
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 11796 6264 11848 6316
rect 6828 6239 6880 6248
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 5448 6128 5500 6180
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 6184 6128 6236 6137
rect 1032 6060 1084 6112
rect 1584 6060 1636 6112
rect 5080 6060 5132 6112
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 8944 6060 8996 6112
rect 10048 6128 10100 6180
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 15384 6264 15436 6316
rect 18144 6264 18196 6316
rect 18788 6264 18840 6316
rect 19616 6307 19668 6316
rect 19616 6273 19625 6307
rect 19625 6273 19659 6307
rect 19659 6273 19668 6307
rect 19616 6264 19668 6273
rect 12900 6196 12952 6205
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 15936 6239 15988 6248
rect 15936 6205 15945 6239
rect 15945 6205 15979 6239
rect 15979 6205 15988 6239
rect 15936 6196 15988 6205
rect 20168 6196 20220 6248
rect 13084 6128 13136 6180
rect 15660 6128 15712 6180
rect 18328 6171 18380 6180
rect 12256 6060 12308 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 18328 6137 18337 6171
rect 18337 6137 18371 6171
rect 18371 6137 18380 6171
rect 18328 6128 18380 6137
rect 18604 6128 18656 6180
rect 17776 6060 17828 6112
rect 24676 6103 24728 6112
rect 24676 6069 24685 6103
rect 24685 6069 24719 6103
rect 24719 6069 24728 6103
rect 24676 6060 24728 6069
rect 26884 6060 26936 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1492 5856 1544 5908
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2780 5899 2832 5908
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 3056 5856 3108 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4896 5856 4948 5908
rect 6460 5856 6512 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 11704 5856 11756 5908
rect 12992 5856 13044 5908
rect 5264 5788 5316 5840
rect 7748 5788 7800 5840
rect 8944 5788 8996 5840
rect 9220 5788 9272 5840
rect 9864 5831 9916 5840
rect 9864 5797 9873 5831
rect 9873 5797 9907 5831
rect 9907 5797 9916 5831
rect 9864 5788 9916 5797
rect 11888 5788 11940 5840
rect 1768 5720 1820 5772
rect 3424 5720 3476 5772
rect 4344 5720 4396 5772
rect 4988 5720 5040 5772
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 7656 5720 7708 5772
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 13820 5763 13872 5772
rect 13820 5729 13829 5763
rect 13829 5729 13863 5763
rect 13863 5729 13872 5763
rect 13820 5720 13872 5729
rect 5080 5652 5132 5704
rect 9956 5652 10008 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11336 5652 11388 5704
rect 14832 5856 14884 5908
rect 15936 5856 15988 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 15384 5788 15436 5840
rect 15752 5788 15804 5840
rect 17132 5788 17184 5840
rect 16488 5720 16540 5772
rect 18604 5788 18656 5840
rect 19524 5831 19576 5840
rect 19524 5797 19533 5831
rect 19533 5797 19567 5831
rect 19567 5797 19576 5831
rect 19524 5788 19576 5797
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 17592 5652 17644 5704
rect 19800 5652 19852 5704
rect 14188 5584 14240 5636
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 18604 5559 18656 5568
rect 18604 5525 18613 5559
rect 18613 5525 18647 5559
rect 18647 5525 18656 5559
rect 18604 5516 18656 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1400 5312 1452 5364
rect 1768 5312 1820 5364
rect 3608 5312 3660 5364
rect 7656 5312 7708 5364
rect 9956 5312 10008 5364
rect 12072 5312 12124 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 15384 5355 15436 5364
rect 13820 5312 13872 5321
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 19800 5355 19852 5364
rect 19800 5321 19809 5355
rect 19809 5321 19843 5355
rect 19843 5321 19852 5355
rect 19800 5312 19852 5321
rect 3884 5244 3936 5296
rect 1124 5108 1176 5160
rect 1952 5108 2004 5160
rect 3608 5108 3660 5160
rect 5264 5244 5316 5296
rect 5540 5176 5592 5228
rect 4896 5108 4948 5160
rect 2044 5040 2096 5092
rect 7748 5244 7800 5296
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 4528 4972 4580 5024
rect 4896 4972 4948 5024
rect 6092 5040 6144 5092
rect 7564 5083 7616 5092
rect 6000 4972 6052 5024
rect 7564 5049 7573 5083
rect 7573 5049 7607 5083
rect 7607 5049 7616 5083
rect 7564 5040 7616 5049
rect 11888 5244 11940 5296
rect 12624 5244 12676 5296
rect 9772 5176 9824 5228
rect 10140 5176 10192 5228
rect 14740 5176 14792 5228
rect 18696 5176 18748 5228
rect 10692 5108 10744 5160
rect 15292 5108 15344 5160
rect 21640 5244 21692 5296
rect 27620 5244 27672 5296
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 11520 4972 11572 5024
rect 14188 5083 14240 5092
rect 14188 5049 14197 5083
rect 14197 5049 14231 5083
rect 14231 5049 14240 5083
rect 14188 5040 14240 5049
rect 14740 5083 14792 5092
rect 14740 5049 14749 5083
rect 14749 5049 14783 5083
rect 14783 5049 14792 5083
rect 14740 5040 14792 5049
rect 15476 4972 15528 5024
rect 17132 5083 17184 5092
rect 17132 5049 17141 5083
rect 17141 5049 17175 5083
rect 17175 5049 17184 5083
rect 17132 5040 17184 5049
rect 18512 5083 18564 5092
rect 18512 5049 18521 5083
rect 18521 5049 18555 5083
rect 18555 5049 18564 5083
rect 18512 5040 18564 5049
rect 18604 5083 18656 5092
rect 18604 5049 18613 5083
rect 18613 5049 18647 5083
rect 18647 5049 18656 5083
rect 18604 5040 18656 5049
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1308 4768 1360 4820
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5172 4768 5224 4820
rect 6460 4700 6512 4752
rect 6920 4700 6972 4752
rect 7564 4768 7616 4820
rect 9772 4768 9824 4820
rect 12256 4768 12308 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 14188 4768 14240 4820
rect 15568 4768 15620 4820
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 9864 4743 9916 4752
rect 9864 4709 9873 4743
rect 9873 4709 9907 4743
rect 9907 4709 9916 4743
rect 9864 4700 9916 4709
rect 10692 4700 10744 4752
rect 1676 4632 1728 4684
rect 2136 4632 2188 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 7932 4632 7984 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8576 4632 8628 4684
rect 10048 4632 10100 4684
rect 15476 4700 15528 4752
rect 16856 4700 16908 4752
rect 17408 4700 17460 4752
rect 18328 4700 18380 4752
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 6276 4564 6328 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 17684 4607 17736 4616
rect 8116 4539 8168 4548
rect 8116 4505 8125 4539
rect 8125 4505 8159 4539
rect 8159 4505 8168 4539
rect 8116 4496 8168 4505
rect 14372 4496 14424 4548
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 17960 4496 18012 4548
rect 18696 4496 18748 4548
rect 11888 4428 11940 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 9220 4267 9272 4276
rect 5632 4156 5684 4208
rect 8576 4156 8628 4208
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 10508 4224 10560 4276
rect 12624 4224 12676 4276
rect 13636 4267 13688 4276
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 16304 4267 16356 4276
rect 16304 4233 16313 4267
rect 16313 4233 16347 4267
rect 16347 4233 16356 4267
rect 16304 4224 16356 4233
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18236 4224 18288 4276
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7932 4088 7984 4140
rect 9588 4088 9640 4140
rect 11888 4088 11940 4140
rect 15384 4156 15436 4208
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 17684 4088 17736 4140
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 24032 4088 24084 4140
rect 5264 4020 5316 4072
rect 13636 4020 13688 4072
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 6000 3952 6052 4004
rect 7380 3952 7432 4004
rect 10048 3995 10100 4004
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 9220 3884 9272 3936
rect 10048 3961 10057 3995
rect 10057 3961 10091 3995
rect 10091 3961 10100 3995
rect 10048 3952 10100 3961
rect 10140 3952 10192 4004
rect 12624 3952 12676 4004
rect 12900 3952 12952 4004
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 14372 3995 14424 4004
rect 14372 3961 14381 3995
rect 14381 3961 14415 3995
rect 14415 3961 14424 3995
rect 14372 3952 14424 3961
rect 14740 3952 14792 4004
rect 16212 3952 16264 4004
rect 16304 3952 16356 4004
rect 18144 3995 18196 4004
rect 18144 3961 18153 3995
rect 18153 3961 18187 3995
rect 18187 3961 18196 3995
rect 18144 3952 18196 3961
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 10692 3884 10744 3936
rect 11336 3884 11388 3936
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 14188 3884 14240 3936
rect 15476 3884 15528 3936
rect 27620 3884 27672 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5632 3680 5684 3732
rect 6000 3680 6052 3732
rect 7380 3723 7432 3732
rect 5908 3612 5960 3664
rect 6460 3612 6512 3664
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 9588 3680 9640 3732
rect 7196 3612 7248 3664
rect 9220 3612 9272 3664
rect 1768 3544 1820 3596
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 6920 3476 6972 3528
rect 7196 3476 7248 3528
rect 8300 3476 8352 3528
rect 9772 3612 9824 3664
rect 10048 3612 10100 3664
rect 11428 3655 11480 3664
rect 11428 3621 11437 3655
rect 11437 3621 11471 3655
rect 11471 3621 11480 3655
rect 11428 3612 11480 3621
rect 12624 3680 12676 3732
rect 14188 3680 14240 3732
rect 14372 3680 14424 3732
rect 14832 3680 14884 3732
rect 15384 3723 15436 3732
rect 12900 3655 12952 3664
rect 12900 3621 12909 3655
rect 12909 3621 12943 3655
rect 12943 3621 12952 3655
rect 12900 3612 12952 3621
rect 13360 3612 13412 3664
rect 14740 3612 14792 3664
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 18144 3680 18196 3732
rect 15476 3612 15528 3664
rect 17592 3655 17644 3664
rect 14280 3544 14332 3596
rect 15568 3587 15620 3596
rect 15568 3553 15577 3587
rect 15577 3553 15611 3587
rect 15611 3553 15620 3587
rect 15568 3544 15620 3553
rect 17132 3587 17184 3596
rect 17132 3553 17141 3587
rect 17141 3553 17175 3587
rect 17175 3553 17184 3587
rect 17132 3544 17184 3553
rect 17592 3621 17601 3655
rect 17601 3621 17635 3655
rect 17635 3621 17644 3655
rect 17592 3612 17644 3621
rect 17408 3544 17460 3596
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 10692 3476 10744 3528
rect 11704 3476 11756 3528
rect 7840 3408 7892 3460
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 10140 3408 10192 3460
rect 12716 3408 12768 3460
rect 18144 3408 18196 3460
rect 6276 3340 6328 3349
rect 9864 3340 9916 3392
rect 17500 3340 17552 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1768 3136 1820 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 6460 3179 6512 3188
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 6920 3136 6972 3188
rect 9220 3136 9272 3188
rect 9772 3136 9824 3188
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 11612 3136 11664 3188
rect 7564 3000 7616 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8760 3000 8812 3052
rect 9864 3068 9916 3120
rect 10140 3068 10192 3120
rect 10968 3068 11020 3120
rect 11520 3000 11572 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 112 2932 164 2984
rect 5632 2932 5684 2984
rect 6000 2932 6052 2984
rect 13360 3136 13412 3188
rect 13452 3136 13504 3188
rect 13728 3068 13780 3120
rect 12900 3000 12952 3052
rect 14556 2932 14608 2984
rect 15568 3136 15620 3188
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 17408 3136 17460 3188
rect 18420 3179 18472 3188
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 17500 2932 17552 2984
rect 4436 2796 4488 2848
rect 5724 2796 5776 2848
rect 8300 2864 8352 2916
rect 8576 2796 8628 2848
rect 8760 2796 8812 2848
rect 11520 2864 11572 2916
rect 15384 2864 15436 2916
rect 14556 2839 14608 2848
rect 14556 2805 14565 2839
rect 14565 2805 14599 2839
rect 14599 2805 14608 2839
rect 14556 2796 14608 2805
rect 15292 2839 15344 2848
rect 15292 2805 15301 2839
rect 15301 2805 15335 2839
rect 15335 2805 15344 2839
rect 15292 2796 15344 2805
rect 16764 2839 16816 2848
rect 16764 2805 16773 2839
rect 16773 2805 16807 2839
rect 16807 2805 16816 2839
rect 16764 2796 16816 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7104 2592 7156 2644
rect 7748 2635 7800 2644
rect 7196 2524 7248 2576
rect 3516 2456 3568 2508
rect 4896 2456 4948 2508
rect 5724 2499 5776 2508
rect 5724 2465 5733 2499
rect 5733 2465 5767 2499
rect 5767 2465 5776 2499
rect 5724 2456 5776 2465
rect 7748 2601 7757 2635
rect 7757 2601 7791 2635
rect 7791 2601 7800 2635
rect 7748 2592 7800 2601
rect 8760 2635 8812 2644
rect 8760 2601 8769 2635
rect 8769 2601 8803 2635
rect 8803 2601 8812 2635
rect 8760 2592 8812 2601
rect 10692 2592 10744 2644
rect 17684 2592 17736 2644
rect 18144 2592 18196 2644
rect 20628 2592 20680 2644
rect 17500 2567 17552 2576
rect 17500 2533 17509 2567
rect 17509 2533 17543 2567
rect 17543 2533 17552 2567
rect 17500 2524 17552 2533
rect 19064 2524 19116 2576
rect 8576 2456 8628 2508
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 11520 2456 11572 2508
rect 13636 2456 13688 2508
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 14556 2388 14608 2440
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 4896 2295 4948 2304
rect 4896 2261 4905 2295
rect 4905 2261 4939 2295
rect 4939 2261 4948 2295
rect 4896 2252 4948 2261
rect 10048 2320 10100 2372
rect 16212 2456 16264 2508
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 23204 2388 23256 2440
rect 24676 2320 24728 2372
rect 9312 2252 9364 2304
rect 9864 2252 9916 2304
rect 14372 2295 14424 2304
rect 14372 2261 14381 2295
rect 14381 2261 14415 2295
rect 14415 2261 14424 2295
rect 14372 2252 14424 2261
rect 23204 2252 23256 2304
rect 26056 2252 26108 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 14556 2048 14608 2100
rect 20260 2048 20312 2100
rect 14372 76 14424 128
rect 23296 76 23348 128
<< metal2 >>
rect 124 27526 520 27554
rect 124 23474 152 27526
rect 492 27520 520 27526
rect 570 27520 626 28000
rect 1766 27520 1822 28000
rect 1872 27526 2176 27554
rect 1872 27520 1900 27526
rect 492 27492 612 27520
rect 1780 27492 1900 27520
rect 1858 26752 1914 26761
rect 1858 26687 1914 26696
rect 1306 25528 1362 25537
rect 1306 25463 1362 25472
rect 1320 23662 1348 25463
rect 1872 24274 1900 26687
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1582 24168 1638 24177
rect 1582 24103 1638 24112
rect 1308 23656 1360 23662
rect 1308 23598 1360 23604
rect 1398 23624 1454 23633
rect 1398 23559 1454 23568
rect 1412 23526 1440 23559
rect 32 23446 152 23474
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 32 9722 60 23446
rect 1596 23186 1624 24103
rect 1872 23866 1900 24210
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1398 22944 1454 22953
rect 1398 22879 1454 22888
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 112 18080 164 18086
rect 112 18022 164 18028
rect 124 17105 152 18022
rect 110 17096 166 17105
rect 110 17031 166 17040
rect 112 16992 164 16998
rect 112 16934 164 16940
rect 124 10713 152 16934
rect 110 10704 166 10713
rect 110 10639 166 10648
rect 20 9716 72 9722
rect 20 9658 72 9664
rect 1032 6112 1084 6118
rect 1032 6054 1084 6060
rect 110 3088 166 3097
rect 110 3023 166 3032
rect 124 2990 152 3023
rect 112 2984 164 2990
rect 112 2926 164 2932
rect 662 82 718 480
rect 1044 82 1072 6054
rect 1136 5166 1164 19246
rect 1412 18834 1440 22879
rect 1596 22778 1624 23122
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1582 21720 1638 21729
rect 1582 21655 1638 21664
rect 1596 21146 1624 21655
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1952 21004 2004 21010
rect 1952 20946 2004 20952
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1596 19514 1624 20295
rect 1964 20262 1992 20946
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1490 19136 1546 19145
rect 1490 19071 1546 19080
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18426 1440 18770
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 1504 15162 1532 19071
rect 1582 18048 1638 18057
rect 1582 17983 1638 17992
rect 1596 17882 1624 17983
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 17105 1624 17682
rect 1964 17241 1992 20198
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 17882 2084 19110
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 1950 17232 2006 17241
rect 1950 17167 2006 17176
rect 1582 17096 1638 17105
rect 1582 17031 1638 17040
rect 1596 16980 1624 17031
rect 1676 16992 1728 16998
rect 1596 16952 1676 16980
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1412 14521 1440 14894
rect 1398 14512 1454 14521
rect 1398 14447 1454 14456
rect 1596 13814 1624 16952
rect 1676 16934 1728 16940
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15638 1716 15846
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1688 15162 1716 15574
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1596 13786 1716 13814
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1596 12345 1624 12378
rect 1582 12336 1638 12345
rect 1308 12300 1360 12306
rect 1582 12271 1638 12280
rect 1308 12242 1360 12248
rect 1320 11082 1348 12242
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 11762 1532 12174
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1308 11076 1360 11082
rect 1308 11018 1360 11024
rect 1124 5160 1176 5166
rect 1124 5102 1176 5108
rect 1320 4826 1348 11018
rect 1688 9568 1716 13786
rect 1780 12850 1808 16730
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16454 1900 16594
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1872 13569 1900 16390
rect 1964 15201 1992 17167
rect 2056 17134 2084 17818
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16425 2084 16934
rect 2042 16416 2098 16425
rect 2042 16351 2098 16360
rect 1950 15192 2006 15201
rect 1950 15127 2006 15136
rect 2148 13814 2176 27526
rect 3054 27532 3110 28000
rect 3054 27520 3056 27532
rect 3108 27520 3110 27532
rect 3884 27532 3936 27538
rect 3056 27474 3108 27480
rect 4342 27520 4398 28000
rect 5630 27554 5686 28000
rect 6918 27554 6974 28000
rect 5630 27526 6040 27554
rect 5630 27520 5686 27526
rect 3884 27474 3936 27480
rect 3068 27443 3096 27474
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 18737 2728 24006
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 2964 18760 3016 18766
rect 2686 18728 2742 18737
rect 2964 18702 3016 18708
rect 2686 18663 2742 18672
rect 2976 18290 3004 18702
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2332 16794 2360 17478
rect 2516 16998 2544 17682
rect 3068 17610 3096 19110
rect 3436 18970 3464 19110
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3528 17882 3556 18226
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16046 2360 16390
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 14822 2360 15982
rect 2516 15910 2544 16594
rect 2884 16250 2912 16594
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2424 15026 2452 15574
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 2056 13786 2176 13814
rect 1858 13560 1914 13569
rect 1858 13495 1914 13504
rect 1964 13462 1992 13738
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 1964 13258 1992 13398
rect 2056 13394 2084 13786
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1964 12646 1992 13194
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 10266 1900 11494
rect 1964 11286 1992 12582
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1964 10470 1992 11222
rect 2056 11014 2084 13126
rect 2148 12714 2176 13670
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1688 9540 1808 9568
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1412 6458 1440 9318
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 6798 1532 8298
rect 1596 8090 1624 8910
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1688 7546 1716 9386
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1412 5370 1440 6394
rect 1504 5914 1532 6734
rect 1596 6118 1624 6802
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1780 5778 1808 9540
rect 1964 9110 1992 10406
rect 2056 9654 2084 10678
rect 2148 10674 2176 11562
rect 2240 11218 2268 14214
rect 2332 13734 2360 14758
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8362 1900 8774
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1872 7410 1900 8298
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1964 6254 1992 8842
rect 2056 8566 2084 9590
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1964 5914 1992 6190
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1780 5370 1808 5714
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4282 1716 4626
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1964 4049 1992 5102
rect 2056 5098 2084 7686
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1766 4040 1822 4049
rect 1766 3975 1822 3984
rect 1950 4040 2006 4049
rect 1950 3975 2006 3984
rect 1780 3602 1808 3975
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3194 1808 3538
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 662 54 1072 82
rect 1950 82 2006 480
rect 2056 82 2084 5034
rect 2148 4690 2176 10610
rect 2240 10538 2268 10950
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2240 10130 2268 10474
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2240 7002 2268 10066
rect 2332 8634 2360 13330
rect 2424 12850 2452 14962
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2516 10248 2544 15846
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2608 13938 2636 15302
rect 2700 14890 2728 15302
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2700 13530 2728 14826
rect 2780 14544 2832 14550
rect 2976 14521 3004 17478
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3160 16114 3188 16526
rect 3436 16454 3464 17614
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3160 14550 3188 15030
rect 3148 14544 3200 14550
rect 2780 14486 2832 14492
rect 2962 14512 3018 14521
rect 2792 13734 2820 14486
rect 3148 14486 3200 14492
rect 2962 14447 3018 14456
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2792 13462 2820 13670
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 3160 12986 3188 13942
rect 3252 13326 3280 15846
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3160 12782 3188 12922
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 10266 3188 12582
rect 3344 11778 3372 15982
rect 3436 15502 3464 16390
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14346 3648 14758
rect 3712 14362 3740 20198
rect 3804 18873 3832 22918
rect 3790 18864 3846 18873
rect 3790 18799 3846 18808
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 15638 3832 16390
rect 3896 16250 3924 27474
rect 4356 23730 4384 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24274 6040 27526
rect 6918 27526 7236 27554
rect 6918 27520 6974 27526
rect 6920 26648 6972 26654
rect 6920 26590 6972 26596
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6656 20262 6684 20946
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3988 18154 4016 19790
rect 5000 19514 5028 19858
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4988 19508 5040 19514
rect 4988 19450 5040 19456
rect 4080 19258 4108 19450
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4080 19242 4200 19258
rect 4080 19236 4212 19242
rect 4080 19230 4160 19236
rect 4160 19178 4212 19184
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 4172 18086 4200 19178
rect 4356 18290 4384 19314
rect 5276 19310 5304 20198
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5092 18426 5120 18838
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4816 18329 4844 18362
rect 4802 18320 4858 18329
rect 4344 18284 4396 18290
rect 4802 18255 4858 18264
rect 4344 18226 4396 18232
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4356 17882 4384 18226
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 4724 17338 4752 17750
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 5184 17202 5212 17546
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5276 16794 5304 18090
rect 5368 17746 5396 18702
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5552 18290 5580 18634
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 20198
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5722 18320 5778 18329
rect 5540 18284 5592 18290
rect 6288 18290 6316 20198
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6564 19514 6592 19858
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 5722 18255 5778 18264
rect 6276 18284 6328 18290
rect 5540 18226 5592 18232
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5552 17270 5580 18226
rect 5736 18222 5764 18255
rect 6276 18226 6328 18232
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5644 17649 5672 17682
rect 6184 17672 6236 17678
rect 5630 17640 5686 17649
rect 6184 17614 6236 17620
rect 5630 17575 5686 17584
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3896 16046 3924 16186
rect 4448 16046 4476 16390
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4448 15706 4476 15982
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 4632 15570 4660 16118
rect 4816 15910 4844 16662
rect 5368 16250 5396 17002
rect 5552 16794 5580 17206
rect 6196 16998 6224 17614
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15638 4844 15846
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4632 15162 4660 15506
rect 4988 15428 5040 15434
rect 4988 15370 5040 15376
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4632 14958 4660 15098
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4356 14618 4384 14826
rect 4632 14618 4660 14894
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4632 14482 4660 14554
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 3608 14340 3660 14346
rect 3712 14334 3924 14362
rect 3608 14282 3660 14288
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3528 13734 3556 13874
rect 3712 13814 3740 14214
rect 3896 14006 3924 14334
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14006 4200 14214
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3896 13870 3924 13942
rect 3884 13864 3936 13870
rect 3712 13786 3832 13814
rect 3884 13806 3936 13812
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3528 12850 3556 13670
rect 3804 13530 3832 13786
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3606 12744 3662 12753
rect 3436 11830 3464 12718
rect 3606 12679 3662 12688
rect 3252 11750 3372 11778
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3252 11354 3280 11750
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3252 10606 3280 11290
rect 3344 10810 3372 11630
rect 3436 11354 3464 11766
rect 3620 11762 3648 12679
rect 3712 12646 3740 13262
rect 4264 12782 4292 13806
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4448 12782 4476 12854
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 4264 12442 4292 12718
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3424 11348 3476 11354
rect 3476 11308 3556 11336
rect 3424 11290 3476 11296
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3148 10260 3200 10266
rect 2516 10220 2636 10248
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9432 2452 9862
rect 2504 9444 2556 9450
rect 2424 9404 2504 9432
rect 2424 9042 2452 9404
rect 2504 9386 2556 9392
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2332 5914 2360 7346
rect 2424 7324 2452 8366
rect 2516 7750 2544 9046
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2504 7336 2556 7342
rect 2424 7296 2504 7324
rect 2504 7278 2556 7284
rect 2516 6934 2544 7278
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2516 6254 2544 6870
rect 2608 6662 2636 10220
rect 3148 10202 3200 10208
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2700 6866 2728 9551
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2792 6254 2820 8570
rect 2976 8430 3004 8774
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 8090 2912 8298
rect 2976 8294 3004 8366
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7206 3004 7890
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6254 3004 7142
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2792 5914 2820 6190
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 1950 54 2084 82
rect 2976 82 3004 6190
rect 3068 5914 3096 10134
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3160 9382 3188 10066
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 6322 3188 9318
rect 3252 9110 3280 10542
rect 3436 10470 3464 10746
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3436 9586 3464 10406
rect 3528 10266 3556 11308
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9382 3464 9522
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3436 8072 3464 9318
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3436 8044 3556 8072
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7410 3372 7890
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7478 3464 7686
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3424 7200 3476 7206
rect 3528 7188 3556 8044
rect 3620 7410 3648 11562
rect 3896 11354 3924 12310
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 8498 3740 10066
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3476 7160 3556 7188
rect 3424 7142 3476 7148
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3436 5778 3464 7142
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3436 5030 3464 5714
rect 3620 5370 3648 7346
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3712 6322 3740 6802
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3620 5166 3648 5306
rect 3896 5302 3924 9862
rect 4080 8838 4108 9862
rect 4172 9178 4200 11154
rect 4264 10266 4292 11698
rect 4448 11694 4476 12242
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11762 4568 12038
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4448 11354 4476 11630
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4448 10606 4476 11290
rect 4528 11212 4580 11218
rect 4816 11200 4844 14758
rect 5000 12782 5028 15370
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 12368 4948 12374
rect 5000 12356 5028 12718
rect 4948 12328 5028 12356
rect 4896 12310 4948 12316
rect 5000 12102 5028 12328
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5092 11336 5120 15914
rect 5552 15910 5580 16526
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6104 16250 6132 16594
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5172 15564 5224 15570
rect 5356 15564 5408 15570
rect 5172 15506 5224 15512
rect 5276 15524 5356 15552
rect 5184 14958 5212 15506
rect 5276 14958 5304 15524
rect 5356 15506 5408 15512
rect 5552 15094 5580 15846
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5276 14346 5304 14894
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5276 13734 5304 14282
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12714 5212 13126
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5184 12306 5212 12650
rect 5276 12646 5304 13670
rect 5460 13530 5488 14350
rect 5828 14346 5856 14894
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5460 12986 5488 13466
rect 6012 13161 6040 14486
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 13802 6132 14418
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 5998 13152 6054 13161
rect 5622 13084 5918 13104
rect 5998 13087 6054 13096
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5184 11694 5212 12242
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5000 11308 5120 11336
rect 4896 11212 4948 11218
rect 4816 11172 4896 11200
rect 4528 11154 4580 11160
rect 4896 11154 4948 11160
rect 4540 10810 4568 11154
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4816 10198 4844 10542
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4908 9926 4936 11154
rect 5000 10033 5028 11308
rect 5184 11286 5212 11630
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5184 10674 5212 11222
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5276 10606 5304 12582
rect 5540 12300 5592 12306
rect 5460 12260 5540 12288
rect 5460 11694 5488 12260
rect 5540 12242 5592 12248
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11688 5500 11694
rect 5552 11676 5580 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5632 11688 5684 11694
rect 5552 11648 5632 11676
rect 5448 11630 5500 11636
rect 5920 11665 5948 11698
rect 5632 11630 5684 11636
rect 5906 11656 5962 11665
rect 5460 10810 5488 11630
rect 5644 11218 5672 11630
rect 5906 11591 5962 11600
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 4986 10024 5042 10033
rect 5092 9994 5120 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 4986 9959 5042 9968
rect 5080 9988 5132 9994
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4264 8838 4292 9454
rect 4356 9042 4384 9658
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4172 7954 4200 8502
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7546 4200 7890
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4264 5914 4292 8774
rect 4356 8634 4384 8978
rect 4540 8838 4568 9590
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4356 7954 4384 8570
rect 4816 8430 4844 8774
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5000 8378 5028 9959
rect 5080 9930 5132 9936
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 5092 9042 5120 9386
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4632 8090 4660 8366
rect 5000 8350 5120 8378
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4632 7886 4660 8026
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4618 6624 4674 6633
rect 4618 6559 4674 6568
rect 4632 6322 4660 6559
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3436 2145 3464 4966
rect 4356 4826 4384 5714
rect 4908 5166 4936 5850
rect 5000 5778 5028 8230
rect 5092 6798 5120 8350
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6458 5120 6734
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5092 5710 5120 6054
rect 5184 5778 5212 10406
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5276 9926 5304 10066
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 7002 5304 9862
rect 5368 9722 5396 10542
rect 6104 10062 6132 13738
rect 6196 13530 6224 16934
rect 6380 16726 6408 17002
rect 6368 16720 6420 16726
rect 6368 16662 6420 16668
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6472 15978 6500 16594
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 13870 6408 14282
rect 6552 14272 6604 14278
rect 6656 14260 6684 20198
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6748 14414 6776 19110
rect 6840 15706 6868 20742
rect 6932 18970 6960 26590
rect 7208 23662 7236 27526
rect 8114 27520 8170 28000
rect 9402 27520 9458 28000
rect 10690 27520 10746 28000
rect 11978 27520 12034 28000
rect 13266 27520 13322 28000
rect 13912 27532 13964 27538
rect 8128 26654 8156 27520
rect 8116 26648 8168 26654
rect 8116 26590 8168 26596
rect 8760 24268 8812 24274
rect 8760 24210 8812 24216
rect 8772 23866 8800 24210
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7104 23520 7156 23526
rect 7024 23480 7104 23508
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6932 17542 6960 18702
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6840 14958 6868 15506
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14482 6868 14894
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6604 14232 6684 14260
rect 6552 14214 6604 14220
rect 6368 13864 6420 13870
rect 6288 13812 6368 13814
rect 6288 13806 6420 13812
rect 6288 13786 6408 13806
rect 6564 13802 6592 14214
rect 6748 13870 6776 14350
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6552 13796 6604 13802
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6288 12306 6316 13786
rect 6552 13738 6604 13744
rect 6564 13394 6592 13738
rect 6932 13734 6960 17478
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6564 12646 6592 13330
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6288 11898 6316 12242
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6288 11354 6316 11834
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6288 10606 6316 11290
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6104 9722 6132 9998
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 5368 9518 5396 9658
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8566 5396 8978
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5460 8090 5488 8842
rect 5552 8634 5580 9046
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5460 7546 5488 8026
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7546 5580 7890
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5368 6662 5396 6938
rect 6012 6934 6040 7754
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6870
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6104 6322 6132 8502
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6866 6224 7142
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6196 6186 6224 6802
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4896 5160 4948 5166
rect 4526 5128 4582 5137
rect 4896 5102 4948 5108
rect 4526 5063 4582 5072
rect 4540 5030 4568 5063
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4908 4690 4936 4966
rect 5184 4826 5212 5714
rect 5276 5302 5304 5782
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5354 5264 5410 5273
rect 5354 5199 5410 5208
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 4282 4936 4626
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5276 3738 5304 4014
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5368 3602 5396 5199
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 3194 5396 3538
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 2310 3556 2450
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3422 2136 3478 2145
rect 3422 2071 3478 2080
rect 3528 1329 3556 2246
rect 4448 1873 4476 2790
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 4908 2310 4936 2450
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4434 1864 4490 1873
rect 4434 1799 4490 1808
rect 3514 1320 3570 1329
rect 3514 1255 3570 1264
rect 3238 82 3294 480
rect 2976 54 3294 82
rect 662 0 718 54
rect 1950 0 2006 54
rect 3238 0 3294 54
rect 4618 82 4674 480
rect 4908 82 4936 2246
rect 5460 1193 5488 6122
rect 6472 5914 6500 11290
rect 6564 9976 6592 12582
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11898 6684 12174
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6748 11218 6776 12038
rect 7024 11898 7052 23480
rect 7104 23462 7156 23468
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7852 21078 7880 21830
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 7944 20262 7972 21014
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7208 19990 7236 20198
rect 8128 19990 8156 20878
rect 8220 20330 8248 21286
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 7196 19984 7248 19990
rect 7196 19926 7248 19932
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 8208 19984 8260 19990
rect 8312 19972 8340 21422
rect 8260 19944 8340 19972
rect 8208 19926 8260 19932
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 7116 18086 7144 18838
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17814 7144 18022
rect 7104 17808 7156 17814
rect 7104 17750 7156 17756
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 15502 7144 16934
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7116 14074 7144 14418
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7208 13954 7236 19382
rect 7668 19242 7696 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7760 19242 7788 19450
rect 8128 19378 8156 19926
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7668 18426 7696 19178
rect 7760 18970 7788 19178
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7116 13926 7236 13954
rect 7116 12782 7144 13926
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13394 7236 13670
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 12306 7144 12718
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11286 6960 11494
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10470 6776 11154
rect 7116 11014 7144 12242
rect 7208 11218 7236 13330
rect 7300 12442 7328 18022
rect 7760 17814 7788 18022
rect 7852 17882 7880 19110
rect 8128 18970 8156 19314
rect 8220 19174 8248 19926
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 7944 18222 7972 18566
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7760 17066 7788 17750
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7668 16046 7696 16526
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7668 15638 7696 15982
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7392 14958 7420 15506
rect 7576 14958 7604 15506
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12714 7420 13330
rect 7380 12708 7432 12714
rect 7380 12650 7432 12656
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7392 11558 7420 12650
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10606 7144 10950
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6828 10124 6880 10130
rect 7012 10124 7064 10130
rect 6880 10084 7012 10112
rect 6828 10066 6880 10072
rect 7012 10066 7064 10072
rect 6736 9988 6788 9994
rect 6564 9948 6736 9976
rect 6736 9930 6788 9936
rect 6748 9586 6776 9930
rect 6840 9722 6868 10066
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 9178 6776 9522
rect 7116 9518 7144 10542
rect 7208 10266 7236 11154
rect 7392 10674 7420 11494
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6564 7206 6592 7958
rect 6840 7886 6868 8366
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 6390 6592 6598
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6840 6254 6868 7822
rect 6932 7750 6960 8366
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5446 1184 5502 1193
rect 5446 1119 5502 1128
rect 4618 54 4936 82
rect 5552 82 5580 5170
rect 6104 5098 6132 5510
rect 6932 5234 6960 5510
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5644 3738 5672 4150
rect 6012 4010 6040 4966
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5920 3670 5948 3946
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2990 6040 3674
rect 6288 3398 6316 4558
rect 6472 4282 6500 4694
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6932 4146 6960 4694
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6472 3194 6500 3606
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3194 6960 3470
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5644 2553 5672 2926
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5630 2544 5686 2553
rect 5736 2514 5764 2790
rect 7116 2650 7144 9318
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 7546 7236 7890
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7300 6458 7328 8230
rect 7392 7449 7420 9998
rect 7378 7440 7434 7449
rect 7378 7375 7434 7384
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 7002 7420 7210
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7392 5914 7420 6802
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 3670 7236 4082
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7392 3738 7420 3946
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 2582 7236 3470
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 5630 2479 5686 2488
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5906 82 5962 480
rect 5552 54 5962 82
rect 4618 0 4674 54
rect 5906 0 5962 54
rect 7286 82 7342 480
rect 7484 82 7512 14826
rect 7576 14822 7604 14894
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7576 13462 7604 14758
rect 7668 14618 7696 15574
rect 7944 15094 7972 18158
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8128 16454 8156 17138
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 15706 8156 16390
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 8036 13814 8064 14962
rect 8220 14958 8248 18566
rect 8496 18358 8524 18770
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8312 15910 8340 16594
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15065 8340 15846
rect 8298 15056 8354 15065
rect 8298 14991 8354 15000
rect 8208 14952 8260 14958
rect 8128 14912 8208 14940
rect 8128 14346 8156 14912
rect 8208 14894 8260 14900
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7840 13184 7892 13190
rect 7944 13172 7972 13806
rect 8036 13786 8156 13814
rect 7892 13144 7972 13172
rect 7840 13126 7892 13132
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7576 11082 7604 11154
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7576 9994 7604 10542
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9178 7604 9386
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8634 7604 9114
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7546 7604 7890
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 5778 7696 7142
rect 7760 6905 7788 11834
rect 7852 9654 7880 13126
rect 8128 12782 8156 13786
rect 8220 13530 8248 14486
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8024 12300 8076 12306
rect 8128 12288 8156 12718
rect 8076 12260 8156 12288
rect 8024 12242 8076 12248
rect 8220 11694 8248 13466
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12306 8340 12718
rect 8588 12306 8616 19246
rect 8680 17678 8708 23462
rect 8760 22092 8812 22098
rect 8760 22034 8812 22040
rect 8772 21554 8800 22034
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8772 21457 8800 21490
rect 8758 21448 8814 21457
rect 8758 21383 8814 21392
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8772 20466 8800 20742
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8760 20324 8812 20330
rect 8864 20312 8892 21286
rect 8812 20284 8892 20312
rect 8760 20266 8812 20272
rect 8772 19990 8800 20266
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8772 17338 8800 18566
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8680 15910 8708 17002
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13938 8708 14350
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8680 13841 8708 13874
rect 8666 13832 8722 13841
rect 8666 13767 8722 13776
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8312 11898 8340 12242
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8128 11014 8156 11630
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7944 10606 7972 10746
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7944 9450 7972 10542
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 10266 8064 10406
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8312 10130 8340 11834
rect 8680 11762 8708 12582
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8312 9722 8340 10066
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8404 9654 8432 10066
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8220 8294 8248 8978
rect 8404 8430 8432 9454
rect 8496 8906 8524 10950
rect 8680 10470 8708 11290
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 10198 8708 10406
rect 8668 10192 8720 10198
rect 8668 10134 8720 10140
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 7818 8248 8230
rect 8404 7954 8432 8366
rect 8588 8090 8616 8910
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7746 6896 7802 6905
rect 7852 6866 7880 7278
rect 8220 7206 8248 7754
rect 8680 7750 8708 8366
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7746 6831 7802 6840
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 6458 7880 6802
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7944 6390 7972 6598
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5846 7788 6054
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7668 5370 7696 5714
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7760 5302 7788 5782
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 4826 7604 5034
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7576 2961 7604 2994
rect 7562 2952 7618 2961
rect 7562 2887 7618 2896
rect 7760 2650 7788 5238
rect 7944 4690 7972 6326
rect 8128 6322 8156 6734
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7944 4146 7972 4626
rect 8116 4548 8168 4554
rect 8220 4536 8248 7142
rect 8680 6934 8708 7686
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8668 6928 8720 6934
rect 8668 6870 8720 6876
rect 8312 4690 8340 6870
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8168 4508 8248 4536
rect 8116 4490 8168 4496
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8128 3942 8156 4490
rect 8588 4214 8616 4626
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8772 4154 8800 17138
rect 8864 13870 8892 18294
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8944 15972 8996 15978
rect 8944 15914 8996 15920
rect 8956 15570 8984 15914
rect 9048 15706 9076 16050
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9140 15638 9168 19110
rect 9232 18290 9260 24006
rect 9416 22778 9444 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 23866 10732 27520
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 23322 9904 23598
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 10152 22438 10180 23122
rect 11992 22778 12020 27520
rect 13280 24177 13308 27520
rect 14554 27532 14610 28000
rect 14554 27520 14556 27532
rect 13912 27474 13964 27480
rect 14608 27520 14610 27532
rect 15750 27520 15806 28000
rect 17038 27520 17094 28000
rect 18326 27554 18382 28000
rect 19614 27554 19670 28000
rect 17144 27526 17356 27554
rect 17144 27520 17172 27526
rect 14556 27474 14608 27480
rect 13266 24168 13322 24177
rect 13266 24103 13322 24112
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 9508 22234 9536 22374
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9784 21690 9812 22374
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9680 21412 9732 21418
rect 9680 21354 9732 21360
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9508 18902 9536 19382
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9312 18692 9364 18698
rect 9312 18634 9364 18640
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9232 17882 9260 18226
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9324 17762 9352 18634
rect 9508 18222 9536 18838
rect 9692 18426 9720 21354
rect 9772 21344 9824 21350
rect 9876 21332 9904 22034
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9824 21304 9904 21332
rect 9772 21286 9824 21292
rect 9784 19990 9812 21286
rect 9968 20602 9996 21830
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 9968 20262 9996 20538
rect 10060 20466 10088 21082
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 10152 20346 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10692 21548 10744 21554
rect 10796 21536 10824 21830
rect 10744 21508 10824 21536
rect 10692 21490 10744 21496
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 10336 20942 10364 21014
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10244 20466 10272 20878
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10060 20318 10180 20346
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9784 18630 9812 19926
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9968 19378 9996 19790
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18698 9996 19178
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9232 17734 9352 17762
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 8852 13864 8904 13870
rect 8904 13812 8984 13814
rect 8852 13806 8984 13812
rect 8864 13786 8984 13806
rect 8956 12782 8984 13786
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 13530 9076 13738
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8864 6225 8892 12378
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8956 10674 8984 12242
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11558 9076 12038
rect 9140 11626 9168 13874
rect 9232 13716 9260 17734
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 17338 9628 17614
rect 9876 17338 9904 17750
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9416 15706 9444 16662
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9508 13938 9536 16526
rect 9968 16182 9996 16730
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9968 15910 9996 16118
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15706 9996 15846
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 9876 14618 9904 15506
rect 9968 15094 9996 15642
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9968 14822 9996 15030
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14618 9996 14758
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9508 13809 9536 13874
rect 9232 13688 9352 13716
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11082 9076 11494
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8956 7342 8984 10610
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 10266 9076 10474
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9140 10130 9168 11562
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9140 9178 9168 9386
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9048 7478 9076 8026
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8956 6662 8984 7278
rect 9048 7002 9076 7414
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 9048 6322 9076 6666
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8850 6216 8906 6225
rect 8850 6151 8906 6160
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5846 8984 6054
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9048 5778 9076 6258
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8680 4126 8800 4154
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7852 3058 7880 3402
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 8128 1737 8156 3878
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 2922 8340 3470
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8588 2514 8616 2790
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8114 1728 8170 1737
rect 8114 1663 8170 1672
rect 7286 54 7512 82
rect 8574 82 8630 480
rect 8680 82 8708 4126
rect 8758 4040 8814 4049
rect 8758 3975 8814 3984
rect 8772 3602 8800 3975
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3058 8800 3538
rect 8956 3233 8984 4966
rect 9232 4282 9260 5782
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9232 3942 9260 4218
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3670 9260 3878
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 8942 3224 8998 3233
rect 9232 3194 9260 3606
rect 8942 3159 8998 3168
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2650 8800 2790
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 9324 2310 9352 13688
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9508 13025 9536 13330
rect 9494 13016 9550 13025
rect 9494 12951 9550 12960
rect 9508 12850 9536 12951
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9784 12646 9812 14350
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 13258 9996 13330
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9968 12442 9996 13194
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11626 9720 12038
rect 10060 11762 10088 20318
rect 10336 20244 10364 20878
rect 10704 20330 10732 21286
rect 10796 20505 10824 21508
rect 10876 21548 10928 21554
rect 10876 21490 10928 21496
rect 10888 21078 10916 21490
rect 11256 21350 11284 22034
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 11716 20992 11744 21354
rect 11796 21004 11848 21010
rect 11716 20964 11796 20992
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20602 11100 20878
rect 11716 20602 11744 20964
rect 11796 20946 11848 20952
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 10782 20496 10838 20505
rect 10782 20431 10838 20440
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10152 20216 10364 20244
rect 10152 19514 10180 20216
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 19990 10732 20266
rect 11716 20058 11744 20538
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 13096 19990 13124 20198
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10152 19174 10180 19450
rect 11440 19174 11468 19722
rect 11624 19242 11652 19926
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10888 18902 10916 19110
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17678 10732 18090
rect 10888 18086 10916 18838
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10796 17814 10824 18022
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16250 10732 17002
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10704 15910 10732 16186
rect 10796 15978 10824 16390
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 10152 14958 10180 15370
rect 10796 15162 10824 15914
rect 10888 15366 10916 18022
rect 11072 17882 11100 18022
rect 11164 17882 11192 18702
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11072 17202 11100 17818
rect 11256 17678 11284 18702
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10980 15706 11008 16050
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14550 10180 14894
rect 10888 14890 10916 15302
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10140 13728 10192 13734
rect 10244 13716 10272 14486
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10192 13688 10272 13716
rect 10140 13670 10192 13676
rect 10152 12646 10180 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13874
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 12306 10180 12582
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9600 11014 9628 11562
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9692 10792 9720 11562
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9784 10810 9812 11222
rect 10060 11150 10088 11698
rect 10152 11558 10180 12242
rect 10336 12209 10364 12310
rect 10876 12232 10928 12238
rect 10322 12200 10378 12209
rect 10876 12174 10928 12180
rect 10322 12135 10378 12144
rect 10888 11898 10916 12174
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9600 10764 9720 10792
rect 9772 10804 9824 10810
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9416 10266 9444 10542
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9508 8566 9536 10542
rect 9600 10470 9628 10764
rect 9772 10746 9824 10752
rect 9678 10704 9734 10713
rect 9678 10639 9734 10648
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 9926 9628 10406
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9692 9586 9720 10639
rect 10152 10538 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10980 11098 11008 15642
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13462 11192 14214
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11256 13326 11284 17614
rect 11440 16998 11468 19110
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11716 16114 11744 19790
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12268 18426 12296 19110
rect 13096 18970 13124 19926
rect 13280 19514 13308 19926
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13372 19378 13400 19790
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13372 18873 13400 19110
rect 13740 18970 13768 19654
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13820 18896 13872 18902
rect 13358 18864 13414 18873
rect 12624 18828 12676 18834
rect 13820 18838 13872 18844
rect 13358 18799 13414 18808
rect 12624 18770 12676 18776
rect 12636 18426 12664 18770
rect 13452 18760 13504 18766
rect 13450 18728 13452 18737
rect 13504 18728 13506 18737
rect 13450 18663 13506 18672
rect 13464 18630 13492 18663
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 11808 18329 11836 18362
rect 11794 18320 11850 18329
rect 11794 18255 11850 18264
rect 11808 18222 11836 18255
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 12636 18086 12664 18362
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11808 16998 11836 17750
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 17202 12020 17546
rect 11980 17196 12032 17202
rect 11900 17156 11980 17184
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11808 16794 11836 16934
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14618 11376 14758
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11624 14550 11652 15438
rect 11716 15434 11744 16050
rect 11808 15638 11836 16730
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11808 15162 11836 15574
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11900 15094 11928 17156
rect 11980 17138 12032 17144
rect 12268 17066 12296 17614
rect 12636 17241 12664 18022
rect 13556 17882 13584 18022
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13648 17610 13676 18294
rect 13740 17814 13768 18566
rect 13832 18086 13860 18838
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 12622 17232 12678 17241
rect 12622 17167 12678 17176
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16726 12940 16934
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 16250 12204 16526
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12268 16114 12296 16662
rect 13188 16454 13216 17070
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11900 14414 11928 15030
rect 12360 15026 12388 15982
rect 13188 15706 13216 16390
rect 13372 16182 13400 16934
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13372 15978 13400 16118
rect 13464 16114 13492 16390
rect 13648 16114 13676 17002
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13740 16250 13768 16662
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13268 15564 13320 15570
rect 13820 15564 13872 15570
rect 13268 15506 13320 15512
rect 13740 15524 13820 15552
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12728 15026 12756 15302
rect 13280 15162 13308 15506
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 10704 11070 11008 11098
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 11070
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9862 9480 9918 9489
rect 9862 9415 9918 9424
rect 9876 9178 9904 9415
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9784 8294 9812 8978
rect 9876 8906 9904 9114
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 10152 8838 10180 10066
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8498 10180 8774
rect 10704 8537 10732 10202
rect 10796 8922 10824 10950
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9178 10916 9998
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10796 8894 10916 8922
rect 10690 8528 10746 8537
rect 10140 8492 10192 8498
rect 10690 8463 10746 8472
rect 10140 8434 10192 8440
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8090 9812 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9692 7546 9720 7890
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9968 7342 9996 7890
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6390 9536 6802
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9784 5234 9812 6938
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10152 6458 10180 6802
rect 10704 6798 10732 8463
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9784 4826 9812 5170
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4758 9904 5782
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9968 5370 9996 5646
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3738 9628 4082
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9772 3664 9824 3670
rect 9876 3652 9904 4694
rect 10060 4690 10088 6122
rect 10152 5710 10180 6258
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5234 10180 5646
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4758 10732 5102
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 4282 10548 4558
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10060 3670 10088 3946
rect 9824 3624 9904 3652
rect 10048 3664 10100 3670
rect 9772 3606 9824 3612
rect 10048 3606 10100 3612
rect 9784 3194 9812 3606
rect 10152 3466 10180 3946
rect 10704 3942 10732 4694
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10796 4049 10824 4558
rect 10888 4154 10916 8894
rect 10980 8498 11008 10406
rect 11072 10198 11100 10474
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11072 8974 11100 9454
rect 11164 9042 11192 9522
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11072 7342 11100 8910
rect 11164 8090 11192 8978
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11348 7342 11376 7686
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11072 7002 11100 7278
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11348 5710 11376 7278
rect 11440 6610 11468 13126
rect 11532 12442 11560 13262
rect 11624 12986 11652 13670
rect 11716 13258 11744 14282
rect 11900 13938 11928 14350
rect 11992 14074 12020 14486
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11808 12986 11836 13398
rect 12636 12986 12664 14214
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12164 12776 12216 12782
rect 12162 12744 12164 12753
rect 12216 12744 12218 12753
rect 12162 12679 12218 12688
rect 12346 12744 12402 12753
rect 12346 12679 12402 12688
rect 12176 12646 12204 12679
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 12360 11830 12388 12679
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12452 11286 12480 11494
rect 12440 11280 12492 11286
rect 12360 11240 12440 11268
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 10470 12020 11154
rect 12070 10568 12126 10577
rect 12070 10503 12126 10512
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 11624 9586 11652 10134
rect 11992 9625 12020 10406
rect 12084 10130 12112 10503
rect 12360 10470 12388 11240
rect 12440 11222 12492 11228
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12544 10674 12572 11086
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 11978 9616 12034 9625
rect 11612 9580 11664 9586
rect 11978 9551 12034 9560
rect 11612 9522 11664 9528
rect 11624 9110 11652 9522
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11624 8634 11652 9046
rect 12360 9042 12388 10406
rect 12438 10024 12494 10033
rect 12438 9959 12494 9968
rect 12452 9926 12480 9959
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 9178 12572 9318
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11624 7886 11652 8570
rect 12360 8362 12388 8978
rect 12636 8974 12664 10950
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8537 12572 8774
rect 12530 8528 12586 8537
rect 12530 8463 12586 8472
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 8090 12572 8230
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11624 7546 11652 7822
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7313 11652 7346
rect 11610 7304 11666 7313
rect 11520 7268 11572 7274
rect 11610 7239 11666 7248
rect 11520 7210 11572 7216
rect 11532 6730 11560 7210
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11440 6582 11652 6610
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10888 4126 11008 4154
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 3126 9904 3334
rect 10704 3194 10732 3470
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10152 2446 10180 3062
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10704 2650 10732 3130
rect 10980 3126 11008 4126
rect 11336 3936 11388 3942
rect 11388 3896 11468 3924
rect 11336 3878 11388 3884
rect 11440 3670 11468 3896
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11440 3194 11468 3606
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 11532 3058 11560 4966
rect 11624 3194 11652 6582
rect 11716 5914 11744 6870
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11808 6322 11836 6802
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11900 5846 11928 7482
rect 12636 7274 12664 7890
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11900 5302 11928 5782
rect 12084 5778 12112 6734
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5370 12112 5714
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 12268 4826 12296 6054
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 12636 4826 12664 5238
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4146 11928 4422
rect 12636 4282 12664 4762
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12636 4010 12664 4218
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3738 12664 3946
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12530 3632 12586 3641
rect 12530 3567 12586 3576
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11716 3058 11744 3470
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11716 2961 11744 2994
rect 11702 2952 11758 2961
rect 11520 2916 11572 2922
rect 11702 2887 11758 2896
rect 11520 2858 11572 2864
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 11532 2514 11560 2858
rect 11794 2544 11850 2553
rect 11520 2508 11572 2514
rect 11794 2479 11850 2488
rect 11520 2450 11572 2456
rect 11808 2446 11836 2479
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 9876 2310 9904 2382
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 8574 54 8708 82
rect 9954 82 10010 480
rect 10060 82 10088 2314
rect 11334 1320 11390 1329
rect 11334 1255 11390 1264
rect 9954 54 10088 82
rect 11242 82 11298 480
rect 11348 82 11376 1255
rect 11242 54 11376 82
rect 12544 82 12572 3567
rect 12728 3466 12756 14962
rect 13464 14550 13492 15370
rect 13740 15026 13768 15524
rect 13820 15506 13872 15512
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 13530 12848 13738
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13188 13462 13216 13874
rect 13464 13530 13492 14486
rect 13648 14346 13676 14758
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12912 12306 12940 12650
rect 13096 12442 13124 13262
rect 13188 12986 13216 13398
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12912 11898 12940 12242
rect 13648 12186 13676 14282
rect 13740 14278 13768 14962
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13832 14074 13860 14486
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13740 13462 13768 13738
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13740 12850 13768 13398
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13464 12158 13676 12186
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10538 12848 10950
rect 13188 10538 13216 11018
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 12820 10198 12848 10474
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12820 9110 12848 10134
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9518 12940 9862
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13082 9480 13138 9489
rect 13082 9415 13138 9424
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8090 13032 8910
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6254 12940 6802
rect 13004 6662 13032 7346
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 13004 5914 13032 6598
rect 13096 6186 13124 9415
rect 13188 9178 13216 10474
rect 13372 10198 13400 11562
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13358 10024 13414 10033
rect 13358 9959 13414 9968
rect 13266 9616 13322 9625
rect 13372 9586 13400 9959
rect 13266 9551 13322 9560
rect 13360 9580 13412 9586
rect 13280 9518 13308 9551
rect 13360 9522 13412 9528
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13188 7410 13216 9114
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8498 13308 8910
rect 13372 8498 13400 9522
rect 13464 9489 13492 12158
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11762 13584 12038
rect 13832 11898 13860 12310
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 10169 13584 11698
rect 13820 11212 13872 11218
rect 13924 11200 13952 27474
rect 14568 27443 14596 27474
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15764 23866 15792 27520
rect 17052 27492 17172 27520
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21049 15332 23462
rect 15290 21040 15346 21049
rect 15290 20975 15346 20984
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 14016 18970 14044 19178
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14016 17814 14044 18906
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 14016 17270 14044 17750
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13872 11172 13952 11200
rect 13820 11154 13872 11160
rect 13832 10470 13860 11154
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13542 10160 13598 10169
rect 13542 10095 13598 10104
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13450 9480 13506 9489
rect 13556 9450 13584 9930
rect 13450 9415 13506 9424
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9110 13492 9318
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8634 13492 9046
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13556 8566 13584 9386
rect 13648 9042 13676 10066
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13740 8974 13768 9998
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13544 8560 13596 8566
rect 13450 8528 13506 8537
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13360 8492 13412 8498
rect 13544 8502 13596 8508
rect 13450 8463 13506 8472
rect 13360 8434 13412 8440
rect 13280 7818 13308 8434
rect 13464 8430 13492 8463
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13556 8362 13584 8502
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13464 6866 13492 7686
rect 13648 7546 13676 7822
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13464 6390 13492 6802
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13464 6118 13492 6326
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12806 4040 12862 4049
rect 12900 4004 12952 4010
rect 12862 3984 12900 3992
rect 12806 3975 12900 3984
rect 12820 3964 12900 3975
rect 12900 3946 12952 3952
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3670 13400 3878
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12912 3058 12940 3606
rect 13372 3194 13400 3606
rect 13464 3194 13492 6054
rect 13648 4282 13676 6734
rect 13832 5896 13860 10406
rect 13924 10033 13952 10474
rect 13910 10024 13966 10033
rect 13910 9959 13966 9968
rect 13924 9926 13952 9959
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13924 8974 13952 9046
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13740 5868 13860 5896
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 4154 13768 5868
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13832 5370 13860 5714
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13832 5273 13860 5306
rect 13818 5264 13874 5273
rect 13818 5199 13874 5208
rect 14016 4690 14044 17070
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14200 16454 14228 16662
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14200 15978 14228 16390
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14108 15162 14136 15914
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14292 13814 14320 20538
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14384 18902 14412 19178
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14464 18148 14516 18154
rect 14464 18090 14516 18096
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14476 17814 14504 18090
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14568 17338 14596 18090
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14384 16046 14412 17206
rect 14660 16794 14688 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14752 16726 14780 18226
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14752 15978 14780 16662
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14200 13786 14320 13814
rect 14200 12753 14228 13786
rect 14186 12744 14242 12753
rect 14186 12679 14242 12688
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14292 12170 14320 12650
rect 14384 12238 14412 12650
rect 14844 12306 14872 18362
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17134 15332 20975
rect 16500 18902 16528 23462
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15488 18426 15516 18770
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 16040 18290 16068 18702
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15396 16998 15424 17682
rect 15580 16998 15608 17682
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15609 15148 15982
rect 15106 15600 15162 15609
rect 15106 15535 15162 15544
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10606 14228 10950
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14108 9625 14136 10202
rect 14292 10033 14320 12106
rect 14384 11898 14412 12174
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11898 15332 12242
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 10713 14504 11630
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14462 10704 14518 10713
rect 14462 10639 14518 10648
rect 14556 10532 14608 10538
rect 14556 10474 14608 10480
rect 14278 10024 14334 10033
rect 14278 9959 14334 9968
rect 14094 9616 14150 9625
rect 14094 9551 14150 9560
rect 14108 8294 14136 9551
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 8838 14228 9454
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 14200 8090 14228 8366
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14108 7256 14136 7958
rect 14188 7268 14240 7274
rect 14108 7228 14188 7256
rect 14108 7002 14136 7228
rect 14188 7210 14240 7216
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14200 5098 14228 5578
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4826 14228 5034
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 13648 4126 13768 4154
rect 13648 4078 13676 4126
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13648 2514 13676 4014
rect 14016 3942 14044 4626
rect 14372 4548 14424 4554
rect 14372 4490 14424 4496
rect 14384 4010 14412 4490
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14016 3233 14044 3878
rect 14200 3738 14228 3878
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14292 3602 14320 3946
rect 14384 3738 14412 3946
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14568 3641 14596 10474
rect 14752 9722 14780 11290
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10266 15424 16934
rect 15580 15026 15608 16934
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15672 15910 15700 16662
rect 15764 16454 15792 18022
rect 15934 17776 15990 17785
rect 15934 17711 15990 17720
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 16658 15884 17614
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15638 15700 15846
rect 15856 15706 15884 16594
rect 15948 16250 15976 17711
rect 16316 17202 16344 18226
rect 16500 17882 16528 18838
rect 16592 18086 16620 18838
rect 17328 18329 17356 27526
rect 17972 27526 18382 27554
rect 17408 23656 17460 23662
rect 17406 23624 17408 23633
rect 17500 23656 17552 23662
rect 17460 23624 17462 23633
rect 17500 23598 17552 23604
rect 17406 23559 17462 23568
rect 17420 23526 17448 23559
rect 17408 23520 17460 23526
rect 17408 23462 17460 23468
rect 17512 20602 17540 23598
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17314 18320 17370 18329
rect 17314 18255 17370 18264
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16316 15978 16344 16526
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 15672 15162 15700 15574
rect 16408 15162 16436 17002
rect 16960 16454 16988 17002
rect 17696 16590 17724 18702
rect 17972 17785 18000 27526
rect 18326 27520 18382 27526
rect 19352 27526 19670 27554
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18340 20505 18368 20742
rect 18326 20496 18382 20505
rect 18326 20431 18382 20440
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 17958 17776 18014 17785
rect 17958 17711 18014 17720
rect 18616 17649 18644 18022
rect 18602 17640 18658 17649
rect 18602 17575 18658 17584
rect 19352 17105 19380 27526
rect 19614 27520 19670 27526
rect 20902 27520 20958 28000
rect 22098 27520 22154 28000
rect 23386 27520 23442 28000
rect 24674 27520 24730 28000
rect 24860 27532 24912 27538
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19430 24168 19486 24177
rect 19430 24103 19486 24112
rect 19444 23594 19472 24103
rect 20916 23866 20944 27520
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19444 18426 19472 23530
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16960 16114 16988 16390
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15672 14872 15700 15098
rect 15934 15056 15990 15065
rect 15934 14991 15936 15000
rect 15988 14991 15990 15000
rect 15936 14962 15988 14968
rect 15752 14884 15804 14890
rect 15672 14844 15752 14872
rect 15672 14532 15700 14844
rect 15752 14826 15804 14832
rect 15752 14544 15804 14550
rect 15672 14504 15752 14532
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15580 13841 15608 14010
rect 15672 14006 15700 14504
rect 15752 14486 15804 14492
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15566 13832 15622 13841
rect 15566 13767 15622 13776
rect 15580 13394 15608 13767
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12986 15608 13330
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 12918 15700 13942
rect 15948 13870 15976 14962
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15856 12782 15884 13330
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 12102 15884 12718
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11694 15884 12038
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15580 11354 15608 11630
rect 15856 11558 15884 11630
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15580 10198 15608 10542
rect 15764 10538 15792 11154
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15488 9722 15516 10134
rect 15672 9722 15700 10406
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15672 9382 15700 9658
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 14660 7478 14688 9046
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15488 8634 15516 9046
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15856 8430 15884 11494
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15474 8256 15530 8265
rect 15474 8191 15530 8200
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 15304 7410 15332 7890
rect 15488 7750 15516 8191
rect 15856 8022 15884 8366
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15948 7818 15976 13806
rect 16132 13394 16160 14214
rect 16500 13870 16528 14894
rect 16592 14482 16620 15846
rect 17696 15638 17724 16526
rect 17788 16250 17816 16662
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17788 15706 17816 16186
rect 18052 16176 18104 16182
rect 18052 16118 18104 16124
rect 18064 15706 18092 16118
rect 18524 16046 18552 16390
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 16868 14550 16896 15438
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16868 13938 16896 14486
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17420 14074 17448 14418
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16500 13530 16528 13806
rect 17512 13682 17540 15098
rect 17880 14890 17908 15438
rect 17972 15162 18000 15506
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17420 13654 17540 13682
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 17316 13456 17368 13462
rect 17316 13398 17368 13404
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16224 12442 16252 12786
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16316 12306 16344 13262
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 16224 10130 16252 11562
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9654 16068 9998
rect 16028 9648 16080 9654
rect 16080 9608 16160 9636
rect 16028 9590 16080 9596
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 16040 9178 16068 9386
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16132 9042 16160 9608
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16408 8265 16436 12922
rect 17328 12714 17356 13398
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 16776 12356 16804 12650
rect 16856 12368 16908 12374
rect 16776 12328 16856 12356
rect 16776 11898 16804 12328
rect 16856 12310 16908 12316
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16960 11898 16988 12242
rect 16764 11892 16816 11898
rect 16948 11892 17000 11898
rect 16816 11852 16896 11880
rect 16764 11834 16816 11840
rect 16868 11286 16896 11852
rect 16948 11834 17000 11840
rect 17420 11762 17448 13654
rect 17604 12850 17632 14554
rect 17880 14482 17908 14826
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 13870 17908 14418
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 18156 13326 18184 14758
rect 18524 14550 18552 14894
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18524 14278 18552 14486
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13530 18276 13670
rect 18524 13530 18552 13738
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18156 12986 18184 13262
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18248 12306 18276 12650
rect 18340 12442 18368 12650
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10674 16528 10950
rect 16776 10674 16804 11086
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16500 10266 16528 10610
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16394 8256 16450 8265
rect 16394 8191 16450 8200
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15476 7744 15528 7750
rect 15396 7704 15476 7732
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 6254 14872 6802
rect 14936 6730 14964 7346
rect 15304 7313 15332 7346
rect 15290 7304 15346 7313
rect 15290 7239 15346 7248
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6322 15424 7704
rect 15476 7686 15528 7692
rect 16316 7274 16344 7958
rect 16500 7954 16528 8910
rect 16776 8498 16804 10610
rect 16868 10470 16896 11222
rect 18064 11014 18092 11630
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17696 10538 17724 10950
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10180 16896 10406
rect 17696 10198 17724 10474
rect 16948 10192 17000 10198
rect 16868 10152 16948 10180
rect 16868 9722 16896 10152
rect 16948 10134 17000 10140
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17788 9926 17816 10746
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9722 17816 9862
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 9382 17816 9658
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 18064 9110 18092 10950
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9450 18184 9862
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18156 9178 18184 9386
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17040 8560 17092 8566
rect 17144 8537 17172 8978
rect 17328 8634 17356 8978
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17040 8502 17092 8508
rect 17130 8528 17186 8537
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 15580 6934 15608 7210
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15488 6458 15516 6734
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5914 14872 6190
rect 15476 6112 15528 6118
rect 15580 6100 15608 6870
rect 15764 6662 15792 7142
rect 16500 7002 16528 7890
rect 16960 7818 16988 8502
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 17052 7478 17080 8502
rect 17130 8463 17186 8472
rect 17144 8276 17172 8463
rect 17328 8430 17356 8570
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17420 8362 17448 8978
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17224 8288 17276 8294
rect 17144 8248 17224 8276
rect 17224 8230 17276 8236
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15528 6072 15608 6100
rect 15476 6054 15528 6060
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 5234 14780 5510
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4010 14780 5034
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14752 3670 14780 3946
rect 14844 3738 14872 5850
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5370 15424 5782
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14740 3664 14792 3670
rect 14554 3632 14610 3641
rect 14280 3596 14332 3602
rect 14740 3606 14792 3612
rect 14554 3567 14610 3576
rect 14280 3538 14332 3544
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14002 3224 14058 3233
rect 14956 3216 15252 3236
rect 14002 3159 14058 3168
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 12622 82 12678 480
rect 12544 54 12678 82
rect 13740 82 13768 3062
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14568 2854 14596 2926
rect 15304 2854 15332 5102
rect 15488 5030 15516 6054
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 5137 15608 5646
rect 15566 5128 15622 5137
rect 15566 5063 15622 5072
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4758 15516 4966
rect 15580 4826 15608 5063
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 4214 15424 4558
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15396 3738 15424 4150
rect 15488 3942 15516 4694
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15488 2990 15516 3606
rect 15568 3596 15620 3602
rect 15672 3584 15700 6122
rect 15764 5846 15792 6598
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15948 5914 15976 6190
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4282 16344 4422
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16316 4010 16344 4218
rect 16500 4146 16528 5714
rect 17144 5098 17172 5782
rect 17132 5092 17184 5098
rect 17132 5034 17184 5040
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4758 16896 4966
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 15620 3556 15700 3584
rect 15568 3538 15620 3544
rect 15580 3194 15608 3538
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 14568 2446 14596 2790
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 13910 82 13966 480
rect 14384 134 14412 2246
rect 14568 2106 14596 2382
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 13740 54 13966 82
rect 14372 128 14424 134
rect 14372 70 14424 76
rect 15290 82 15346 480
rect 15396 82 15424 2858
rect 16224 2514 16252 3946
rect 16500 3738 16528 4082
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 17132 3596 17184 3602
rect 17236 3584 17264 8230
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17604 7177 17632 7278
rect 17590 7168 17646 7177
rect 17590 7103 17646 7112
rect 17880 6866 17908 8570
rect 18156 8498 18184 8774
rect 18248 8634 18276 9046
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18616 8634 18644 8978
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7886 18184 8230
rect 18248 8004 18276 8298
rect 18328 8016 18380 8022
rect 18248 7976 18328 8004
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18248 7750 18276 7976
rect 18328 7958 18380 7964
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7478 18276 7686
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 18156 6730 18184 7210
rect 18248 6934 18276 7414
rect 18340 7274 18368 7822
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18236 6928 18288 6934
rect 18340 6905 18368 7210
rect 18432 7206 18460 7346
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18510 7168 18566 7177
rect 18510 7103 18566 7112
rect 18524 7002 18552 7103
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18236 6870 18288 6876
rect 18326 6896 18382 6905
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5030 17632 5646
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 4282 17448 4694
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17604 3670 17632 4966
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 4146 17724 4558
rect 17788 4282 17816 6054
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17972 3738 18000 4490
rect 18156 4010 18184 6258
rect 18248 5914 18276 6870
rect 18326 6831 18382 6840
rect 18616 6730 18644 7346
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18340 4758 18368 6122
rect 18616 5846 18644 6122
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18616 5574 18644 5782
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18616 5098 18644 5510
rect 18708 5234 18736 8502
rect 18800 7970 18828 15914
rect 19352 14618 19380 17031
rect 19444 15026 19472 18362
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 22112 15162 22140 27520
rect 23400 23866 23428 27520
rect 23754 26616 23810 26625
rect 23754 26551 23810 26560
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22848 20602 22876 20946
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 19982 14512 20038 14521
rect 19800 14476 19852 14482
rect 19982 14447 20038 14456
rect 19800 14418 19852 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18892 12850 18920 13874
rect 19352 13734 19380 14282
rect 19812 14074 19840 14418
rect 19996 14074 20024 14447
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19984 13864 20036 13870
rect 20088 13852 20116 14214
rect 20036 13824 20116 13852
rect 19984 13806 20036 13812
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19168 12646 19196 13398
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12714 19472 13126
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11830 18920 12174
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18892 11665 18920 11766
rect 18878 11656 18934 11665
rect 19168 11626 19196 12378
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 18878 11591 18934 11600
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 11286 19012 11494
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10674 19104 11086
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 19168 10538 19196 11222
rect 19352 11150 19380 12242
rect 19444 11540 19472 12650
rect 19536 12646 19564 13262
rect 19892 12912 19944 12918
rect 19892 12854 19944 12860
rect 19904 12714 19932 12854
rect 20088 12850 20116 13824
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19892 12708 19944 12714
rect 20076 12708 20128 12714
rect 19944 12668 20024 12696
rect 19892 12650 19944 12656
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19536 12209 19564 12582
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19996 12442 20024 12668
rect 20076 12650 20128 12656
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19522 12200 19578 12209
rect 19522 12135 19578 12144
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11898 19840 12038
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19524 11552 19576 11558
rect 19444 11512 19524 11540
rect 19524 11494 19576 11500
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18892 8090 18920 9998
rect 19076 9926 19104 10474
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19168 9722 19196 10134
rect 19352 10062 19380 11086
rect 19536 10742 19564 11494
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19892 11008 19944 11014
rect 19996 10996 20024 11562
rect 20088 11286 20116 12650
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19944 10968 20024 10996
rect 19892 10950 19944 10956
rect 19904 10810 19932 10950
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 20088 10742 20116 11222
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19352 9586 19380 9998
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 9722 19932 9862
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19340 8832 19392 8838
rect 19444 8820 19472 9522
rect 19984 9512 20036 9518
rect 20036 9472 20116 9500
rect 19984 9454 20036 9460
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 8906 19564 9318
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19392 8792 19472 8820
rect 19340 8774 19392 8780
rect 19352 8294 19380 8774
rect 20088 8430 20116 9472
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19340 8288 19392 8294
rect 19444 8265 19472 8298
rect 19524 8288 19576 8294
rect 19340 8230 19392 8236
rect 19430 8256 19486 8265
rect 19524 8230 19576 8236
rect 19430 8191 19486 8200
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 19536 8022 19564 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19524 8016 19576 8022
rect 18800 7942 19104 7970
rect 19524 7958 19576 7964
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18800 6730 18828 7210
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18800 6322 18828 6666
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18970 6216 19026 6225
rect 18970 6151 19026 6160
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18524 4826 18552 5034
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18248 4010 18276 4218
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18156 3738 18184 3946
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 18432 3602 18460 4082
rect 18524 4049 18552 4762
rect 18708 4554 18736 5170
rect 18696 4548 18748 4554
rect 18696 4490 18748 4496
rect 18510 4040 18566 4049
rect 18510 3975 18566 3984
rect 17184 3556 17264 3584
rect 17408 3596 17460 3602
rect 17132 3538 17184 3544
rect 17408 3538 17460 3544
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 17144 3194 17172 3538
rect 17420 3194 17448 3538
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17512 2990 17540 3334
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 7286 0 7342 54
rect 8574 0 8630 54
rect 9954 0 10010 54
rect 11242 0 11298 54
rect 12622 0 12678 54
rect 13910 0 13966 54
rect 15290 54 15424 82
rect 16578 82 16634 480
rect 16776 82 16804 2790
rect 17512 2582 17540 2926
rect 18156 2650 18184 3402
rect 18432 3194 18460 3538
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 16578 54 16804 82
rect 17696 82 17724 2586
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 18892 2446 18920 2479
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 17958 82 18014 480
rect 17696 54 18014 82
rect 18984 82 19012 6151
rect 19076 2582 19104 7942
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6458 19288 6734
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19536 5846 19564 7822
rect 20088 7818 20116 8366
rect 20180 8090 20208 8978
rect 20272 8430 20300 14554
rect 20916 13433 20944 14758
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21100 14074 21128 14418
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13814 21128 14010
rect 21376 13938 21404 14758
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21100 13802 21312 13814
rect 21100 13796 21324 13802
rect 21100 13786 21272 13796
rect 21100 13530 21128 13786
rect 21272 13738 21324 13744
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20902 13424 20958 13433
rect 20902 13359 20958 13368
rect 20916 12306 20944 13359
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11762 20392 12038
rect 20916 11830 20944 12242
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11354 20392 11698
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10538 20760 10746
rect 21008 10742 21036 11086
rect 21100 10810 21128 11222
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20640 9926 20668 10474
rect 21100 10198 21128 10746
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20904 10124 20956 10130
rect 21192 10112 21220 13670
rect 21376 13530 21404 13874
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21560 12850 21588 13398
rect 21744 13326 21772 13670
rect 21836 13462 21864 14350
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21560 11082 21588 12786
rect 21744 12442 21772 13262
rect 21836 12986 21864 13398
rect 22020 13326 22048 13738
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22008 13320 22060 13326
rect 22388 13297 22416 13330
rect 22008 13262 22060 13268
rect 22374 13288 22430 13297
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 21836 11898 21864 12310
rect 22020 12238 22048 13262
rect 22374 13223 22430 13232
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22020 11898 22048 12174
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 21836 11218 21864 11834
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22112 11354 22140 11698
rect 22756 11626 22784 12174
rect 22848 11762 22876 12174
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22204 11286 22232 11562
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21560 10606 21588 11018
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 22296 10169 22324 11494
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22572 10810 22600 11154
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22756 10606 22784 11562
rect 22940 10742 22968 23462
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23400 12986 23428 13330
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 23676 10266 23704 22510
rect 23768 12782 23796 26551
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21010 24716 27520
rect 25962 27532 26018 28000
rect 25962 27520 25964 27532
rect 24860 27474 24912 27480
rect 26016 27520 26018 27532
rect 27250 27520 27306 28000
rect 25964 27474 26016 27480
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 24780 22778 24808 23423
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24122 18320 24178 18329
rect 24122 18255 24178 18264
rect 24136 16658 24164 18255
rect 24214 17776 24270 17785
rect 24214 17711 24270 17720
rect 24228 17134 24256 17711
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24766 17368 24822 17377
rect 24766 17303 24822 17312
rect 24780 17270 24808 17303
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24136 16250 24164 16594
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24872 13814 24900 27474
rect 25976 27443 26004 27474
rect 25134 25120 25190 25129
rect 25134 25055 25190 25064
rect 25148 23866 25176 25055
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23662 25176 23802
rect 25136 23656 25188 23662
rect 27264 23633 27292 27520
rect 25136 23598 25188 23604
rect 27250 23624 27306 23633
rect 27250 23559 27306 23568
rect 27618 22536 27674 22545
rect 27618 22471 27674 22480
rect 27632 21457 27660 22471
rect 27618 21448 27674 21457
rect 27618 21383 27674 21392
rect 25134 18864 25190 18873
rect 25134 18799 25190 18808
rect 25148 18426 25176 18799
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25148 18222 25176 18362
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27632 16289 27660 16390
rect 27618 16280 27674 16289
rect 27618 16215 27674 16224
rect 25134 14240 25190 14249
rect 25134 14175 25190 14184
rect 25148 14074 25176 14175
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25148 13870 25176 14010
rect 24780 13786 24900 13814
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 22282 10160 22338 10169
rect 21364 10124 21416 10130
rect 21192 10084 21364 10112
rect 20904 10066 20956 10072
rect 22282 10095 22338 10104
rect 23572 10124 23624 10130
rect 21364 10066 21416 10072
rect 23572 10066 23624 10072
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20548 8294 20576 8978
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 20180 7206 20208 7890
rect 20548 7857 20576 8230
rect 20534 7848 20590 7857
rect 20534 7783 20590 7792
rect 20548 7342 20576 7783
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19628 6322 19656 6802
rect 20180 6458 20208 7142
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19628 6225 19656 6258
rect 20180 6254 20208 6394
rect 20168 6248 20220 6254
rect 19614 6216 19670 6225
rect 20168 6190 20220 6196
rect 19614 6151 19670 6160
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 5370 19840 5646
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20640 2650 20668 9862
rect 20916 9450 20944 10066
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 21376 9178 21404 10066
rect 23584 9654 23612 10066
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20916 7546 20944 7890
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20916 7449 20944 7482
rect 20902 7440 20958 7449
rect 20902 7375 20958 7384
rect 21652 5302 21680 9318
rect 24228 8430 24256 13126
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 13786
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24766 11384 24822 11393
rect 24766 11319 24822 11328
rect 24780 11082 24808 11319
rect 24872 11218 24900 12038
rect 24964 11558 24992 12242
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24768 11076 24820 11082
rect 24768 11018 24820 11024
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24872 10810 24900 11154
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24596 10130 24624 10406
rect 24584 10124 24636 10130
rect 24636 10084 24716 10112
rect 24584 10066 24636 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 10084
rect 24964 10033 24992 11494
rect 24950 10024 25006 10033
rect 24950 9959 25006 9968
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9761 24808 9862
rect 24766 9752 24822 9761
rect 24676 9716 24728 9722
rect 24766 9687 24822 9696
rect 24676 9658 24728 9664
rect 24766 8800 24822 8809
rect 24289 8732 24585 8752
rect 24766 8735 24822 8744
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24780 8634 24808 8735
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 27618 6896 27674 6905
rect 24676 6860 24728 6866
rect 27618 6831 27674 6840
rect 24676 6802 24728 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6118 24716 6802
rect 27632 6458 27660 6831
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 26884 6112 26936 6118
rect 26884 6054 26936 6060
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24044 4049 24072 4082
rect 24030 4040 24086 4049
rect 24030 3975 24086 3984
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 2310 23244 2382
rect 24676 2372 24728 2378
rect 24676 2314 24728 2320
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 20260 2100 20312 2106
rect 20260 2042 20312 2048
rect 19246 82 19302 480
rect 18984 54 19302 82
rect 20272 82 20300 2042
rect 22006 1864 22062 1873
rect 22006 1799 22062 1808
rect 20626 82 20682 480
rect 20272 54 20682 82
rect 15290 0 15346 54
rect 16578 0 16634 54
rect 17958 0 18014 54
rect 19246 0 19302 54
rect 20626 0 20682 54
rect 21914 82 21970 480
rect 22020 82 22048 1799
rect 21914 54 22048 82
rect 23294 128 23350 480
rect 23294 76 23296 128
rect 23348 76 23350 128
rect 21914 0 21970 54
rect 23294 0 23350 76
rect 24582 82 24638 480
rect 24688 82 24716 2314
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 24582 54 24716 82
rect 25962 82 26018 480
rect 26068 82 26096 2246
rect 25962 54 26096 82
rect 26896 82 26924 6054
rect 27618 5400 27674 5409
rect 27618 5335 27674 5344
rect 27632 5302 27660 5335
rect 27620 5296 27672 5302
rect 27620 5238 27672 5244
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3777 27660 3878
rect 27618 3768 27674 3777
rect 27618 3703 27674 3712
rect 27618 1728 27674 1737
rect 27618 1663 27674 1672
rect 27632 785 27660 1663
rect 27618 776 27674 785
rect 27618 711 27674 720
rect 27250 82 27306 480
rect 26896 54 27306 82
rect 24582 0 24638 54
rect 25962 0 26018 54
rect 27250 0 27306 54
<< via2 >>
rect 1858 26696 1914 26752
rect 1306 25472 1362 25528
rect 1582 24112 1638 24168
rect 1398 23568 1454 23624
rect 1398 22888 1454 22944
rect 110 17040 166 17096
rect 110 10648 166 10704
rect 110 3032 166 3088
rect 1582 21664 1638 21720
rect 1582 20304 1638 20360
rect 1490 19080 1546 19136
rect 1582 17992 1638 18048
rect 1950 17176 2006 17232
rect 1582 17040 1638 17096
rect 1398 14456 1454 14512
rect 1582 12280 1638 12336
rect 2042 16360 2098 16416
rect 1950 15136 2006 15192
rect 2686 18672 2742 18728
rect 1858 13504 1914 13560
rect 1766 3984 1822 4040
rect 1950 3984 2006 4040
rect 2962 14456 3018 14512
rect 3790 18808 3846 18864
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 4802 18264 4858 18320
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5722 18264 5778 18320
rect 5630 17584 5686 17640
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 3606 12688 3662 12744
rect 2686 9560 2742 9616
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5998 13096 6054 13152
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5906 11600 5962 11656
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4986 9968 5042 10024
rect 4618 6568 4674 6624
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 4526 5072 4582 5128
rect 5354 5208 5410 5264
rect 3422 2080 3478 2136
rect 4434 1808 4490 1864
rect 3514 1264 3570 1320
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5446 1128 5502 1184
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5630 2488 5686 2544
rect 7378 7384 7434 7440
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 8298 15000 8354 15056
rect 8758 21392 8814 21448
rect 8666 13776 8722 13832
rect 7746 6840 7802 6896
rect 7562 2896 7618 2952
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 13266 24112 13322 24168
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 8850 6160 8906 6216
rect 8114 1672 8170 1728
rect 8758 3984 8814 4040
rect 8942 3168 8998 3224
rect 9494 12960 9550 13016
rect 10782 20440 10838 20496
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10322 12144 10378 12200
rect 9678 10648 9734 10704
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 13358 18808 13414 18864
rect 13450 18708 13452 18728
rect 13452 18708 13504 18728
rect 13504 18708 13506 18728
rect 13450 18672 13506 18708
rect 11794 18264 11850 18320
rect 12622 17176 12678 17232
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9862 9424 9918 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10690 8472 10746 8528
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 12162 12724 12164 12744
rect 12164 12724 12216 12744
rect 12216 12724 12218 12744
rect 12162 12688 12218 12724
rect 12346 12688 12402 12744
rect 12070 10512 12126 10568
rect 11978 9560 12034 9616
rect 12438 9968 12494 10024
rect 12530 8472 12586 8528
rect 11610 7248 11666 7304
rect 10782 3984 10838 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12530 3576 12586 3632
rect 11702 2896 11758 2952
rect 11794 2488 11850 2544
rect 11334 1264 11390 1320
rect 13082 9424 13138 9480
rect 13358 9968 13414 10024
rect 13266 9560 13322 9616
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15290 20984 15346 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 13542 10104 13598 10160
rect 13450 9424 13506 9480
rect 13450 8472 13506 8528
rect 12806 3984 12862 4040
rect 13910 9968 13966 10024
rect 13818 5208 13874 5264
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14186 12688 14242 12744
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15106 15544 15162 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14462 10648 14518 10704
rect 14278 9968 14334 10024
rect 14094 9560 14150 9616
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15934 17720 15990 17776
rect 17406 23604 17408 23624
rect 17408 23604 17460 23624
rect 17460 23604 17462 23624
rect 17406 23568 17462 23604
rect 17314 18264 17370 18320
rect 18326 20440 18382 20496
rect 17958 17720 18014 17776
rect 18602 17584 18658 17640
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19430 24112 19486 24168
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19338 17040 19394 17096
rect 15934 15020 15990 15056
rect 15934 15000 15936 15020
rect 15936 15000 15988 15020
rect 15988 15000 15990 15020
rect 15566 13776 15622 13832
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15474 8200 15530 8256
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 16394 8200 16450 8256
rect 15290 7248 15346 7304
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 17130 8472 17186 8528
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14554 3576 14610 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14002 3168 14058 3224
rect 15566 5072 15622 5128
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17590 7112 17646 7168
rect 18510 7112 18566 7168
rect 18326 6840 18382 6896
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 23754 26560 23810 26616
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19982 14456 20038 14512
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18878 11600 18934 11656
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19522 12144 19578 12200
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 8200 19486 8256
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 18970 6160 19026 6216
rect 18510 3984 18566 4040
rect 18878 2488 18934 2544
rect 20902 13368 20958 13424
rect 22374 13232 22430 13288
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 23432 24822 23488
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 18264 24178 18320
rect 24214 17720 24270 17776
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17312 24822 17368
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25134 25064 25190 25120
rect 27250 23568 27306 23624
rect 27618 22480 27674 22536
rect 27618 21392 27674 21448
rect 25134 18808 25190 18864
rect 27618 16224 27674 16280
rect 25134 14184 25190 14240
rect 22282 10104 22338 10160
rect 20534 7792 20590 7848
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19614 6160 19670 6216
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20902 7384 20958 7440
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11328 24822 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24950 9968 25006 10024
rect 24766 9696 24822 9752
rect 24766 8744 24822 8800
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 27618 6840 27674 6896
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24030 3984 24086 4040
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 22006 1808 22062 1864
rect 27618 5344 27674 5400
rect 27618 3712 27674 3768
rect 27618 1672 27674 1728
rect 27618 720 27674 776
<< metal3 >>
rect 0 27208 480 27328
rect 62 26754 122 27208
rect 27520 27072 28000 27192
rect 1853 26754 1919 26757
rect 62 26752 1919 26754
rect 62 26696 1858 26752
rect 1914 26696 1919 26752
rect 62 26694 1919 26696
rect 1853 26691 1919 26694
rect 23749 26618 23815 26621
rect 27662 26618 27722 27072
rect 23749 26616 27722 26618
rect 23749 26560 23754 26616
rect 23810 26560 27722 26616
rect 23749 26558 27722 26560
rect 23749 26555 23815 26558
rect 0 25984 480 26104
rect 62 25530 122 25984
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 27520 25576 28000 25696
rect 19610 25535 19930 25536
rect 1301 25530 1367 25533
rect 62 25528 1367 25530
rect 62 25472 1306 25528
rect 1362 25472 1367 25528
rect 62 25470 1367 25472
rect 1301 25467 1367 25470
rect 25129 25122 25195 25125
rect 27662 25122 27722 25576
rect 25129 25120 27722 25122
rect 25129 25064 25134 25120
rect 25190 25064 27722 25120
rect 25129 25062 27722 25064
rect 25129 25059 25195 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24624 480 24744
rect 62 24170 122 24624
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 1577 24170 1643 24173
rect 62 24168 1643 24170
rect 62 24112 1582 24168
rect 1638 24112 1643 24168
rect 62 24110 1643 24112
rect 1577 24107 1643 24110
rect 13261 24170 13327 24173
rect 19425 24170 19491 24173
rect 13261 24168 19491 24170
rect 13261 24112 13266 24168
rect 13322 24112 19430 24168
rect 19486 24112 19491 24168
rect 13261 24110 19491 24112
rect 13261 24107 13327 24110
rect 19425 24107 19491 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 27520 23944 28000 24064
rect 24277 23903 24597 23904
rect 1393 23626 1459 23629
rect 1526 23626 1532 23628
rect 1393 23624 1532 23626
rect 1393 23568 1398 23624
rect 1454 23568 1532 23624
rect 1393 23566 1532 23568
rect 1393 23563 1459 23566
rect 1526 23564 1532 23566
rect 1596 23564 1602 23628
rect 17401 23626 17467 23629
rect 27245 23626 27311 23629
rect 17401 23624 27311 23626
rect 17401 23568 17406 23624
rect 17462 23568 27250 23624
rect 27306 23568 27311 23624
rect 17401 23566 27311 23568
rect 17401 23563 17467 23566
rect 27245 23563 27311 23566
rect 0 23400 480 23520
rect 24761 23490 24827 23493
rect 27662 23490 27722 23944
rect 24761 23488 27722 23490
rect 24761 23432 24766 23488
rect 24822 23432 27722 23488
rect 24761 23430 27722 23432
rect 24761 23427 24827 23430
rect 10277 23424 10597 23425
rect 62 22946 122 23400
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 1393 22946 1459 22949
rect 62 22944 1459 22946
rect 62 22888 1398 22944
rect 1454 22888 1459 22944
rect 62 22886 1459 22888
rect 1393 22883 1459 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 27520 22536 28000 22568
rect 27520 22480 27618 22536
rect 27674 22480 28000 22536
rect 27520 22448 28000 22480
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1577 21722 1643 21725
rect 62 21720 1643 21722
rect 62 21664 1582 21720
rect 1638 21664 1643 21720
rect 62 21662 1643 21664
rect 1577 21659 1643 21662
rect 8753 21450 8819 21453
rect 27613 21450 27679 21453
rect 8753 21448 27679 21450
rect 8753 21392 8758 21448
rect 8814 21392 27618 21448
rect 27674 21392 27679 21448
rect 8753 21390 27679 21392
rect 8753 21387 8819 21390
rect 27613 21387 27679 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27654 21178 27660 21180
rect 27248 21118 27660 21178
rect 15285 21042 15351 21045
rect 27248 21042 27308 21118
rect 27654 21116 27660 21118
rect 27724 21116 27730 21180
rect 15285 21040 27308 21042
rect 15285 20984 15290 21040
rect 15346 20984 27308 21040
rect 15285 20982 27308 20984
rect 15285 20979 15351 20982
rect 0 20816 480 20936
rect 27520 20908 28000 20936
rect 27520 20844 27660 20908
rect 27724 20844 28000 20908
rect 27520 20816 28000 20844
rect 62 20362 122 20816
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10777 20498 10843 20501
rect 18321 20498 18387 20501
rect 10777 20496 18387 20498
rect 10777 20440 10782 20496
rect 10838 20440 18326 20496
rect 18382 20440 18387 20496
rect 10777 20438 18387 20440
rect 10777 20435 10843 20438
rect 18321 20435 18387 20438
rect 1577 20362 1643 20365
rect 62 20360 1643 20362
rect 62 20304 1582 20360
rect 1638 20304 1643 20360
rect 62 20302 1643 20304
rect 1577 20299 1643 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19592 480 19712
rect 5610 19616 5930 19617
rect 62 19138 122 19592
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19320 28000 19440
rect 1485 19138 1551 19141
rect 62 19136 1551 19138
rect 62 19080 1490 19136
rect 1546 19080 1551 19136
rect 62 19078 1551 19080
rect 1485 19075 1551 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 3785 18866 3851 18869
rect 13353 18866 13419 18869
rect 3785 18864 13419 18866
rect 3785 18808 3790 18864
rect 3846 18808 13358 18864
rect 13414 18808 13419 18864
rect 3785 18806 13419 18808
rect 3785 18803 3851 18806
rect 13353 18803 13419 18806
rect 25129 18866 25195 18869
rect 27662 18866 27722 19320
rect 25129 18864 27722 18866
rect 25129 18808 25134 18864
rect 25190 18808 27722 18864
rect 25129 18806 27722 18808
rect 25129 18803 25195 18806
rect 2681 18730 2747 18733
rect 13445 18730 13511 18733
rect 2681 18728 13511 18730
rect 2681 18672 2686 18728
rect 2742 18672 13450 18728
rect 13506 18672 13511 18728
rect 2681 18670 13511 18672
rect 2681 18667 2747 18670
rect 13445 18667 13511 18670
rect 5610 18528 5930 18529
rect 0 18368 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 62 18050 122 18368
rect 4797 18322 4863 18325
rect 5717 18322 5783 18325
rect 4797 18320 5783 18322
rect 4797 18264 4802 18320
rect 4858 18264 5722 18320
rect 5778 18264 5783 18320
rect 4797 18262 5783 18264
rect 4797 18259 4863 18262
rect 5717 18259 5783 18262
rect 11789 18322 11855 18325
rect 17309 18322 17375 18325
rect 24117 18322 24183 18325
rect 11789 18320 24183 18322
rect 11789 18264 11794 18320
rect 11850 18264 17314 18320
rect 17370 18264 24122 18320
rect 24178 18264 24183 18320
rect 11789 18262 24183 18264
rect 11789 18259 11855 18262
rect 17309 18259 17375 18262
rect 24117 18259 24183 18262
rect 1577 18050 1643 18053
rect 62 18048 1643 18050
rect 62 17992 1582 18048
rect 1638 17992 1643 18048
rect 62 17990 1643 17992
rect 1577 17987 1643 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 15929 17778 15995 17781
rect 17953 17778 18019 17781
rect 24209 17778 24275 17781
rect 15929 17776 24275 17778
rect 15929 17720 15934 17776
rect 15990 17720 17958 17776
rect 18014 17720 24214 17776
rect 24270 17720 24275 17776
rect 15929 17718 24275 17720
rect 15929 17715 15995 17718
rect 17953 17715 18019 17718
rect 24209 17715 24275 17718
rect 27520 17688 28000 17808
rect 5625 17642 5691 17645
rect 18597 17642 18663 17645
rect 5625 17640 18663 17642
rect 5625 17584 5630 17640
rect 5686 17584 18602 17640
rect 18658 17584 18663 17640
rect 5625 17582 18663 17584
rect 5625 17579 5691 17582
rect 18597 17579 18663 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 24761 17370 24827 17373
rect 27662 17370 27722 17688
rect 24761 17368 27722 17370
rect 24761 17312 24766 17368
rect 24822 17312 27722 17368
rect 24761 17310 27722 17312
rect 24761 17307 24827 17310
rect 1945 17234 2011 17237
rect 12617 17234 12683 17237
rect 1945 17232 12683 17234
rect 1945 17176 1950 17232
rect 2006 17176 12622 17232
rect 12678 17176 12683 17232
rect 1945 17174 12683 17176
rect 1945 17171 2011 17174
rect 12617 17171 12683 17174
rect 0 17096 480 17128
rect 0 17040 110 17096
rect 166 17040 480 17096
rect 0 17008 480 17040
rect 1577 17098 1643 17101
rect 19333 17098 19399 17101
rect 1577 17096 19399 17098
rect 1577 17040 1582 17096
rect 1638 17040 19338 17096
rect 19394 17040 19399 17096
rect 1577 17038 19399 17040
rect 1577 17035 1643 17038
rect 19333 17035 19399 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 2037 16418 2103 16421
rect 62 16416 2103 16418
rect 62 16360 2042 16416
rect 2098 16360 2103 16416
rect 62 16358 2103 16360
rect 62 15904 122 16358
rect 2037 16355 2103 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 16280 28000 16312
rect 27520 16224 27618 16280
rect 27674 16224 28000 16280
rect 27520 16192 28000 16224
rect 0 15784 480 15904
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 9622 15540 9628 15604
rect 9692 15602 9698 15604
rect 15101 15602 15167 15605
rect 9692 15600 15167 15602
rect 9692 15544 15106 15600
rect 15162 15544 15167 15600
rect 9692 15542 15167 15544
rect 9692 15540 9698 15542
rect 15101 15539 15167 15542
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 1945 15194 2011 15197
rect 62 15192 2011 15194
rect 62 15136 1950 15192
rect 2006 15136 2011 15192
rect 62 15134 2011 15136
rect 62 14680 122 15134
rect 1945 15131 2011 15134
rect 8293 15058 8359 15061
rect 15929 15058 15995 15061
rect 8293 15056 15995 15058
rect 8293 15000 8298 15056
rect 8354 15000 15934 15056
rect 15990 15000 15995 15056
rect 8293 14998 15995 15000
rect 8293 14995 8359 14998
rect 15929 14995 15995 14998
rect 10277 14720 10597 14721
rect 0 14560 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 27520 14696 28000 14816
rect 19610 14655 19930 14656
rect 1393 14514 1459 14517
rect 2957 14514 3023 14517
rect 19977 14514 20043 14517
rect 1393 14512 20043 14514
rect 1393 14456 1398 14512
rect 1454 14456 2962 14512
rect 3018 14456 19982 14512
rect 20038 14456 20043 14512
rect 1393 14454 20043 14456
rect 1393 14451 1459 14454
rect 2957 14451 3023 14454
rect 19977 14451 20043 14454
rect 25129 14242 25195 14245
rect 27662 14242 27722 14696
rect 25129 14240 27722 14242
rect 25129 14184 25134 14240
rect 25190 14184 27722 14240
rect 25129 14182 27722 14184
rect 25129 14179 25195 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 8661 13834 8727 13837
rect 15561 13834 15627 13837
rect 8661 13832 15627 13834
rect 8661 13776 8666 13832
rect 8722 13776 15566 13832
rect 15622 13776 15627 13832
rect 8661 13774 15627 13776
rect 8661 13771 8727 13774
rect 15561 13771 15627 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 1853 13562 1919 13565
rect 62 13560 4170 13562
rect 62 13504 1858 13560
rect 1914 13504 4170 13560
rect 62 13502 4170 13504
rect 62 13320 122 13502
rect 1853 13499 1919 13502
rect 4110 13426 4170 13502
rect 20897 13426 20963 13429
rect 4110 13424 20963 13426
rect 4110 13368 20902 13424
rect 20958 13368 20963 13424
rect 4110 13366 20963 13368
rect 20897 13363 20963 13366
rect 0 13200 480 13320
rect 22369 13290 22435 13293
rect 13770 13288 22435 13290
rect 13770 13232 22374 13288
rect 22430 13232 22435 13288
rect 13770 13230 22435 13232
rect 5993 13154 6059 13157
rect 13770 13154 13830 13230
rect 22369 13227 22435 13230
rect 5993 13152 13830 13154
rect 5993 13096 5998 13152
rect 6054 13096 13830 13152
rect 5993 13094 13830 13096
rect 5993 13091 6059 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13184
rect 24277 13023 24597 13024
rect 9489 13018 9555 13021
rect 9622 13018 9628 13020
rect 9489 13016 9628 13018
rect 9489 12960 9494 13016
rect 9550 12960 9628 13016
rect 9489 12958 9628 12960
rect 9489 12955 9555 12958
rect 9622 12956 9628 12958
rect 9692 12956 9698 13020
rect 3601 12746 3667 12749
rect 12157 12746 12223 12749
rect 3601 12744 12223 12746
rect 3601 12688 3606 12744
rect 3662 12688 12162 12744
rect 12218 12688 12223 12744
rect 3601 12686 12223 12688
rect 3601 12683 3667 12686
rect 12157 12683 12223 12686
rect 12341 12746 12407 12749
rect 14181 12746 14247 12749
rect 27662 12746 27722 13064
rect 12341 12744 27722 12746
rect 12341 12688 12346 12744
rect 12402 12688 14186 12744
rect 14242 12688 27722 12744
rect 12341 12686 27722 12688
rect 12341 12683 12407 12686
rect 14181 12683 14247 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 54 12276 60 12340
rect 124 12338 130 12340
rect 1577 12338 1643 12341
rect 124 12336 1643 12338
rect 124 12280 1582 12336
rect 1638 12280 1643 12336
rect 124 12278 1643 12280
rect 124 12276 130 12278
rect 1577 12275 1643 12278
rect 10317 12202 10383 12205
rect 19517 12202 19583 12205
rect 10317 12200 19583 12202
rect 10317 12144 10322 12200
rect 10378 12144 19522 12200
rect 19578 12144 19583 12200
rect 10317 12142 19583 12144
rect 10317 12139 10383 12142
rect 19517 12139 19583 12142
rect 0 12068 480 12096
rect 0 12004 60 12068
rect 124 12004 480 12068
rect 0 11976 480 12004
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 5901 11658 5967 11661
rect 18873 11658 18939 11661
rect 5901 11656 18939 11658
rect 5901 11600 5906 11656
rect 5962 11600 18878 11656
rect 18934 11600 18939 11656
rect 5901 11598 18939 11600
rect 5901 11595 5967 11598
rect 18873 11595 18939 11598
rect 27520 11568 28000 11688
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 24761 11386 24827 11389
rect 27662 11386 27722 11568
rect 24761 11384 27722 11386
rect 24761 11328 24766 11384
rect 24822 11328 27722 11384
rect 24761 11326 27722 11328
rect 24761 11323 24827 11326
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10704 480 10736
rect 0 10648 110 10704
rect 166 10648 480 10704
rect 0 10616 480 10648
rect 9673 10706 9739 10709
rect 14457 10706 14523 10709
rect 9673 10704 14523 10706
rect 9673 10648 9678 10704
rect 9734 10648 14462 10704
rect 14518 10648 14523 10704
rect 9673 10646 14523 10648
rect 9673 10643 9739 10646
rect 14457 10643 14523 10646
rect 4102 10508 4108 10572
rect 4172 10570 4178 10572
rect 12065 10570 12131 10573
rect 4172 10568 12131 10570
rect 4172 10512 12070 10568
rect 12126 10512 12131 10568
rect 4172 10510 12131 10512
rect 4172 10508 4178 10510
rect 12065 10507 12131 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 13537 10162 13603 10165
rect 22277 10162 22343 10165
rect 13537 10160 22343 10162
rect 13537 10104 13542 10160
rect 13598 10104 22282 10160
rect 22338 10104 22343 10160
rect 13537 10102 22343 10104
rect 13537 10099 13603 10102
rect 22277 10099 22343 10102
rect 4981 10026 5047 10029
rect 12433 10026 12499 10029
rect 4981 10024 12499 10026
rect 4981 9968 4986 10024
rect 5042 9968 12438 10024
rect 12494 9968 12499 10024
rect 4981 9966 12499 9968
rect 4981 9963 5047 9966
rect 12433 9963 12499 9966
rect 13353 10026 13419 10029
rect 13905 10026 13971 10029
rect 13353 10024 13971 10026
rect 13353 9968 13358 10024
rect 13414 9968 13910 10024
rect 13966 9968 13971 10024
rect 13353 9966 13971 9968
rect 13353 9963 13419 9966
rect 13905 9963 13971 9966
rect 14273 10026 14339 10029
rect 24945 10026 25011 10029
rect 14273 10024 25011 10026
rect 14273 9968 14278 10024
rect 14334 9968 24950 10024
rect 25006 9968 25011 10024
rect 14273 9966 25011 9968
rect 14273 9963 14339 9966
rect 24945 9963 25011 9966
rect 27520 10028 28000 10056
rect 27520 9964 27660 10028
rect 27724 9964 28000 10028
rect 27520 9936 28000 9964
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 24761 9754 24827 9757
rect 27654 9754 27660 9756
rect 24761 9752 27660 9754
rect 24761 9696 24766 9752
rect 24822 9696 27660 9752
rect 24761 9694 27660 9696
rect 24761 9691 24827 9694
rect 27654 9692 27660 9694
rect 27724 9692 27730 9756
rect 54 9590 60 9654
rect 124 9652 130 9654
rect 124 9618 674 9652
rect 2681 9618 2747 9621
rect 11973 9618 12039 9621
rect 124 9616 12039 9618
rect 124 9592 2686 9616
rect 124 9590 130 9592
rect 614 9560 2686 9592
rect 2742 9560 11978 9616
rect 12034 9560 12039 9616
rect 614 9558 12039 9560
rect 2681 9555 2747 9558
rect 11973 9555 12039 9558
rect 13261 9618 13327 9621
rect 14089 9618 14155 9621
rect 13261 9616 14155 9618
rect 13261 9560 13266 9616
rect 13322 9560 14094 9616
rect 14150 9560 14155 9616
rect 13261 9558 14155 9560
rect 13261 9555 13327 9558
rect 14089 9555 14155 9558
rect 0 9484 480 9512
rect 0 9420 60 9484
rect 124 9420 480 9484
rect 0 9392 480 9420
rect 9857 9482 9923 9485
rect 13077 9482 13143 9485
rect 13445 9482 13511 9485
rect 9857 9480 13511 9482
rect 9857 9424 9862 9480
rect 9918 9424 13082 9480
rect 13138 9424 13450 9480
rect 13506 9424 13511 9480
rect 9857 9422 13511 9424
rect 9857 9419 9923 9422
rect 13077 9419 13143 9422
rect 13445 9419 13511 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 24761 8802 24827 8805
rect 27654 8802 27660 8804
rect 24761 8800 27660 8802
rect 24761 8744 24766 8800
rect 24822 8744 27660 8800
rect 24761 8742 27660 8744
rect 24761 8739 24827 8742
rect 27654 8740 27660 8742
rect 27724 8740 27730 8804
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 10685 8530 10751 8533
rect 12525 8530 12591 8533
rect 13445 8530 13511 8533
rect 17125 8530 17191 8533
rect 10685 8528 17191 8530
rect 10685 8472 10690 8528
rect 10746 8472 12530 8528
rect 12586 8472 13450 8528
rect 13506 8472 17130 8528
rect 17186 8472 17191 8528
rect 10685 8470 17191 8472
rect 10685 8467 10751 8470
rect 12525 8467 12591 8470
rect 13445 8467 13511 8470
rect 17125 8467 17191 8470
rect 27520 8532 28000 8560
rect 27520 8468 27660 8532
rect 27724 8468 28000 8532
rect 27520 8440 28000 8468
rect 0 8168 480 8288
rect 15469 8258 15535 8261
rect 16389 8258 16455 8261
rect 19425 8258 19491 8261
rect 15469 8256 19491 8258
rect 15469 8200 15474 8256
rect 15530 8200 16394 8256
rect 16450 8200 19430 8256
rect 19486 8200 19491 8256
rect 15469 8198 19491 8200
rect 15469 8195 15535 8198
rect 16389 8195 16455 8198
rect 19425 8195 19491 8198
rect 10277 8192 10597 8193
rect 62 7850 122 8168
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 20529 7850 20595 7853
rect 62 7848 20595 7850
rect 62 7792 20534 7848
rect 20590 7792 20595 7848
rect 62 7790 20595 7792
rect 20529 7787 20595 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 7373 7442 7439 7445
rect 20897 7442 20963 7445
rect 7373 7440 20963 7442
rect 7373 7384 7378 7440
rect 7434 7384 20902 7440
rect 20958 7384 20963 7440
rect 7373 7382 20963 7384
rect 7373 7379 7439 7382
rect 20897 7379 20963 7382
rect 11605 7306 11671 7309
rect 15285 7306 15351 7309
rect 11605 7304 15351 7306
rect 11605 7248 11610 7304
rect 11666 7248 15290 7304
rect 15346 7248 15351 7304
rect 11605 7246 15351 7248
rect 11605 7243 11671 7246
rect 15285 7243 15351 7246
rect 17585 7170 17651 7173
rect 18505 7170 18571 7173
rect 17585 7168 18571 7170
rect 17585 7112 17590 7168
rect 17646 7112 18510 7168
rect 18566 7112 18571 7168
rect 17585 7110 18571 7112
rect 17585 7107 17651 7110
rect 18505 7107 18571 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6900 480 6928
rect 0 6836 60 6900
rect 124 6836 480 6900
rect 0 6808 480 6836
rect 7741 6898 7807 6901
rect 18321 6898 18387 6901
rect 7741 6896 18387 6898
rect 7741 6840 7746 6896
rect 7802 6840 18326 6896
rect 18382 6840 18387 6896
rect 7741 6838 18387 6840
rect 7741 6835 7807 6838
rect 18321 6835 18387 6838
rect 27520 6896 28000 6928
rect 27520 6840 27618 6896
rect 27674 6840 28000 6896
rect 27520 6808 28000 6840
rect 54 6564 60 6628
rect 124 6626 130 6628
rect 4613 6626 4679 6629
rect 124 6624 4679 6626
rect 124 6568 4618 6624
rect 4674 6568 4679 6624
rect 124 6566 4679 6568
rect 124 6564 130 6566
rect 4613 6563 4679 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 8845 6218 8911 6221
rect 18965 6218 19031 6221
rect 19609 6218 19675 6221
rect 8845 6216 19675 6218
rect 8845 6160 8850 6216
rect 8906 6160 18970 6216
rect 19026 6160 19614 6216
rect 19670 6160 19675 6216
rect 8845 6158 19675 6160
rect 8845 6155 8911 6158
rect 18965 6155 19031 6158
rect 19609 6155 19675 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5584 480 5704
rect 62 5130 122 5584
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 27520 5400 28000 5432
rect 27520 5344 27618 5400
rect 27674 5344 28000 5400
rect 27520 5312 28000 5344
rect 5349 5266 5415 5269
rect 13813 5266 13879 5269
rect 4110 5264 13879 5266
rect 4110 5208 5354 5264
rect 5410 5208 13818 5264
rect 13874 5208 13879 5264
rect 4110 5206 13879 5208
rect 4110 5130 4170 5206
rect 5349 5203 5415 5206
rect 13813 5203 13879 5206
rect 62 5070 4170 5130
rect 4521 5130 4587 5133
rect 15561 5130 15627 5133
rect 4521 5128 15627 5130
rect 4521 5072 4526 5128
rect 4582 5072 15566 5128
rect 15622 5072 15627 5128
rect 4521 5070 15627 5072
rect 4521 5067 4587 5070
rect 15561 5067 15627 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4360 480 4480
rect 5610 4384 5930 4385
rect 62 4042 122 4360
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 1761 4042 1827 4045
rect 62 4040 1827 4042
rect 62 3984 1766 4040
rect 1822 3984 1827 4040
rect 62 3982 1827 3984
rect 1761 3979 1827 3982
rect 1945 4042 2011 4045
rect 8753 4042 8819 4045
rect 10777 4042 10843 4045
rect 12801 4042 12867 4045
rect 1945 4040 4170 4042
rect 1945 3984 1950 4040
rect 2006 3984 4170 4040
rect 1945 3982 4170 3984
rect 1945 3979 2011 3982
rect 4110 3634 4170 3982
rect 8753 4040 12867 4042
rect 8753 3984 8758 4040
rect 8814 3984 10782 4040
rect 10838 3984 12806 4040
rect 12862 3984 12867 4040
rect 8753 3982 12867 3984
rect 8753 3979 8819 3982
rect 10777 3979 10843 3982
rect 12801 3979 12867 3982
rect 18505 4042 18571 4045
rect 24025 4042 24091 4045
rect 18505 4040 24091 4042
rect 18505 3984 18510 4040
rect 18566 3984 24030 4040
rect 24086 3984 24091 4040
rect 18505 3982 24091 3984
rect 18505 3979 18571 3982
rect 24025 3979 24091 3982
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27520 3768 28000 3800
rect 27520 3712 27618 3768
rect 27674 3712 28000 3768
rect 27520 3680 28000 3712
rect 12525 3634 12591 3637
rect 14549 3634 14615 3637
rect 4110 3632 14615 3634
rect 4110 3576 12530 3632
rect 12586 3576 14554 3632
rect 14610 3576 14615 3632
rect 4110 3574 14615 3576
rect 12525 3571 12591 3574
rect 14549 3571 14615 3574
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 8937 3226 9003 3229
rect 13997 3226 14063 3229
rect 8937 3224 14063 3226
rect 8937 3168 8942 3224
rect 8998 3168 14002 3224
rect 14058 3168 14063 3224
rect 8937 3166 14063 3168
rect 8937 3163 9003 3166
rect 13997 3163 14063 3166
rect 0 3088 480 3120
rect 0 3032 110 3088
rect 166 3032 480 3088
rect 0 3000 480 3032
rect 7557 2954 7623 2957
rect 11697 2954 11763 2957
rect 7557 2952 11763 2954
rect 7557 2896 7562 2952
rect 7618 2896 11702 2952
rect 11758 2896 11763 2952
rect 7557 2894 11763 2896
rect 7557 2891 7623 2894
rect 11697 2891 11763 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5625 2546 5691 2549
rect 11789 2546 11855 2549
rect 5625 2544 11855 2546
rect 5625 2488 5630 2544
rect 5686 2488 11794 2544
rect 11850 2488 11855 2544
rect 5625 2486 11855 2488
rect 5625 2483 5691 2486
rect 11789 2483 11855 2486
rect 18873 2546 18939 2549
rect 18873 2544 27722 2546
rect 18873 2488 18878 2544
rect 18934 2488 27722 2544
rect 18873 2486 27722 2488
rect 18873 2483 18939 2486
rect 27662 2304 27722 2486
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 27520 2184 28000 2304
rect 24277 2143 24597 2144
rect 3417 2138 3483 2141
rect 62 2136 3483 2138
rect 62 2080 3422 2136
rect 3478 2080 3483 2136
rect 62 2078 3483 2080
rect 62 1896 122 2078
rect 3417 2075 3483 2078
rect 0 1776 480 1896
rect 4429 1866 4495 1869
rect 22001 1866 22067 1869
rect 4429 1864 22067 1866
rect 4429 1808 4434 1864
rect 4490 1808 22006 1864
rect 22062 1808 22067 1864
rect 4429 1806 22067 1808
rect 4429 1803 4495 1806
rect 22001 1803 22067 1806
rect 8109 1730 8175 1733
rect 27613 1730 27679 1733
rect 8109 1728 27679 1730
rect 8109 1672 8114 1728
rect 8170 1672 27618 1728
rect 27674 1672 27679 1728
rect 8109 1670 27679 1672
rect 8109 1667 8175 1670
rect 27613 1667 27679 1670
rect 3509 1322 3575 1325
rect 11329 1322 11395 1325
rect 3509 1320 11395 1322
rect 3509 1264 3514 1320
rect 3570 1264 11334 1320
rect 11390 1264 11395 1320
rect 3509 1262 11395 1264
rect 3509 1259 3575 1262
rect 11329 1259 11395 1262
rect 5441 1186 5507 1189
rect 62 1184 5507 1186
rect 62 1128 5446 1184
rect 5502 1128 5507 1184
rect 62 1126 5507 1128
rect 62 672 122 1126
rect 5441 1123 5507 1126
rect 27520 776 28000 808
rect 27520 720 27618 776
rect 27674 720 28000 776
rect 27520 688 28000 720
rect 0 552 480 672
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 1532 23564 1596 23628
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 27660 21116 27724 21180
rect 27660 20844 27724 20908
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 9628 15540 9692 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 9628 12956 9692 13020
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 60 12276 124 12340
rect 60 12004 124 12068
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 4108 10508 4172 10572
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 27660 9964 27724 10028
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 27660 9692 27724 9756
rect 60 9590 124 9654
rect 60 9420 124 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 27660 8740 27724 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 27660 8468 27724 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 60 6836 124 6900
rect 60 6564 124 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 1531 23628 1597 23629
rect 1531 23564 1532 23628
rect 1596 23564 1597 23628
rect 1531 23563 1597 23564
rect 59 12340 125 12341
rect 59 12276 60 12340
rect 124 12276 125 12340
rect 59 12275 125 12276
rect 62 12069 122 12275
rect 59 12068 125 12069
rect 59 12004 60 12068
rect 124 12004 125 12068
rect 59 12003 125 12004
rect 1534 10658 1594 23563
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9627 15604 9693 15605
rect 9627 15540 9628 15604
rect 9692 15540 9693 15604
rect 9627 15539 9693 15540
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 9630 13021 9690 15539
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9627 13020 9693 13021
rect 9627 12956 9628 13020
rect 9692 12956 9693 13020
rect 9627 12955 9693 12956
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 59 9654 125 9655
rect 59 9590 60 9654
rect 124 9590 125 9654
rect 59 9589 125 9590
rect 62 9485 122 9589
rect 59 9484 125 9485
rect 59 9420 60 9484
rect 124 9420 125 9484
rect 59 9419 125 9420
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 59 6900 125 6901
rect 59 6836 60 6900
rect 124 6836 125 6900
rect 59 6835 125 6836
rect 62 6629 122 6835
rect 59 6628 125 6629
rect 59 6564 60 6628
rect 124 6564 125 6628
rect 59 6563 125 6564
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 27659 21180 27725 21181
rect 27659 21116 27660 21180
rect 27724 21116 27725 21180
rect 27659 21115 27725 21116
rect 27662 20909 27722 21115
rect 27659 20908 27725 20909
rect 27659 20844 27660 20908
rect 27724 20844 27725 20908
rect 27659 20843 27725 20844
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 27659 10028 27725 10029
rect 27659 9964 27660 10028
rect 27724 9964 27725 10028
rect 27659 9963 27725 9964
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 27662 9757 27722 9963
rect 27659 9756 27725 9757
rect 27659 9692 27660 9756
rect 27724 9692 27725 9756
rect 27659 9691 27725 9692
rect 27659 8804 27725 8805
rect 27659 8740 27660 8804
rect 27724 8740 27725 8804
rect 27659 8739 27725 8740
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 27662 8533 27722 8739
rect 27659 8532 27725 8533
rect 27659 8468 27660 8532
rect 27724 8468 27725 8532
rect 27659 8467 27725 8468
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 1446 10422 1682 10658
rect 4022 10572 4258 10658
rect 4022 10508 4108 10572
rect 4108 10508 4172 10572
rect 4172 10508 4258 10572
rect 4022 10422 4258 10508
<< metal5 >>
rect 1404 10658 4300 10700
rect 1404 10422 1446 10658
rect 1682 10422 4022 10658
rect 4258 10422 4300 10658
rect 1404 10380 4300 10422
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_14 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_0_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_42
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_43 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _226_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_69
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_81
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7820 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _208_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_109
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_inv_8  _204_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_134 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_171
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_190
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_190
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_194
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_226
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_238
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_38
timestamp 1586364061
transform 1 0 4600 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_2  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_66
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 590 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__C
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_161
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_274
timestamp 1586364061
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_49
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_53
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_66
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_70
timestamp 1586364061
transform 1 0 7544 0 -1 4896
box -38 -48 406 592
use scs8hd_or3_4  _101_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_74
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_97
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 590 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_23
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_104
timestamp 1586364061
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_172
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_9
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_14
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _173_
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_35
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _135_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_70
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_130
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_140
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_157
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_169
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_188
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_206
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_253
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_12
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_77
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_139
timestamp 1586364061
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_171
timestamp 1586364061
transform 1 0 16836 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_194
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_258
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_270
timestamp 1586364061
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_49
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_223
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_85
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_148
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_152
timestamp 1586364061
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_195
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_266
timestamp 1586364061
transform 1 0 25576 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _134_
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _107_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_221
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_275
timestamp 1586364061
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_14
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_or3_4  _155_
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_42
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_86
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 21344 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_222
timestamp 1586364061
transform 1 0 21528 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_246
timestamp 1586364061
transform 1 0 23736 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_nor4_4  _182_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__C
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_69
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_or3_4  _147_
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_or2_4  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_or2_4  _116_
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 682 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_225
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_237
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_249
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_8  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_259
timestamp 1586364061
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_271
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use scs8hd_or2_4  _089_
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _185_
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_120
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_161
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_190
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 22080 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_224
timestamp 1586364061
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_252
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_14
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _178_
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__178__D
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_90
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_158
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 22448 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_241
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 314 592
use scs8hd_or2_4  _126_
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 6900 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_87
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_261
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_273
timestamp 1586364061
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_18
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_38
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_115
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_187
timestamp 1586364061
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_191
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_204
timestamp 1586364061
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_222
timestamp 1586364061
transform 1 0 21528 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_225
timestamp 1586364061
transform 1 0 21804 0 -1 12512
box -38 -48 130 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_235
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_257
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__C
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__B
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__D
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _187_
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_95
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_99
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 1050 592
use scs8hd_buf_1  _127_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_116
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_155
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_170
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_185
timestamp 1586364061
transform 1 0 18124 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_194
timestamp 1586364061
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_198
timestamp 1586364061
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_228
timestamp 1586364061
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_264
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_276
timestamp 1586364061
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1472 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _175_
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_24
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__C
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _188_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__188__D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_or2_4  _136_
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_99
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_213
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 590 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_274
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _171_
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_1  _137_
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__B
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 20976 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_225
timestamp 1586364061
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_237
timestamp 1586364061
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_249
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_261
timestamp 1586364061
transform 1 0 25116 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_273
timestamp 1586364061
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_169
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_209
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_224
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_13
timestamp 1586364061
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_17
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_55
timestamp 1586364061
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_124
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_128
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_6  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_181
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_12
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _144_
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_94
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_126
timestamp 1586364061
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_130
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_181
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_227
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_17
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_49
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_116
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_131
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_127
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_149
timestamp 1586364061
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_171
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_200
timestamp 1586364061
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_259
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2300 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_74
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_133
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_174
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_198
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_182
timestamp 1586364061
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_50
timestamp 1586364061
transform 1 0 5704 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_30_58
timestamp 1586364061
transform 1 0 6440 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_96
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_100
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_113
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_132
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_187
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _180_
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_60
timestamp 1586364061
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_90
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_108
timestamp 1586364061
transform 1 0 11040 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_145
timestamp 1586364061
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_67
timestamp 1586364061
transform 1 0 7268 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_121
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_138
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_42
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_60
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_buf_1  _163_
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_67
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_88
timestamp 1586364061
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_84
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_107
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 866 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_109
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 590 592
use scs8hd_decap_4  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_124
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_137
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_148
timestamp 1586364061
transform 1 0 14720 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_165
timestamp 1586364061
transform 1 0 16284 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_177
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_243
timestamp 1586364061
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_238
timestamp 1586364061
transform 1 0 23000 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_250
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_262
timestamp 1586364061
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_68
timestamp 1586364061
transform 1 0 7360 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_80
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_84
timestamp 1586364061
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_91
timestamp 1586364061
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 774 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_76
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_102
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_106
timestamp 1586364061
transform 1 0 10856 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_113
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_137
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 8832 0 1 22304
box -38 -48 406 592
use scs8hd_decap_8  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_82
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_100
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_104
timestamp 1586364061
transform 1 0 10672 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _248_
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_259
timestamp 1586364061
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_263
timestamp 1586364061
transform 1 0 25300 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_275
timestamp 1586364061
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_18
timestamp 1586364061
transform 1 0 2760 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_30
timestamp 1586364061
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_99
timestamp 1586364061
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_111
timestamp 1586364061
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_135
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_147
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_50
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_65
timestamp 1586364061
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_69
timestamp 1586364061
transform 1 0 7452 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_76
timestamp 1586364061
transform 1 0 8096 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_77
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_89
timestamp 1586364061
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_81
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_85
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_81
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_93
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_109
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_150
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_154
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_178
timestamp 1586364061
transform 1 0 17480 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _247_
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_225
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 570 27520 626 28000 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 552 480 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 688 28000 808 6 address[2]
port 2 nsew default input
rlabel metal2 s 3238 0 3294 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 1766 27520 1822 28000 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[5]
port 5 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 address[6]
port 6 nsew default input
rlabel metal2 s 4618 0 4674 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal3 s 0 4360 480 4480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 bottom_right_grid_pin_13_
port 9 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 bottom_right_grid_pin_15_
port 10 nsew default input
rlabel metal3 s 27520 2184 28000 2304 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 bottom_right_grid_pin_3_
port 12 nsew default input
rlabel metal3 s 0 3000 480 3120 6 bottom_right_grid_pin_5_
port 13 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 bottom_right_grid_pin_7_
port 14 nsew default input
rlabel metal2 s 5906 0 5962 480 6 bottom_right_grid_pin_9_
port 15 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 27520 6808 28000 6928 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_out[0]
port 25 nsew default tristate
rlabel metal2 s 9402 27520 9458 28000 6 chanx_left_out[1]
port 26 nsew default tristate
rlabel metal3 s 27520 8440 28000 8560 6 chanx_left_out[2]
port 27 nsew default tristate
rlabel metal3 s 27520 9936 28000 10056 6 chanx_left_out[3]
port 28 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 chanx_left_out[4]
port 29 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[5]
port 30 nsew default tristate
rlabel metal3 s 27520 11568 28000 11688 6 chanx_left_out[6]
port 31 nsew default tristate
rlabel metal2 s 10690 27520 10746 28000 6 chanx_left_out[7]
port 32 nsew default tristate
rlabel metal2 s 11978 27520 12034 28000 6 chanx_left_out[8]
port 33 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 13266 27520 13322 28000 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal3 s 27520 14696 28000 14816 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal3 s 27520 16192 28000 16312 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 15750 27520 15806 28000 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 19246 0 19302 480 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 20626 0 20682 480 6 chany_top_in[2]
port 54 nsew default input
rlabel metal3 s 27520 19320 28000 19440 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal3 s 27520 20816 28000 20936 6 chany_top_in[6]
port 58 nsew default input
rlabel metal3 s 27520 22448 28000 22568 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 21914 0 21970 480 6 chany_top_in[8]
port 60 nsew default input
rlabel metal3 s 27520 23944 28000 24064 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 23386 27520 23442 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 23294 0 23350 480 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 1950 0 2006 480 6 data_in
port 70 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 71 nsew default input
rlabel metal2 s 24674 27520 24730 28000 6 left_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 0 23400 480 23520 6 left_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 25962 27520 26018 28000 6 top_left_grid_pin_13_
port 74 nsew default input
rlabel metal2 s 27250 0 27306 480 6 top_right_grid_pin_11_
port 75 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 top_right_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 0 27208 480 27328 6 top_right_grid_pin_15_
port 77 nsew default input
rlabel metal2 s 25962 0 26018 480 6 top_right_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 0 24624 480 24744 6 top_right_grid_pin_3_
port 79 nsew default input
rlabel metal3 s 0 25984 480 26104 6 top_right_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 27520 25576 28000 25696 6 top_right_grid_pin_7_
port 81 nsew default input
rlabel metal2 s 27250 27520 27306 28000 6 top_right_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
