magic
tech EFS8A
magscale 1 2
timestamp 1602873834
<< locali >>
rect 2547 20961 2582 20995
rect 4019 18785 4146 18819
rect 4019 16609 4146 16643
rect 4439 14569 4445 14603
rect 4439 14501 4473 14569
rect 13863 12257 13898 12291
rect 9229 12155 9263 12257
rect 9781 11543 9815 11713
rect 12081 11543 12115 11713
rect 13645 11543 13679 11849
rect 5175 11305 5181 11339
rect 5175 11237 5209 11305
rect 14139 11169 14174 11203
rect 9873 10489 9965 10523
rect 13277 9367 13311 9673
rect 8861 9027 8895 9129
rect 1443 7905 1478 7939
rect 7941 7905 8066 7939
rect 10793 7735 10827 7905
rect 9229 7191 9263 7429
rect 17411 6953 17417 6987
rect 17411 6885 17445 6953
rect 20855 6817 20982 6851
rect 2421 6171 2455 6409
rect 16859 5865 16865 5899
rect 16859 5797 16893 5865
rect 22511 5729 22546 5763
rect 12449 3451 12483 3689
rect 1547 3145 1685 3179
rect 19073 2975 19107 3145
<< viali >>
rect 1593 24361 1627 24395
rect 1409 24225 1443 24259
rect 1593 23817 1627 23851
rect 2697 23817 2731 23851
rect 2053 23681 2087 23715
rect 1409 23613 1443 23647
rect 2513 23613 2547 23647
rect 3157 23477 3191 23511
rect 1685 22933 1719 22967
rect 1593 21641 1627 21675
rect 1409 21437 1443 21471
rect 2053 21301 2087 21335
rect 1593 21097 1627 21131
rect 2651 21097 2685 21131
rect 1409 20961 1443 20995
rect 2513 20961 2547 20995
rect 2237 20553 2271 20587
rect 1476 20349 1510 20383
rect 1547 20213 1581 20247
rect 1869 20213 1903 20247
rect 2605 20213 2639 20247
rect 1593 20009 1627 20043
rect 2651 20009 2685 20043
rect 1409 19873 1443 19907
rect 2580 19873 2614 19907
rect 1593 19465 1627 19499
rect 2329 19465 2363 19499
rect 2651 19465 2685 19499
rect 3341 19465 3375 19499
rect 1409 19261 1443 19295
rect 2548 19261 2582 19295
rect 2973 19261 3007 19295
rect 2053 19125 2087 19159
rect 3525 19125 3559 19159
rect 1593 18921 1627 18955
rect 4215 18921 4249 18955
rect 1409 18785 1443 18819
rect 1961 18785 1995 18819
rect 2513 18785 2547 18819
rect 3985 18785 4019 18819
rect 2697 18649 2731 18683
rect 4859 18377 4893 18411
rect 2053 18173 2087 18207
rect 2881 18173 2915 18207
rect 3341 18173 3375 18207
rect 4788 18173 4822 18207
rect 5273 18173 5307 18207
rect 2973 18105 3007 18139
rect 1685 18037 1719 18071
rect 2513 18037 2547 18071
rect 4077 18037 4111 18071
rect 5733 18037 5767 18071
rect 3341 17833 3375 17867
rect 5779 17833 5813 17867
rect 2237 17697 2271 17731
rect 4721 17697 4755 17731
rect 5676 17697 5710 17731
rect 4077 17629 4111 17663
rect 6653 17629 6687 17663
rect 1961 17493 1995 17527
rect 2789 17493 2823 17527
rect 7435 17289 7469 17323
rect 2789 17221 2823 17255
rect 6193 17221 6227 17255
rect 3341 17153 3375 17187
rect 3617 17153 3651 17187
rect 5273 17153 5307 17187
rect 2329 17085 2363 17119
rect 7364 17085 7398 17119
rect 7757 17085 7791 17119
rect 3157 17017 3191 17051
rect 3433 17017 3467 17051
rect 5365 17017 5399 17051
rect 5917 17017 5951 17051
rect 1961 16949 1995 16983
rect 4353 16949 4387 16983
rect 5089 16949 5123 16983
rect 8309 16949 8343 16983
rect 2329 16745 2363 16779
rect 5273 16745 5307 16779
rect 2605 16677 2639 16711
rect 5365 16677 5399 16711
rect 8125 16677 8159 16711
rect 1476 16609 1510 16643
rect 3985 16609 4019 16643
rect 6009 16609 6043 16643
rect 6964 16609 6998 16643
rect 1961 16541 1995 16575
rect 2513 16541 2547 16575
rect 2789 16541 2823 16575
rect 8033 16541 8067 16575
rect 8309 16541 8343 16575
rect 3433 16473 3467 16507
rect 7067 16473 7101 16507
rect 1547 16405 1581 16439
rect 4215 16405 4249 16439
rect 7481 16405 7515 16439
rect 8953 16405 8987 16439
rect 1593 16201 1627 16235
rect 3065 16201 3099 16235
rect 6561 16201 6595 16235
rect 9597 16201 9631 16235
rect 4629 16133 4663 16167
rect 2789 16065 2823 16099
rect 3709 16065 3743 16099
rect 5917 16065 5951 16099
rect 7573 16065 7607 16099
rect 8401 15997 8435 16031
rect 2145 15929 2179 15963
rect 2237 15929 2271 15963
rect 3525 15929 3559 15963
rect 3778 15929 3812 15963
rect 4353 15929 4387 15963
rect 5273 15929 5307 15963
rect 5365 15929 5399 15963
rect 6929 15929 6963 15963
rect 7021 15929 7055 15963
rect 8722 15929 8756 15963
rect 5089 15861 5123 15895
rect 6285 15861 6319 15895
rect 7941 15861 7975 15895
rect 8309 15861 8343 15895
rect 9321 15861 9355 15895
rect 3249 15657 3283 15691
rect 3709 15657 3743 15691
rect 5825 15657 5859 15691
rect 1685 15589 1719 15623
rect 4813 15589 4847 15623
rect 6653 15589 6687 15623
rect 8033 15589 8067 15623
rect 5457 15521 5491 15555
rect 7941 15521 7975 15555
rect 8677 15521 8711 15555
rect 1593 15453 1627 15487
rect 6285 15453 6319 15487
rect 6561 15453 6595 15487
rect 6837 15453 6871 15487
rect 7481 15453 7515 15487
rect 2145 15385 2179 15419
rect 2605 15317 2639 15351
rect 2881 15317 2915 15351
rect 1685 15113 1719 15147
rect 2881 15113 2915 15147
rect 3525 15113 3559 15147
rect 4905 15113 4939 15147
rect 9597 15113 9631 15147
rect 2513 15045 2547 15079
rect 5825 15045 5859 15079
rect 1961 14977 1995 15011
rect 4353 14977 4387 15011
rect 6561 14977 6595 15011
rect 7113 14977 7147 15011
rect 7205 14909 7239 14943
rect 8217 14909 8251 14943
rect 8677 14909 8711 14943
rect 2053 14841 2087 14875
rect 3709 14841 3743 14875
rect 3801 14841 3835 14875
rect 5273 14841 5307 14875
rect 5365 14841 5399 14875
rect 8998 14841 9032 14875
rect 8493 14773 8527 14807
rect 4445 14569 4479 14603
rect 4997 14569 5031 14603
rect 5365 14569 5399 14603
rect 7205 14569 7239 14603
rect 10609 14569 10643 14603
rect 1777 14501 1811 14535
rect 2329 14501 2363 14535
rect 6187 14501 6221 14535
rect 8211 14501 8245 14535
rect 10010 14501 10044 14535
rect 6745 14433 6779 14467
rect 8769 14433 8803 14467
rect 1685 14365 1719 14399
rect 2973 14365 3007 14399
rect 4077 14365 4111 14399
rect 5825 14365 5859 14399
rect 7849 14365 7883 14399
rect 9689 14365 9723 14399
rect 5641 14297 5675 14331
rect 2605 14229 2639 14263
rect 3709 14229 3743 14263
rect 7757 14229 7791 14263
rect 9045 14229 9079 14263
rect 10885 14229 10919 14263
rect 1685 14025 1719 14059
rect 7849 14025 7883 14059
rect 11437 14025 11471 14059
rect 9873 13957 9907 13991
rect 2421 13889 2455 13923
rect 6285 13889 6319 13923
rect 3433 13821 3467 13855
rect 4261 13821 4295 13855
rect 6837 13821 6871 13855
rect 7389 13821 7423 13855
rect 8493 13821 8527 13855
rect 9045 13821 9079 13855
rect 9321 13821 9355 13855
rect 10333 13821 10367 13855
rect 10425 13821 10459 13855
rect 10885 13821 10919 13855
rect 2145 13753 2179 13787
rect 2237 13753 2271 13787
rect 3801 13753 3835 13787
rect 4169 13753 4203 13787
rect 4623 13753 4657 13787
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 5825 13685 5859 13719
rect 6653 13685 6687 13719
rect 6929 13685 6963 13719
rect 8401 13685 8435 13719
rect 8585 13685 8619 13719
rect 10517 13685 10551 13719
rect 1547 13481 1581 13515
rect 7665 13481 7699 13515
rect 10333 13481 10367 13515
rect 4261 13413 4295 13447
rect 6187 13413 6221 13447
rect 9045 13413 9079 13447
rect 10701 13413 10735 13447
rect 1476 13345 1510 13379
rect 2789 13345 2823 13379
rect 7573 13345 7607 13379
rect 8033 13345 8067 13379
rect 9689 13345 9723 13379
rect 11253 13345 11287 13379
rect 2421 13277 2455 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 5825 13277 5859 13311
rect 10057 13277 10091 13311
rect 12265 13277 12299 13311
rect 2145 13209 2179 13243
rect 6745 13209 6779 13243
rect 8677 13209 8711 13243
rect 11437 13209 11471 13243
rect 3893 13141 3927 13175
rect 7021 13141 7055 13175
rect 9413 13141 9447 13175
rect 9827 13141 9861 13175
rect 9965 13141 9999 13175
rect 1593 12937 1627 12971
rect 2237 12937 2271 12971
rect 3801 12937 3835 12971
rect 7941 12937 7975 12971
rect 9873 12937 9907 12971
rect 5089 12869 5123 12903
rect 2697 12801 2731 12835
rect 5917 12801 5951 12835
rect 6561 12801 6595 12835
rect 9413 12801 9447 12835
rect 9597 12801 9631 12835
rect 3960 12733 3994 12767
rect 4353 12733 4387 12767
rect 5181 12733 5215 12767
rect 5733 12733 5767 12767
rect 7021 12733 7055 12767
rect 8493 12733 8527 12767
rect 9321 12733 9355 12767
rect 10333 12733 10367 12767
rect 10609 12733 10643 12767
rect 11069 12733 11103 12767
rect 11253 12733 11287 12767
rect 12516 12733 12550 12767
rect 12909 12733 12943 12767
rect 2421 12665 2455 12699
rect 2513 12665 2547 12699
rect 6837 12665 6871 12699
rect 11897 12665 11931 12699
rect 3433 12597 3467 12631
rect 4031 12597 4065 12631
rect 6285 12597 6319 12631
rect 8401 12597 8435 12631
rect 10517 12597 10551 12631
rect 12587 12597 12621 12631
rect 1961 12393 1995 12427
rect 5273 12393 5307 12427
rect 6469 12393 6503 12427
rect 6653 12393 6687 12427
rect 11069 12393 11103 12427
rect 13001 12393 13035 12427
rect 2329 12325 2363 12359
rect 2605 12325 2639 12359
rect 4261 12325 4295 12359
rect 4813 12325 4847 12359
rect 5641 12325 5675 12359
rect 8033 12325 8067 12359
rect 8401 12325 8435 12359
rect 1476 12257 1510 12291
rect 6653 12257 6687 12291
rect 7021 12257 7055 12291
rect 8493 12257 8527 12291
rect 9229 12257 9263 12291
rect 10333 12257 10367 12291
rect 11713 12257 11747 12291
rect 12817 12257 12851 12291
rect 13829 12257 13863 12291
rect 2513 12189 2547 12223
rect 2789 12189 2823 12223
rect 4169 12189 4203 12223
rect 9689 12189 9723 12223
rect 11253 12189 11287 12223
rect 12541 12189 12575 12223
rect 13967 12189 14001 12223
rect 3433 12121 3467 12155
rect 9137 12121 9171 12155
rect 9229 12121 9263 12155
rect 1547 12053 1581 12087
rect 3893 12053 3927 12087
rect 7665 12053 7699 12087
rect 8677 12053 8711 12087
rect 9413 12053 9447 12087
rect 10793 12053 10827 12087
rect 13277 12053 13311 12087
rect 3157 11849 3191 11883
rect 4261 11849 4295 11883
rect 5917 11849 5951 11883
rect 8125 11849 8159 11883
rect 13645 11849 13679 11883
rect 13829 11849 13863 11883
rect 2789 11781 2823 11815
rect 7757 11781 7791 11815
rect 10793 11781 10827 11815
rect 12265 11781 12299 11815
rect 12725 11781 12759 11815
rect 13461 11781 13495 11815
rect 1777 11713 1811 11747
rect 2421 11713 2455 11747
rect 3617 11713 3651 11747
rect 5181 11713 5215 11747
rect 6285 11713 6319 11747
rect 6837 11713 6871 11747
rect 9781 11713 9815 11747
rect 10885 11713 10919 11747
rect 12081 11713 12115 11747
rect 12596 11713 12630 11747
rect 12817 11713 12851 11747
rect 8493 11645 8527 11679
rect 8861 11645 8895 11679
rect 9413 11645 9447 11679
rect 9597 11645 9631 11679
rect 1869 11577 1903 11611
rect 3341 11577 3375 11611
rect 3433 11577 3467 11611
rect 4905 11577 4939 11611
rect 4997 11577 5031 11611
rect 7158 11577 7192 11611
rect 10517 11645 10551 11679
rect 10664 11645 10698 11679
rect 11253 11577 11287 11611
rect 12449 11645 12483 11679
rect 14064 11645 14098 11679
rect 14473 11645 14507 11679
rect 14151 11577 14185 11611
rect 15025 11577 15059 11611
rect 4721 11509 4755 11543
rect 6561 11509 6595 11543
rect 8677 11509 8711 11543
rect 9781 11509 9815 11543
rect 10057 11509 10091 11543
rect 10425 11509 10459 11543
rect 11805 11509 11839 11543
rect 12081 11509 12115 11543
rect 13093 11509 13127 11543
rect 13645 11509 13679 11543
rect 1593 11305 1627 11339
rect 3617 11305 3651 11339
rect 4721 11305 4755 11339
rect 5181 11305 5215 11339
rect 5733 11305 5767 11339
rect 8033 11305 8067 11339
rect 10149 11305 10183 11339
rect 11989 11305 12023 11339
rect 12357 11305 12391 11339
rect 2053 11237 2087 11271
rect 2605 11237 2639 11271
rect 6974 11237 7008 11271
rect 9505 11237 9539 11271
rect 7573 11169 7607 11203
rect 8585 11169 8619 11203
rect 9965 11169 9999 11203
rect 10609 11169 10643 11203
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 13185 11169 13219 11203
rect 14105 11169 14139 11203
rect 15368 11169 15402 11203
rect 1961 11101 1995 11135
rect 4813 11101 4847 11135
rect 6653 11101 6687 11135
rect 8401 11101 8435 11135
rect 11713 11101 11747 11135
rect 12541 11101 12575 11135
rect 6561 11033 6595 11067
rect 8769 11033 8803 11067
rect 15439 11033 15473 11067
rect 2881 10965 2915 10999
rect 3341 10965 3375 10999
rect 9137 10965 9171 10999
rect 14243 10965 14277 10999
rect 3433 10761 3467 10795
rect 10425 10761 10459 10795
rect 11069 10761 11103 10795
rect 13645 10761 13679 10795
rect 3157 10693 3191 10727
rect 9505 10693 9539 10727
rect 10241 10693 10275 10727
rect 14657 10693 14691 10727
rect 2789 10625 2823 10659
rect 6285 10625 6319 10659
rect 10333 10625 10367 10659
rect 11345 10625 11379 10659
rect 3652 10557 3686 10591
rect 4077 10557 4111 10591
rect 4537 10557 4571 10591
rect 4997 10557 5031 10591
rect 7113 10557 7147 10591
rect 7389 10557 7423 10591
rect 8401 10557 8435 10591
rect 8861 10557 8895 10591
rect 10112 10557 10146 10591
rect 12265 10557 12299 10591
rect 12725 10557 12759 10591
rect 14197 10557 14231 10591
rect 15025 10557 15059 10591
rect 15244 10557 15278 10591
rect 15669 10557 15703 10591
rect 16256 10557 16290 10591
rect 16681 10557 16715 10591
rect 2145 10489 2179 10523
rect 2237 10489 2271 10523
rect 5318 10489 5352 10523
rect 6561 10489 6595 10523
rect 9965 10489 9999 10523
rect 16037 10489 16071 10523
rect 1961 10421 1995 10455
rect 3755 10421 3789 10455
rect 4813 10421 4847 10455
rect 5917 10421 5951 10455
rect 6929 10421 6963 10455
rect 8033 10421 8067 10455
rect 8493 10421 8527 10455
rect 11713 10421 11747 10455
rect 12909 10421 12943 10455
rect 14381 10421 14415 10455
rect 15347 10421 15381 10455
rect 16359 10421 16393 10455
rect 2697 10217 2731 10251
rect 4215 10217 4249 10251
rect 4721 10217 4755 10251
rect 5365 10217 5399 10251
rect 6745 10217 6779 10251
rect 9137 10217 9171 10251
rect 11161 10217 11195 10251
rect 1777 10149 1811 10183
rect 8769 10149 8803 10183
rect 3893 10081 3927 10115
rect 4123 10081 4157 10115
rect 5273 10081 5307 10115
rect 5825 10081 5859 10115
rect 8033 10081 8067 10115
rect 10149 10081 10183 10115
rect 11437 10081 11471 10115
rect 11805 10081 11839 10115
rect 13093 10081 13127 10115
rect 13277 10081 13311 10115
rect 16380 10081 16414 10115
rect 1685 10013 1719 10047
rect 6837 10013 6871 10047
rect 7849 10013 7883 10047
rect 8401 10013 8435 10047
rect 9689 10013 9723 10047
rect 11989 10013 12023 10047
rect 13553 10013 13587 10047
rect 15301 10013 15335 10047
rect 2237 9945 2271 9979
rect 2973 9945 3007 9979
rect 4997 9877 5031 9911
rect 7573 9877 7607 9911
rect 8171 9877 8205 9911
rect 8309 9877 8343 9911
rect 9505 9877 9539 9911
rect 10793 9877 10827 9911
rect 12541 9877 12575 9911
rect 16451 9877 16485 9911
rect 5089 9673 5123 9707
rect 8861 9673 8895 9707
rect 10609 9673 10643 9707
rect 11621 9673 11655 9707
rect 13277 9673 13311 9707
rect 3157 9605 3191 9639
rect 8539 9605 8573 9639
rect 8677 9605 8711 9639
rect 2145 9537 2179 9571
rect 2421 9537 2455 9571
rect 7573 9537 7607 9571
rect 8125 9537 8159 9571
rect 8769 9537 8803 9571
rect 10425 9537 10459 9571
rect 3617 9469 3651 9503
rect 4169 9469 4203 9503
rect 4721 9469 4755 9503
rect 5825 9469 5859 9503
rect 6653 9469 6687 9503
rect 7481 9469 7515 9503
rect 8401 9469 8435 9503
rect 10793 9469 10827 9503
rect 11253 9469 11287 9503
rect 12449 9469 12483 9503
rect 12909 9469 12943 9503
rect 2237 9401 2271 9435
rect 5181 9401 5215 9435
rect 13185 9401 13219 9435
rect 13829 9605 13863 9639
rect 14013 9537 14047 9571
rect 14105 9469 14139 9503
rect 15485 9469 15519 9503
rect 15669 9469 15703 9503
rect 15577 9401 15611 9435
rect 1593 9333 1627 9367
rect 3433 9333 3467 9367
rect 3893 9333 3927 9367
rect 9781 9333 9815 9367
rect 11989 9333 12023 9367
rect 13277 9333 13311 9367
rect 13553 9333 13587 9367
rect 16589 9333 16623 9367
rect 5365 9129 5399 9163
rect 7573 9129 7607 9163
rect 7941 9129 7975 9163
rect 8861 9129 8895 9163
rect 9137 9129 9171 9163
rect 10793 9129 10827 9163
rect 2329 9061 2363 9095
rect 2421 9061 2455 9095
rect 4439 9061 4473 9095
rect 6009 9061 6043 9095
rect 12909 9061 12943 9095
rect 15485 9061 15519 9095
rect 4077 8993 4111 9027
rect 8677 8993 8711 9027
rect 8861 8993 8895 9027
rect 9689 8993 9723 9027
rect 11437 8993 11471 9027
rect 16865 8993 16899 9027
rect 17944 8993 17978 9027
rect 18924 8993 18958 9027
rect 2605 8925 2639 8959
rect 5641 8925 5675 8959
rect 5917 8925 5951 8959
rect 8769 8925 8803 8959
rect 12817 8925 12851 8959
rect 13461 8925 13495 8959
rect 15393 8925 15427 8959
rect 16037 8925 16071 8959
rect 19349 8925 19383 8959
rect 3709 8857 3743 8891
rect 6469 8857 6503 8891
rect 9873 8857 9907 8891
rect 11161 8857 11195 8891
rect 1777 8789 1811 8823
rect 2145 8789 2179 8823
rect 3249 8789 3283 8823
rect 4997 8789 5031 8823
rect 12449 8789 12483 8823
rect 14013 8789 14047 8823
rect 17049 8789 17083 8823
rect 18015 8789 18049 8823
rect 19027 8789 19061 8823
rect 6285 8585 6319 8619
rect 6561 8585 6595 8619
rect 8125 8585 8159 8619
rect 9413 8585 9447 8619
rect 10057 8585 10091 8619
rect 13369 8585 13403 8619
rect 15117 8585 15151 8619
rect 15485 8585 15519 8619
rect 16957 8585 16991 8619
rect 18245 8585 18279 8619
rect 18521 8585 18555 8619
rect 2329 8517 2363 8551
rect 8447 8517 8481 8551
rect 8585 8517 8619 8551
rect 19211 8517 19245 8551
rect 5549 8449 5583 8483
rect 6837 8449 6871 8483
rect 7757 8449 7791 8483
rect 8677 8449 8711 8483
rect 8769 8449 8803 8483
rect 9781 8449 9815 8483
rect 3249 8381 3283 8415
rect 10793 8381 10827 8415
rect 11345 8381 11379 8415
rect 11529 8381 11563 8415
rect 12449 8381 12483 8415
rect 13645 8381 13679 8415
rect 14197 8381 14231 8415
rect 15853 8381 15887 8415
rect 16037 8381 16071 8415
rect 18061 8381 18095 8415
rect 18889 8381 18923 8415
rect 19119 8381 19153 8415
rect 19533 8381 19567 8415
rect 1777 8313 1811 8347
rect 1869 8313 1903 8347
rect 3065 8313 3099 8347
rect 3611 8313 3645 8347
rect 5273 8313 5307 8347
rect 5365 8313 5399 8347
rect 8309 8313 8343 8347
rect 11805 8313 11839 8347
rect 12265 8313 12299 8347
rect 12770 8313 12804 8347
rect 14105 8313 14139 8347
rect 14518 8313 14552 8347
rect 15945 8313 15979 8347
rect 2697 8245 2731 8279
rect 4169 8245 4203 8279
rect 4537 8245 4571 8279
rect 5089 8245 5123 8279
rect 7389 8245 7423 8279
rect 10701 8245 10735 8279
rect 1961 8041 1995 8075
rect 3893 8041 3927 8075
rect 4169 8041 4203 8075
rect 5273 8041 5307 8075
rect 8677 8041 8711 8075
rect 12449 8041 12483 8075
rect 12817 8041 12851 8075
rect 13921 8041 13955 8075
rect 14289 8041 14323 8075
rect 19119 8041 19153 8075
rect 3157 7973 3191 8007
rect 6095 7973 6129 8007
rect 10609 7973 10643 8007
rect 11437 7973 11471 8007
rect 13093 7973 13127 8007
rect 13645 7973 13679 8007
rect 15393 7973 15427 8007
rect 15485 7973 15519 8007
rect 1409 7905 1443 7939
rect 2697 7905 2731 7939
rect 2973 7905 3007 7939
rect 4353 7905 4387 7939
rect 4629 7905 4663 7939
rect 7021 7905 7055 7939
rect 9137 7905 9171 7939
rect 9505 7905 9539 7939
rect 9873 7905 9907 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 11253 7905 11287 7939
rect 11621 7905 11655 7939
rect 17969 7905 18003 7939
rect 19016 7905 19050 7939
rect 23648 7905 23682 7939
rect 1547 7837 1581 7871
rect 3433 7837 3467 7871
rect 5733 7837 5767 7871
rect 7941 7837 7975 7871
rect 8401 7837 8435 7871
rect 10020 7837 10054 7871
rect 10241 7837 10275 7871
rect 6653 7769 6687 7803
rect 11989 7837 12023 7871
rect 13001 7837 13035 7871
rect 15025 7837 15059 7871
rect 16037 7837 16071 7871
rect 18153 7837 18187 7871
rect 2237 7701 2271 7735
rect 5549 7701 5583 7735
rect 7573 7701 7607 7735
rect 8171 7701 8205 7735
rect 8309 7701 8343 7735
rect 10149 7701 10183 7735
rect 10793 7701 10827 7735
rect 23719 7701 23753 7735
rect 2973 7497 3007 7531
rect 4721 7497 4755 7531
rect 5089 7497 5123 7531
rect 6653 7497 6687 7531
rect 7941 7497 7975 7531
rect 10130 7497 10164 7531
rect 11069 7497 11103 7531
rect 12173 7497 12207 7531
rect 12725 7497 12759 7531
rect 15301 7497 15335 7531
rect 2697 7429 2731 7463
rect 8677 7429 8711 7463
rect 9229 7429 9263 7463
rect 10241 7429 10275 7463
rect 13645 7429 13679 7463
rect 16773 7429 16807 7463
rect 1593 7361 1627 7395
rect 4353 7361 4387 7395
rect 5917 7361 5951 7395
rect 7205 7361 7239 7395
rect 8309 7361 8343 7395
rect 8769 7361 8803 7395
rect 1961 7293 1995 7327
rect 3617 7293 3651 7327
rect 4169 7293 4203 7327
rect 8548 7293 8582 7327
rect 5273 7225 5307 7259
rect 5365 7225 5399 7259
rect 6929 7225 6963 7259
rect 7021 7225 7055 7259
rect 8401 7225 8435 7259
rect 10333 7361 10367 7395
rect 9965 7293 9999 7327
rect 12817 7293 12851 7327
rect 13829 7293 13863 7327
rect 14381 7293 14415 7327
rect 15393 7293 15427 7327
rect 15945 7293 15979 7327
rect 16405 7293 16439 7327
rect 16957 7293 16991 7327
rect 17417 7293 17451 7327
rect 18153 7293 18187 7327
rect 19660 7293 19694 7327
rect 20085 7293 20119 7327
rect 20688 7293 20722 7327
rect 21716 7293 21750 7327
rect 22109 7293 22143 7327
rect 10701 7225 10735 7259
rect 11529 7225 11563 7259
rect 14565 7225 14599 7259
rect 16129 7225 16163 7259
rect 18061 7225 18095 7259
rect 20775 7225 20809 7259
rect 3433 7157 3467 7191
rect 6193 7157 6227 7191
rect 9045 7157 9079 7191
rect 9229 7157 9263 7191
rect 9505 7157 9539 7191
rect 9873 7157 9907 7191
rect 11897 7157 11931 7191
rect 13001 7157 13035 7191
rect 13369 7157 13403 7191
rect 14841 7157 14875 7191
rect 17141 7157 17175 7191
rect 17877 7157 17911 7191
rect 19073 7157 19107 7191
rect 19763 7157 19797 7191
rect 21097 7157 21131 7191
rect 21787 7157 21821 7191
rect 23857 7157 23891 7191
rect 3065 6953 3099 6987
rect 6377 6953 6411 6987
rect 7573 6953 7607 6987
rect 9137 6953 9171 6987
rect 9413 6953 9447 6987
rect 10333 6953 10367 6987
rect 12725 6953 12759 6987
rect 13093 6953 13127 6987
rect 16221 6953 16255 6987
rect 17417 6953 17451 6987
rect 17969 6953 18003 6987
rect 18245 6953 18279 6987
rect 2053 6885 2087 6919
rect 2145 6885 2179 6919
rect 5819 6885 5853 6919
rect 8033 6885 8067 6919
rect 9689 6885 9723 6919
rect 15622 6885 15656 6919
rect 18981 6885 19015 6919
rect 2697 6817 2731 6851
rect 4112 6817 4146 6851
rect 7205 6817 7239 6851
rect 8180 6817 8214 6851
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 12357 6817 12391 6851
rect 13645 6817 13679 6851
rect 14105 6817 14139 6851
rect 17049 6817 17083 6851
rect 20821 6817 20855 6851
rect 21960 6817 21994 6851
rect 24593 6817 24627 6851
rect 5457 6749 5491 6783
rect 8401 6749 8435 6783
rect 10057 6749 10091 6783
rect 11621 6749 11655 6783
rect 11989 6749 12023 6783
rect 14289 6749 14323 6783
rect 15301 6749 15335 6783
rect 18889 6749 18923 6783
rect 21051 6749 21085 6783
rect 3709 6681 3743 6715
rect 4629 6681 4663 6715
rect 8493 6681 8527 6715
rect 9854 6681 9888 6715
rect 11391 6681 11425 6715
rect 19441 6681 19475 6715
rect 1593 6613 1627 6647
rect 4215 6613 4249 6647
rect 4905 6613 4939 6647
rect 6837 6613 6871 6647
rect 7941 6613 7975 6647
rect 8309 6613 8343 6647
rect 9965 6613 9999 6647
rect 10793 6613 10827 6647
rect 11529 6613 11563 6647
rect 22063 6613 22097 6647
rect 24777 6613 24811 6647
rect 2421 6409 2455 6443
rect 2697 6409 2731 6443
rect 4353 6409 4387 6443
rect 5825 6409 5859 6443
rect 7389 6409 7423 6443
rect 8474 6409 8508 6443
rect 10038 6409 10072 6443
rect 11713 6409 11747 6443
rect 13461 6409 13495 6443
rect 14197 6409 14231 6443
rect 16221 6409 16255 6443
rect 16773 6409 16807 6443
rect 17877 6409 17911 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 22017 6409 22051 6443
rect 24593 6409 24627 6443
rect 2237 6341 2271 6375
rect 1685 6273 1719 6307
rect 7757 6341 7791 6375
rect 8585 6341 8619 6375
rect 10149 6341 10183 6375
rect 3157 6273 3191 6307
rect 8677 6273 8711 6307
rect 10241 6273 10275 6307
rect 12541 6273 12575 6307
rect 13921 6273 13955 6307
rect 15301 6273 15335 6307
rect 16957 6273 16991 6307
rect 18797 6273 18831 6307
rect 4905 6205 4939 6239
rect 8125 6205 8159 6239
rect 9413 6205 9447 6239
rect 9781 6205 9815 6239
rect 14013 6205 14047 6239
rect 15025 6205 15059 6239
rect 19993 6205 20027 6239
rect 21256 6205 21290 6239
rect 21649 6205 21683 6239
rect 22236 6205 22270 6239
rect 22661 6205 22695 6239
rect 23740 6205 23774 6239
rect 24133 6205 24167 6239
rect 1777 6137 1811 6171
rect 2421 6137 2455 6171
rect 3065 6137 3099 6171
rect 3519 6137 3553 6171
rect 5267 6137 5301 6171
rect 6469 6137 6503 6171
rect 8309 6137 8343 6171
rect 9873 6137 9907 6171
rect 12265 6137 12299 6171
rect 12633 6137 12667 6171
rect 13185 6137 13219 6171
rect 14749 6137 14783 6171
rect 15393 6137 15427 6171
rect 15945 6137 15979 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 19625 6137 19659 6171
rect 22339 6137 22373 6171
rect 4077 6069 4111 6103
rect 4813 6069 4847 6103
rect 6193 6069 6227 6103
rect 6837 6069 6871 6103
rect 8953 6069 8987 6103
rect 10517 6069 10551 6103
rect 10977 6069 11011 6103
rect 11345 6069 11379 6103
rect 17417 6069 17451 6103
rect 20913 6069 20947 6103
rect 21327 6069 21361 6103
rect 23811 6069 23845 6103
rect 2513 5865 2547 5899
rect 4537 5865 4571 5899
rect 5457 5865 5491 5899
rect 7021 5865 7055 5899
rect 8401 5865 8435 5899
rect 10793 5865 10827 5899
rect 11621 5865 11655 5899
rect 13461 5865 13495 5899
rect 15117 5865 15151 5899
rect 15853 5865 15887 5899
rect 16865 5865 16899 5899
rect 17417 5865 17451 5899
rect 18153 5865 18187 5899
rect 19717 5865 19751 5899
rect 1685 5797 1719 5831
rect 2237 5797 2271 5831
rect 3249 5797 3283 5831
rect 9689 5797 9723 5831
rect 11253 5797 11287 5831
rect 12126 5797 12160 5831
rect 18429 5797 18463 5831
rect 23627 5797 23661 5831
rect 4144 5729 4178 5763
rect 5365 5729 5399 5763
rect 5917 5729 5951 5763
rect 7205 5729 7239 5763
rect 7481 5729 7515 5763
rect 9505 5729 9539 5763
rect 11805 5729 11839 5763
rect 13093 5729 13127 5763
rect 13645 5729 13679 5763
rect 14105 5729 14139 5763
rect 15301 5729 15335 5763
rect 18981 5729 19015 5763
rect 21005 5729 21039 5763
rect 22477 5729 22511 5763
rect 23524 5729 23558 5763
rect 1593 5661 1627 5695
rect 8493 5661 8527 5695
rect 9045 5661 9079 5695
rect 9836 5661 9870 5695
rect 10057 5661 10091 5695
rect 14381 5661 14415 5695
rect 16497 5661 16531 5695
rect 18337 5661 18371 5695
rect 19809 5661 19843 5695
rect 3525 5593 3559 5627
rect 4215 5593 4249 5627
rect 12725 5593 12759 5627
rect 5273 5525 5307 5559
rect 8033 5525 8067 5559
rect 9965 5525 9999 5559
rect 10149 5525 10183 5559
rect 15485 5525 15519 5559
rect 21189 5525 21223 5559
rect 22615 5525 22649 5559
rect 7941 5321 7975 5355
rect 9873 5321 9907 5355
rect 17877 5321 17911 5355
rect 19073 5321 19107 5355
rect 20729 5321 20763 5355
rect 4445 5253 4479 5287
rect 5089 5253 5123 5287
rect 6653 5253 6687 5287
rect 11345 5253 11379 5287
rect 13645 5253 13679 5287
rect 15117 5253 15151 5287
rect 24133 5253 24167 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 6285 5185 6319 5219
rect 8677 5185 8711 5219
rect 10241 5185 10275 5219
rect 12541 5185 12575 5219
rect 13185 5185 13219 5219
rect 15301 5185 15335 5219
rect 15945 5185 15979 5219
rect 18153 5185 18187 5219
rect 18797 5185 18831 5219
rect 21189 5185 21223 5219
rect 3341 5117 3375 5151
rect 3433 5117 3467 5151
rect 3893 5117 3927 5151
rect 5181 5117 5215 5151
rect 5733 5117 5767 5151
rect 7113 5117 7147 5151
rect 7389 5117 7423 5151
rect 9045 5117 9079 5151
rect 9321 5117 9355 5151
rect 10609 5117 10643 5151
rect 10793 5117 10827 5151
rect 14013 5117 14047 5151
rect 16957 5117 16991 5151
rect 19717 5117 19751 5151
rect 21097 5117 21131 5151
rect 21281 5117 21315 5151
rect 23949 5117 23983 5151
rect 24501 5117 24535 5151
rect 25120 5117 25154 5151
rect 1777 5049 1811 5083
rect 2697 5049 2731 5083
rect 4169 5049 4203 5083
rect 8309 5049 8343 5083
rect 9505 5049 9539 5083
rect 11069 5049 11103 5083
rect 12633 5049 12667 5083
rect 14565 5049 14599 5083
rect 15393 5049 15427 5083
rect 18245 5049 18279 5083
rect 19625 5049 19659 5083
rect 23397 5049 23431 5083
rect 5273 4981 5307 5015
rect 6929 4981 6963 5015
rect 11897 4981 11931 5015
rect 12265 4981 12299 5015
rect 14197 4981 14231 5015
rect 16497 4981 16531 5015
rect 19441 4981 19475 5015
rect 22477 4981 22511 5015
rect 25191 4981 25225 5015
rect 25513 4981 25547 5015
rect 1685 4777 1719 4811
rect 2053 4777 2087 4811
rect 3525 4777 3559 4811
rect 5365 4777 5399 4811
rect 5825 4777 5859 4811
rect 7849 4777 7883 4811
rect 9045 4777 9079 4811
rect 9413 4777 9447 4811
rect 10701 4777 10735 4811
rect 11805 4777 11839 4811
rect 12265 4777 12299 4811
rect 18705 4777 18739 4811
rect 2145 4709 2179 4743
rect 4439 4709 4473 4743
rect 6330 4709 6364 4743
rect 9781 4709 9815 4743
rect 9873 4709 9907 4743
rect 11161 4709 11195 4743
rect 12541 4709 12575 4743
rect 13645 4709 13679 4743
rect 15622 4709 15656 4743
rect 16497 4709 16531 4743
rect 18153 4709 18187 4743
rect 18521 4709 18555 4743
rect 2789 4641 2823 4675
rect 4077 4641 4111 4675
rect 6009 4641 6043 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 8309 4641 8343 4675
rect 13921 4641 13955 4675
rect 15301 4641 15335 4675
rect 16221 4641 16255 4675
rect 17141 4641 17175 4675
rect 18613 4641 18647 4675
rect 19073 4641 19107 4675
rect 21005 4641 21039 4675
rect 22569 4641 22603 4675
rect 23708 4641 23742 4675
rect 24720 4641 24754 4675
rect 10057 4573 10091 4607
rect 11253 4573 11287 4607
rect 12449 4573 12483 4607
rect 20913 4573 20947 4607
rect 24823 4573 24857 4607
rect 13001 4505 13035 4539
rect 22753 4505 22787 4539
rect 3893 4437 3927 4471
rect 4997 4437 5031 4471
rect 6929 4437 6963 4471
rect 14105 4437 14139 4471
rect 15117 4437 15151 4471
rect 17325 4437 17359 4471
rect 23811 4437 23845 4471
rect 1777 4233 1811 4267
rect 6653 4233 6687 4267
rect 7113 4233 7147 4267
rect 8677 4233 8711 4267
rect 18981 4233 19015 4267
rect 22569 4233 22603 4267
rect 24823 4233 24857 4267
rect 25513 4233 25547 4267
rect 10885 4165 10919 4199
rect 14289 4165 14323 4199
rect 17785 4165 17819 4199
rect 2789 4097 2823 4131
rect 3249 4097 3283 4131
rect 11437 4097 11471 4131
rect 12449 4097 12483 4131
rect 15485 4097 15519 4131
rect 16681 4097 16715 4131
rect 19257 4097 19291 4131
rect 2053 4029 2087 4063
rect 5457 4029 5491 4063
rect 5641 4029 5675 4063
rect 7481 4029 7515 4063
rect 7849 4029 7883 4063
rect 8125 4029 8159 4063
rect 8309 4029 8343 4063
rect 9137 4029 9171 4063
rect 10977 4029 11011 4063
rect 11161 4029 11195 4063
rect 18061 4029 18095 4063
rect 19809 4029 19843 4063
rect 19901 4029 19935 4063
rect 21465 4029 21499 4063
rect 23740 4029 23774 4063
rect 24133 4029 24167 4063
rect 24720 4029 24754 4063
rect 25145 4029 25179 4063
rect 3157 3961 3191 3995
rect 3611 3961 3645 3995
rect 5089 3961 5123 3995
rect 5917 3961 5951 3995
rect 9499 3961 9533 3995
rect 11897 3961 11931 3995
rect 12265 3961 12299 3995
rect 12811 3961 12845 3995
rect 15025 3961 15059 3995
rect 15393 3961 15427 3995
rect 15847 3961 15881 3995
rect 18382 3961 18416 3995
rect 19625 3961 19659 3995
rect 21373 3961 21407 3995
rect 24501 3961 24535 3995
rect 4169 3893 4203 3927
rect 4537 3893 4571 3927
rect 6193 3893 6227 3927
rect 9045 3893 9079 3927
rect 10057 3893 10091 3927
rect 10333 3893 10367 3927
rect 13369 3893 13403 3927
rect 14013 3893 14047 3927
rect 14473 3893 14507 3927
rect 16405 3893 16439 3927
rect 17049 3893 17083 3927
rect 17417 3893 17451 3927
rect 20821 3893 20855 3927
rect 21189 3893 21223 3927
rect 23811 3893 23845 3927
rect 1547 3689 1581 3723
rect 1961 3689 1995 3723
rect 2329 3689 2363 3723
rect 3525 3689 3559 3723
rect 3801 3689 3835 3723
rect 5273 3689 5307 3723
rect 7665 3689 7699 3723
rect 9137 3689 9171 3723
rect 11161 3689 11195 3723
rect 12449 3689 12483 3723
rect 14289 3689 14323 3723
rect 15025 3689 15059 3723
rect 18061 3689 18095 3723
rect 18705 3689 18739 3723
rect 2605 3621 2639 3655
rect 4169 3621 4203 3655
rect 4261 3621 4295 3655
rect 4813 3621 4847 3655
rect 6003 3621 6037 3655
rect 8211 3621 8245 3655
rect 9781 3621 9815 3655
rect 9873 3621 9907 3655
rect 11713 3621 11747 3655
rect 1476 3553 1510 3587
rect 2513 3485 2547 3519
rect 5641 3485 5675 3519
rect 7849 3485 7883 3519
rect 11621 3485 11655 3519
rect 12265 3485 12299 3519
rect 13185 3621 13219 3655
rect 13277 3621 13311 3655
rect 15669 3621 15703 3655
rect 17233 3621 17267 3655
rect 18981 3621 19015 3655
rect 21005 3553 21039 3587
rect 22569 3553 22603 3587
rect 24225 3553 24259 3587
rect 13461 3485 13495 3519
rect 14749 3485 14783 3519
rect 15577 3485 15611 3519
rect 16221 3485 16255 3519
rect 17141 3485 17175 3519
rect 17417 3485 17451 3519
rect 18889 3485 18923 3519
rect 19165 3485 19199 3519
rect 20913 3485 20947 3519
rect 22477 3485 22511 3519
rect 24041 3485 24075 3519
rect 3065 3417 3099 3451
rect 7297 3417 7331 3451
rect 10333 3417 10367 3451
rect 12449 3417 12483 3451
rect 6561 3349 6595 3383
rect 6837 3349 6871 3383
rect 8769 3349 8803 3383
rect 10701 3349 10735 3383
rect 12633 3349 12667 3383
rect 12909 3349 12943 3383
rect 19809 3349 19843 3383
rect 1685 3145 1719 3179
rect 4307 3145 4341 3179
rect 6653 3145 6687 3179
rect 9505 3145 9539 3179
rect 9781 3145 9815 3179
rect 14197 3145 14231 3179
rect 15577 3145 15611 3179
rect 19073 3145 19107 3179
rect 19257 3145 19291 3179
rect 20821 3145 20855 3179
rect 24225 3145 24259 3179
rect 24915 3145 24949 3179
rect 3065 3077 3099 3111
rect 3801 3077 3835 3111
rect 7941 3077 7975 3111
rect 8309 3077 8343 3111
rect 17233 3077 17267 3111
rect 2513 3009 2547 3043
rect 5273 3009 5307 3043
rect 6285 3009 6319 3043
rect 6929 3009 6963 3043
rect 8493 3009 8527 3043
rect 9965 3009 9999 3043
rect 11253 3009 11287 3043
rect 13461 3009 13495 3043
rect 14289 3009 14323 3043
rect 16221 3009 16255 3043
rect 16497 3009 16531 3043
rect 18337 3009 18371 3043
rect 18981 3009 19015 3043
rect 19901 3077 19935 3111
rect 1476 2941 1510 2975
rect 4236 2941 4270 2975
rect 5917 2941 5951 2975
rect 15209 2941 15243 2975
rect 19073 2941 19107 2975
rect 19809 2941 19843 2975
rect 20361 2941 20395 2975
rect 21465 2941 21499 2975
rect 23397 2941 23431 2975
rect 23673 2941 23707 2975
rect 24844 2941 24878 2975
rect 25237 2941 25271 2975
rect 1961 2873 1995 2907
rect 2605 2873 2639 2907
rect 5089 2873 5123 2907
rect 5365 2873 5399 2907
rect 7021 2873 7055 2907
rect 7573 2873 7607 2907
rect 8585 2873 8619 2907
rect 9137 2873 9171 2907
rect 10327 2873 10361 2907
rect 12817 2873 12851 2907
rect 12909 2873 12943 2907
rect 14610 2873 14644 2907
rect 16313 2873 16347 2907
rect 18429 2873 18463 2907
rect 19625 2873 19659 2907
rect 21373 2873 21407 2907
rect 22477 2873 22511 2907
rect 2329 2805 2363 2839
rect 3525 2805 3559 2839
rect 4721 2805 4755 2839
rect 10885 2805 10919 2839
rect 11621 2805 11655 2839
rect 11897 2805 11931 2839
rect 13829 2805 13863 2839
rect 16037 2805 16071 2839
rect 17877 2805 17911 2839
rect 21189 2805 21223 2839
rect 23857 2805 23891 2839
rect 1547 2601 1581 2635
rect 4399 2601 4433 2635
rect 6285 2601 6319 2635
rect 7941 2601 7975 2635
rect 8631 2601 8665 2635
rect 10793 2601 10827 2635
rect 11161 2601 11195 2635
rect 11345 2601 11379 2635
rect 14013 2601 14047 2635
rect 15301 2601 15335 2635
rect 17693 2601 17727 2635
rect 19349 2601 19383 2635
rect 2329 2533 2363 2567
rect 2605 2533 2639 2567
rect 3157 2533 3191 2567
rect 5181 2533 5215 2567
rect 5457 2533 5491 2567
rect 6745 2533 6779 2567
rect 7113 2533 7147 2567
rect 9597 2533 9631 2567
rect 9965 2533 9999 2567
rect 12357 2533 12391 2567
rect 12817 2533 12851 2567
rect 16589 2533 16623 2567
rect 16865 2533 16899 2567
rect 18521 2533 18555 2567
rect 21189 2533 21223 2567
rect 1476 2465 1510 2499
rect 3893 2465 3927 2499
rect 4328 2465 4362 2499
rect 6009 2465 6043 2499
rect 8560 2465 8594 2499
rect 8953 2465 8987 2499
rect 14933 2465 14967 2499
rect 15577 2465 15611 2499
rect 17417 2465 17451 2499
rect 19073 2465 19107 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21281 2465 21315 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 25697 2465 25731 2499
rect 2513 2397 2547 2431
rect 3525 2397 3559 2431
rect 5365 2397 5399 2431
rect 7021 2397 7055 2431
rect 7665 2397 7699 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 14381 2397 14415 2431
rect 16129 2397 16163 2431
rect 16773 2397 16807 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 20913 2397 20947 2431
rect 4813 2329 4847 2363
rect 13645 2329 13679 2363
rect 20085 2329 20119 2363
rect 24225 2329 24259 2363
rect 1869 2261 1903 2295
rect 8309 2261 8343 2295
rect 12081 2261 12115 2295
rect 15761 2261 15795 2295
rect 19717 2261 19751 2295
rect 22937 2261 22971 2295
rect 25329 2261 25363 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1578 24392 1584 24404
rect 1539 24364 1584 24392
rect 1578 24352 1584 24364
rect 1636 24352 1642 24404
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 1486 24256 1492 24268
rect 1443 24228 1492 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 1486 24216 1492 24228
rect 1544 24216 1550 24268
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1118 23808 1124 23860
rect 1176 23848 1182 23860
rect 1581 23851 1639 23857
rect 1581 23848 1593 23851
rect 1176 23820 1593 23848
rect 1176 23808 1182 23820
rect 1581 23817 1593 23820
rect 1627 23817 1639 23851
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 1581 23811 1639 23817
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 1486 23672 1492 23724
rect 1544 23712 1550 23724
rect 2041 23715 2099 23721
rect 2041 23712 2053 23715
rect 1544 23684 2053 23712
rect 1544 23672 1550 23684
rect 2041 23681 2053 23684
rect 2087 23712 2099 23715
rect 3418 23712 3424 23724
rect 2087 23684 3424 23712
rect 2087 23681 2099 23684
rect 2041 23675 2099 23681
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 1394 23644 1400 23656
rect 1355 23616 1400 23644
rect 1394 23604 1400 23616
rect 1452 23604 1458 23656
rect 2501 23647 2559 23653
rect 2501 23613 2513 23647
rect 2547 23644 2559 23647
rect 2547 23616 3188 23644
rect 2547 23613 2559 23616
rect 2501 23607 2559 23613
rect 3160 23517 3188 23616
rect 3145 23511 3203 23517
rect 3145 23477 3157 23511
rect 3191 23508 3203 23511
rect 4890 23508 4896 23520
rect 3191 23480 4896 23508
rect 3191 23477 3203 23480
rect 3145 23471 3203 23477
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1394 22924 1400 22976
rect 1452 22964 1458 22976
rect 1673 22967 1731 22973
rect 1673 22964 1685 22967
rect 1452 22936 1685 22964
rect 1452 22924 1458 22936
rect 1673 22933 1685 22936
rect 1719 22964 1731 22967
rect 1946 22964 1952 22976
rect 1719 22936 1952 22964
rect 1719 22933 1731 22936
rect 1673 22927 1731 22933
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 2084 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2056 21344 2084 21440
rect 2038 21332 2044 21344
rect 1999 21304 2044 21332
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1486 21088 1492 21140
rect 1544 21128 1550 21140
rect 1581 21131 1639 21137
rect 1581 21128 1593 21131
rect 1544 21100 1593 21128
rect 1544 21088 1550 21100
rect 1581 21097 1593 21100
rect 1627 21097 1639 21131
rect 1581 21091 1639 21097
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 2639 21131 2697 21137
rect 2639 21128 2651 21131
rect 2096 21100 2651 21128
rect 2096 21088 2102 21100
rect 2639 21097 2651 21100
rect 2685 21097 2697 21131
rect 2639 21091 2697 21097
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 2222 20992 2228 21004
rect 1443 20964 2228 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 2222 20952 2228 20964
rect 2280 20952 2286 21004
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 2590 20992 2596 21004
rect 2547 20964 2596 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 2590 20952 2596 20964
rect 2648 20952 2654 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 1464 20383 1522 20389
rect 1464 20349 1476 20383
rect 1510 20380 1522 20383
rect 1510 20352 1900 20380
rect 1510 20349 1522 20352
rect 1464 20343 1522 20349
rect 1872 20256 1900 20352
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1535 20247 1593 20253
rect 1535 20244 1547 20247
rect 1452 20216 1547 20244
rect 1452 20204 1458 20216
rect 1535 20213 1547 20216
rect 1581 20213 1593 20247
rect 1854 20244 1860 20256
rect 1815 20216 1860 20244
rect 1535 20207 1593 20213
rect 1854 20204 1860 20216
rect 1912 20204 1918 20256
rect 2590 20244 2596 20256
rect 2551 20216 2596 20244
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 2222 20000 2228 20052
rect 2280 20040 2286 20052
rect 2639 20043 2697 20049
rect 2639 20040 2651 20043
rect 2280 20012 2651 20040
rect 2280 20000 2286 20012
rect 2639 20009 2651 20012
rect 2685 20009 2697 20043
rect 2639 20003 2697 20009
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2314 19904 2320 19916
rect 1443 19876 2320 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2568 19907 2626 19913
rect 2568 19873 2580 19907
rect 2614 19904 2626 19907
rect 3326 19904 3332 19916
rect 2614 19876 3332 19904
rect 2614 19873 2626 19876
rect 2568 19867 2626 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 2314 19456 2320 19468
rect 2372 19496 2378 19508
rect 2639 19499 2697 19505
rect 2639 19496 2651 19499
rect 2372 19468 2651 19496
rect 2372 19456 2378 19468
rect 2639 19465 2651 19468
rect 2685 19465 2697 19499
rect 3326 19496 3332 19508
rect 3287 19468 3332 19496
rect 2639 19459 2697 19465
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1443 19264 2084 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2056 19168 2084 19264
rect 2130 19252 2136 19304
rect 2188 19292 2194 19304
rect 2536 19295 2594 19301
rect 2536 19292 2548 19295
rect 2188 19264 2548 19292
rect 2188 19252 2194 19264
rect 2536 19261 2548 19264
rect 2582 19292 2594 19295
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2582 19264 2973 19292
rect 2582 19261 2594 19264
rect 2536 19255 2594 19261
rect 2961 19261 2973 19264
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 3326 19184 3332 19236
rect 3384 19224 3390 19236
rect 4798 19224 4804 19236
rect 3384 19196 4804 19224
rect 3384 19184 3390 19196
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 3510 19156 3516 19168
rect 3471 19128 3516 19156
rect 3510 19116 3516 19128
rect 3568 19116 3574 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 106 18912 112 18964
rect 164 18952 170 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 164 18924 1593 18952
rect 164 18912 170 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 4203 18955 4261 18961
rect 4203 18952 4215 18955
rect 2096 18924 4215 18952
rect 2096 18912 2102 18924
rect 4203 18921 4215 18924
rect 4249 18921 4261 18955
rect 4203 18915 4261 18921
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18816 1458 18828
rect 1949 18819 2007 18825
rect 1949 18816 1961 18819
rect 1452 18788 1961 18816
rect 1452 18776 1458 18788
rect 1949 18785 1961 18788
rect 1995 18785 2007 18819
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 1949 18779 2007 18785
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 3970 18816 3976 18828
rect 3931 18788 3976 18816
rect 3970 18776 3976 18788
rect 4028 18776 4034 18828
rect 14 18640 20 18692
rect 72 18680 78 18692
rect 2685 18683 2743 18689
rect 2685 18680 2697 18683
rect 72 18652 2697 18680
rect 72 18640 78 18652
rect 2685 18649 2697 18652
rect 2731 18649 2743 18683
rect 2685 18643 2743 18649
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 4847 18411 4905 18417
rect 4847 18408 4859 18411
rect 3476 18380 4859 18408
rect 3476 18368 3482 18380
rect 4847 18377 4859 18380
rect 4893 18377 4905 18411
rect 4847 18371 4905 18377
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18204 2099 18207
rect 2869 18207 2927 18213
rect 2087 18176 2544 18204
rect 2087 18173 2099 18176
rect 2041 18167 2099 18173
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 2516 18077 2544 18176
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3326 18204 3332 18216
rect 2915 18176 3332 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 4776 18207 4834 18213
rect 4776 18173 4788 18207
rect 4822 18204 4834 18207
rect 5261 18207 5319 18213
rect 5261 18204 5273 18207
rect 4822 18176 5273 18204
rect 4822 18173 4834 18176
rect 4776 18167 4834 18173
rect 5261 18173 5273 18176
rect 5307 18204 5319 18207
rect 5994 18204 6000 18216
rect 5307 18176 6000 18204
rect 5307 18173 5319 18176
rect 5261 18167 5319 18173
rect 5994 18164 6000 18176
rect 6052 18164 6058 18216
rect 2958 18136 2964 18148
rect 2919 18108 2964 18136
rect 2958 18096 2964 18108
rect 3016 18096 3022 18148
rect 2501 18071 2559 18077
rect 2501 18037 2513 18071
rect 2547 18068 2559 18071
rect 2682 18068 2688 18080
rect 2547 18040 2688 18068
rect 2547 18037 2559 18040
rect 2501 18031 2559 18037
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 3970 18068 3976 18080
rect 3108 18040 3976 18068
rect 3108 18028 3114 18040
rect 3970 18028 3976 18040
rect 4028 18068 4034 18080
rect 4065 18071 4123 18077
rect 4065 18068 4077 18071
rect 4028 18040 4077 18068
rect 4028 18028 4034 18040
rect 4065 18037 4077 18040
rect 4111 18037 4123 18071
rect 4065 18031 4123 18037
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 5721 18071 5779 18077
rect 5721 18068 5733 18071
rect 5316 18040 5733 18068
rect 5316 18028 5322 18040
rect 5721 18037 5733 18040
rect 5767 18037 5779 18071
rect 5721 18031 5779 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 3510 17864 3516 17876
rect 3375 17836 3516 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 5767 17867 5825 17873
rect 5767 17864 5779 17867
rect 4948 17836 5779 17864
rect 4948 17824 4954 17836
rect 5767 17833 5779 17836
rect 5813 17833 5825 17867
rect 5767 17827 5825 17833
rect 2222 17728 2228 17740
rect 2183 17700 2228 17728
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 4982 17728 4988 17740
rect 4755 17700 4988 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 4982 17688 4988 17700
rect 5040 17688 5046 17740
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 5664 17731 5722 17737
rect 5664 17728 5676 17731
rect 5592 17700 5676 17728
rect 5592 17688 5598 17700
rect 5664 17697 5676 17700
rect 5710 17697 5722 17731
rect 5664 17691 5722 17697
rect 3418 17620 3424 17672
rect 3476 17660 3482 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3476 17632 4077 17660
rect 3476 17620 3482 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 5224 17632 6653 17660
rect 5224 17620 5230 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1820 17496 1961 17524
rect 1820 17484 1826 17496
rect 1949 17493 1961 17496
rect 1995 17493 2007 17527
rect 1949 17487 2007 17493
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 2777 17527 2835 17533
rect 2777 17524 2789 17527
rect 2556 17496 2789 17524
rect 2556 17484 2562 17496
rect 2777 17493 2789 17496
rect 2823 17524 2835 17527
rect 3878 17524 3884 17536
rect 2823 17496 3884 17524
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 7423 17323 7481 17329
rect 7423 17320 7435 17323
rect 2004 17292 7435 17320
rect 2004 17280 2010 17292
rect 7423 17289 7435 17292
rect 7469 17289 7481 17323
rect 7423 17283 7481 17289
rect 2777 17255 2835 17261
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 3234 17252 3240 17264
rect 2823 17224 3240 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 2792 17116 2820 17215
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 5534 17252 5540 17264
rect 4126 17224 5540 17252
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17184 3387 17187
rect 3510 17184 3516 17196
rect 3375 17156 3516 17184
rect 3375 17153 3387 17156
rect 3329 17147 3387 17153
rect 3510 17144 3516 17156
rect 3568 17144 3574 17196
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 4126 17184 4154 17224
rect 5534 17212 5540 17224
rect 5592 17252 5598 17264
rect 6181 17255 6239 17261
rect 6181 17252 6193 17255
rect 5592 17224 6193 17252
rect 5592 17212 5598 17224
rect 6181 17221 6193 17224
rect 6227 17221 6239 17255
rect 6181 17215 6239 17221
rect 5258 17184 5264 17196
rect 3660 17156 4154 17184
rect 5219 17156 5264 17184
rect 3660 17144 3666 17156
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 2363 17088 2820 17116
rect 7352 17119 7410 17125
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 7352 17085 7364 17119
rect 7398 17116 7410 17119
rect 7558 17116 7564 17128
rect 7398 17088 7564 17116
rect 7398 17085 7410 17088
rect 7352 17079 7410 17085
rect 7558 17076 7564 17088
rect 7616 17116 7622 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7616 17088 7757 17116
rect 7616 17076 7622 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 3145 17051 3203 17057
rect 3145 17017 3157 17051
rect 3191 17048 3203 17051
rect 3418 17048 3424 17060
rect 3191 17020 3424 17048
rect 3191 17017 3203 17020
rect 3145 17011 3203 17017
rect 3418 17008 3424 17020
rect 3476 17008 3482 17060
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 5905 17051 5963 17057
rect 5408 17020 5453 17048
rect 5408 17008 5414 17020
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 5994 17048 6000 17060
rect 5951 17020 6000 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 5994 17008 6000 17020
rect 6052 17008 6058 17060
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 2924 16952 4353 16980
rect 2924 16940 2930 16952
rect 4341 16949 4353 16952
rect 4387 16980 4399 16983
rect 4982 16980 4988 16992
rect 4387 16952 4988 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5077 16983 5135 16989
rect 5077 16949 5089 16983
rect 5123 16980 5135 16983
rect 5368 16980 5396 17008
rect 5123 16952 5396 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 8110 16940 8116 16992
rect 8168 16980 8174 16992
rect 8297 16983 8355 16989
rect 8297 16980 8309 16983
rect 8168 16952 8309 16980
rect 8168 16940 8174 16952
rect 8297 16949 8309 16952
rect 8343 16949 8355 16983
rect 8297 16943 8355 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2314 16776 2320 16788
rect 2227 16748 2320 16776
rect 2314 16736 2320 16748
rect 2372 16776 2378 16788
rect 2866 16776 2872 16788
rect 2372 16748 2872 16776
rect 2372 16736 2378 16748
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 5258 16776 5264 16788
rect 5219 16748 5264 16776
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 2593 16711 2651 16717
rect 2593 16677 2605 16711
rect 2639 16708 2651 16711
rect 2958 16708 2964 16720
rect 2639 16680 2964 16708
rect 2639 16677 2651 16680
rect 2593 16671 2651 16677
rect 2958 16668 2964 16680
rect 3016 16668 3022 16720
rect 4430 16708 4436 16720
rect 3436 16680 4436 16708
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1578 16640 1584 16652
rect 1510 16612 1584 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2222 16572 2228 16584
rect 1995 16544 2228 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2498 16572 2504 16584
rect 2459 16544 2504 16572
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 2130 16464 2136 16516
rect 2188 16504 2194 16516
rect 2792 16504 2820 16535
rect 3436 16513 3464 16680
rect 4430 16668 4436 16680
rect 4488 16668 4494 16720
rect 5350 16708 5356 16720
rect 5311 16680 5356 16708
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 8018 16668 8024 16720
rect 8076 16708 8082 16720
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 8076 16680 8125 16708
rect 8076 16668 8082 16680
rect 8113 16677 8125 16680
rect 8159 16677 8171 16711
rect 8113 16671 8171 16677
rect 3970 16640 3976 16652
rect 3931 16612 3976 16640
rect 3970 16600 3976 16612
rect 4028 16600 4034 16652
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16640 6055 16643
rect 6270 16640 6276 16652
rect 6043 16612 6276 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6952 16643 7010 16649
rect 6952 16640 6964 16643
rect 6604 16612 6964 16640
rect 6604 16600 6610 16612
rect 6952 16609 6964 16612
rect 6998 16609 7010 16643
rect 6952 16603 7010 16609
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16572 8079 16575
rect 8110 16572 8116 16584
rect 8067 16544 8116 16572
rect 8067 16541 8079 16544
rect 8021 16535 8079 16541
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 8297 16575 8355 16581
rect 8297 16541 8309 16575
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 3421 16507 3479 16513
rect 3421 16504 3433 16507
rect 2188 16476 3433 16504
rect 2188 16464 2194 16476
rect 3421 16473 3433 16476
rect 3467 16473 3479 16507
rect 3421 16467 3479 16473
rect 3694 16464 3700 16516
rect 3752 16504 3758 16516
rect 7055 16507 7113 16513
rect 7055 16504 7067 16507
rect 3752 16476 7067 16504
rect 3752 16464 3758 16476
rect 7055 16473 7067 16476
rect 7101 16473 7113 16507
rect 7055 16467 7113 16473
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 8312 16504 8340 16535
rect 7616 16476 8340 16504
rect 7616 16464 7622 16476
rect 1535 16439 1593 16445
rect 1535 16405 1547 16439
rect 1581 16436 1593 16439
rect 2406 16436 2412 16448
rect 1581 16408 2412 16436
rect 1581 16405 1593 16408
rect 1535 16399 1593 16405
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 4203 16439 4261 16445
rect 4203 16436 4215 16439
rect 2556 16408 4215 16436
rect 2556 16396 2562 16408
rect 4203 16405 4215 16408
rect 4249 16405 4261 16439
rect 4203 16399 4261 16405
rect 7469 16439 7527 16445
rect 7469 16405 7481 16439
rect 7515 16436 7527 16439
rect 7926 16436 7932 16448
rect 7515 16408 7932 16436
rect 7515 16405 7527 16408
rect 7469 16399 7527 16405
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 8570 16396 8576 16448
rect 8628 16436 8634 16448
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8628 16408 8953 16436
rect 8628 16396 8634 16408
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 3016 16204 3065 16232
rect 3016 16192 3022 16204
rect 3053 16201 3065 16204
rect 3099 16201 3111 16235
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 3053 16195 3111 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 8168 16204 9597 16232
rect 8168 16192 8174 16204
rect 9585 16201 9597 16204
rect 9631 16201 9643 16235
rect 9585 16195 9643 16201
rect 3970 16164 3976 16176
rect 2583 16136 3976 16164
rect 106 16056 112 16108
rect 164 16096 170 16108
rect 2583 16096 2611 16136
rect 3970 16124 3976 16136
rect 4028 16164 4034 16176
rect 4617 16167 4675 16173
rect 4617 16164 4629 16167
rect 4028 16136 4629 16164
rect 4028 16124 4034 16136
rect 4617 16133 4629 16136
rect 4663 16133 4675 16167
rect 4617 16127 4675 16133
rect 164 16068 2611 16096
rect 2777 16099 2835 16105
rect 164 16056 170 16068
rect 2777 16065 2789 16099
rect 2823 16096 2835 16099
rect 3510 16096 3516 16108
rect 2823 16068 3516 16096
rect 2823 16065 2835 16068
rect 2777 16059 2835 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 3694 16096 3700 16108
rect 3655 16068 3700 16096
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16096 5963 16099
rect 5994 16096 6000 16108
rect 5951 16068 6000 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 8570 16028 8576 16040
rect 8435 16000 8576 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 2130 15960 2136 15972
rect 2091 15932 2136 15960
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 2225 15963 2283 15969
rect 2225 15929 2237 15963
rect 2271 15960 2283 15963
rect 2314 15960 2320 15972
rect 2271 15932 2320 15960
rect 2271 15929 2283 15932
rect 2225 15923 2283 15929
rect 2314 15920 2320 15932
rect 2372 15920 2378 15972
rect 3510 15960 3516 15972
rect 3471 15932 3516 15960
rect 3510 15920 3516 15932
rect 3568 15960 3574 15972
rect 3766 15963 3824 15969
rect 3766 15960 3778 15963
rect 3568 15932 3778 15960
rect 3568 15920 3574 15932
rect 3766 15929 3778 15932
rect 3812 15929 3824 15963
rect 4338 15960 4344 15972
rect 4299 15932 4344 15960
rect 3766 15923 3824 15929
rect 4338 15920 4344 15932
rect 4396 15960 4402 15972
rect 5258 15960 5264 15972
rect 4396 15932 5264 15960
rect 4396 15920 4402 15932
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 5353 15963 5411 15969
rect 5353 15929 5365 15963
rect 5399 15960 5411 15963
rect 6917 15963 6975 15969
rect 5399 15932 6316 15960
rect 5399 15929 5411 15932
rect 5353 15923 5411 15929
rect 5077 15895 5135 15901
rect 5077 15861 5089 15895
rect 5123 15892 5135 15895
rect 5368 15892 5396 15923
rect 6288 15904 6316 15932
rect 6917 15929 6929 15963
rect 6963 15929 6975 15963
rect 6917 15923 6975 15929
rect 7009 15963 7067 15969
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 7834 15960 7840 15972
rect 7055 15932 7840 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 6270 15892 6276 15904
rect 5123 15864 5396 15892
rect 6231 15864 6276 15892
rect 5123 15861 5135 15864
rect 5077 15855 5135 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 6932 15892 6960 15923
rect 7834 15920 7840 15932
rect 7892 15920 7898 15972
rect 8710 15963 8768 15969
rect 8710 15929 8722 15963
rect 8756 15929 8768 15963
rect 8710 15923 8768 15929
rect 6880 15864 6960 15892
rect 7929 15895 7987 15901
rect 6880 15852 6886 15864
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 8018 15892 8024 15904
rect 7975 15864 8024 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 8297 15895 8355 15901
rect 8297 15861 8309 15895
rect 8343 15892 8355 15895
rect 8386 15892 8392 15904
rect 8343 15864 8392 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 8386 15852 8392 15864
rect 8444 15892 8450 15904
rect 8725 15892 8753 15923
rect 9306 15892 9312 15904
rect 8444 15864 8753 15892
rect 9267 15864 9312 15892
rect 8444 15852 8450 15864
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2556 15660 3249 15688
rect 2556 15648 2562 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3694 15688 3700 15700
rect 3655 15660 3700 15688
rect 3237 15651 3295 15657
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5813 15691 5871 15697
rect 5813 15688 5825 15691
rect 5316 15660 5825 15688
rect 5316 15648 5322 15660
rect 5813 15657 5825 15660
rect 5859 15657 5871 15691
rect 5813 15651 5871 15657
rect 1670 15620 1676 15632
rect 1631 15592 1676 15620
rect 1670 15580 1676 15592
rect 1728 15580 1734 15632
rect 3510 15580 3516 15632
rect 3568 15620 3574 15632
rect 4801 15623 4859 15629
rect 4801 15620 4813 15623
rect 3568 15592 4813 15620
rect 3568 15580 3574 15592
rect 4801 15589 4813 15592
rect 4847 15589 4859 15623
rect 6638 15620 6644 15632
rect 6599 15592 6644 15620
rect 4801 15583 4859 15589
rect 6638 15580 6644 15592
rect 6696 15580 6702 15632
rect 8018 15620 8024 15632
rect 7979 15592 8024 15620
rect 8018 15580 8024 15592
rect 8076 15580 8082 15632
rect 2406 15512 2412 15564
rect 2464 15552 2470 15564
rect 5442 15552 5448 15564
rect 2464 15524 4154 15552
rect 5403 15524 5448 15552
rect 2464 15512 2470 15524
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 2774 15484 2780 15496
rect 1627 15456 2780 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 4126 15484 4154 15524
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 7926 15552 7932 15564
rect 7839 15524 7932 15552
rect 7926 15512 7932 15524
rect 7984 15552 7990 15564
rect 8665 15555 8723 15561
rect 8665 15552 8677 15555
rect 7984 15524 8677 15552
rect 7984 15512 7990 15524
rect 8665 15521 8677 15524
rect 8711 15552 8723 15555
rect 9306 15552 9312 15564
rect 8711 15524 9312 15552
rect 8711 15521 8723 15524
rect 8665 15515 8723 15521
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 6273 15487 6331 15493
rect 6273 15484 6285 15487
rect 4126 15456 6285 15484
rect 6273 15453 6285 15456
rect 6319 15484 6331 15487
rect 6549 15487 6607 15493
rect 6549 15484 6561 15487
rect 6319 15456 6561 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 6549 15453 6561 15456
rect 6595 15453 6607 15487
rect 6822 15484 6828 15496
rect 6783 15456 6828 15484
rect 6549 15447 6607 15453
rect 6822 15444 6828 15456
rect 6880 15484 6886 15496
rect 7469 15487 7527 15493
rect 7469 15484 7481 15487
rect 6880 15456 7481 15484
rect 6880 15444 6886 15456
rect 7469 15453 7481 15456
rect 7515 15453 7527 15487
rect 7469 15447 7527 15453
rect 1854 15376 1860 15428
rect 1912 15416 1918 15428
rect 2130 15416 2136 15428
rect 1912 15388 2136 15416
rect 1912 15376 1918 15388
rect 2130 15376 2136 15388
rect 2188 15376 2194 15428
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15348 2651 15351
rect 2682 15348 2688 15360
rect 2639 15320 2688 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 2866 15348 2872 15360
rect 2827 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2832 15116 2881 15144
rect 2832 15104 2838 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 3513 15147 3571 15153
rect 3513 15113 3525 15147
rect 3559 15144 3571 15147
rect 3786 15144 3792 15156
rect 3559 15116 3792 15144
rect 3559 15113 3571 15116
rect 3513 15107 3571 15113
rect 2130 15036 2136 15088
rect 2188 15076 2194 15088
rect 2501 15079 2559 15085
rect 2501 15076 2513 15079
rect 2188 15048 2513 15076
rect 2188 15036 2194 15048
rect 2501 15045 2513 15048
rect 2547 15045 2559 15079
rect 2884 15076 2912 15107
rect 3786 15104 3792 15116
rect 3844 15144 3850 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 3844 15116 4905 15144
rect 3844 15104 3850 15116
rect 4893 15113 4905 15116
rect 4939 15144 4951 15147
rect 5442 15144 5448 15156
rect 4939 15116 5448 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5442 15104 5448 15116
rect 5500 15144 5506 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 5500 15116 9597 15144
rect 5500 15104 5506 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 5166 15076 5172 15088
rect 2884 15048 5172 15076
rect 2501 15039 2559 15045
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 5813 15079 5871 15085
rect 5813 15045 5825 15079
rect 5859 15076 5871 15079
rect 6822 15076 6828 15088
rect 5859 15048 6828 15076
rect 5859 15045 5871 15048
rect 5813 15039 5871 15045
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2314 15008 2320 15020
rect 1995 14980 2320 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2314 14968 2320 14980
rect 2372 15008 2378 15020
rect 2866 15008 2872 15020
rect 2372 14980 2872 15008
rect 2372 14968 2378 14980
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 4338 15008 4344 15020
rect 4299 14980 4344 15008
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6638 15008 6644 15020
rect 6595 14980 6644 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 6638 14968 6644 14980
rect 6696 15008 6702 15020
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 6696 14980 7113 15008
rect 6696 14968 6702 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 7190 14940 7196 14952
rect 7151 14912 7196 14940
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14940 8263 14943
rect 8662 14940 8668 14952
rect 8251 14912 8668 14940
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 2041 14875 2099 14881
rect 2041 14841 2053 14875
rect 2087 14872 2099 14875
rect 2682 14872 2688 14884
rect 2087 14844 2688 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3694 14872 3700 14884
rect 3655 14844 3700 14872
rect 3694 14832 3700 14844
rect 3752 14832 3758 14884
rect 3786 14832 3792 14884
rect 3844 14872 3850 14884
rect 5258 14872 5264 14884
rect 3844 14844 3889 14872
rect 5219 14844 5264 14872
rect 3844 14832 3850 14844
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 7208 14872 7236 14900
rect 5408 14844 7236 14872
rect 8986 14875 9044 14881
rect 5408 14832 5414 14844
rect 8986 14841 8998 14875
rect 9032 14841 9044 14875
rect 8986 14835 9044 14841
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 8444 14776 8493 14804
rect 8444 14764 8450 14776
rect 8481 14773 8493 14776
rect 8527 14804 8539 14807
rect 9001 14804 9029 14835
rect 9858 14804 9864 14816
rect 8527 14776 9864 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4982 14600 4988 14612
rect 4943 14572 4988 14600
rect 4433 14563 4491 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5350 14600 5356 14612
rect 5311 14572 5356 14600
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 6454 14600 6460 14612
rect 6190 14572 6460 14600
rect 1762 14532 1768 14544
rect 1723 14504 1768 14532
rect 1762 14492 1768 14504
rect 1820 14492 1826 14544
rect 2314 14532 2320 14544
rect 2275 14504 2320 14532
rect 2314 14492 2320 14504
rect 2372 14492 2378 14544
rect 6190 14541 6218 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7190 14600 7196 14612
rect 7103 14572 7196 14600
rect 7190 14560 7196 14572
rect 7248 14600 7254 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 7248 14572 10609 14600
rect 7248 14560 7254 14572
rect 10597 14569 10609 14572
rect 10643 14569 10655 14603
rect 10597 14563 10655 14569
rect 6175 14535 6233 14541
rect 6175 14501 6187 14535
rect 6221 14501 6233 14535
rect 6175 14495 6233 14501
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 8199 14535 8257 14541
rect 6328 14504 7880 14532
rect 6328 14492 6334 14504
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 2740 14436 6745 14464
rect 2740 14424 2746 14436
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 7852 14464 7880 14504
rect 8199 14501 8211 14535
rect 8245 14532 8257 14535
rect 8386 14532 8392 14544
rect 8245 14504 8392 14532
rect 8245 14501 8257 14504
rect 8199 14495 8257 14501
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 9998 14535 10056 14541
rect 9998 14532 10010 14535
rect 9916 14504 10010 14532
rect 9916 14492 9922 14504
rect 9998 14501 10010 14504
rect 10044 14501 10056 14535
rect 9998 14495 10056 14501
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 7852 14436 8769 14464
rect 6733 14427 6791 14433
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 1670 14396 1676 14408
rect 1583 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14396 1734 14408
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 1728 14368 2973 14396
rect 1728 14356 1734 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 2961 14359 3019 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5258 14356 5264 14408
rect 5316 14356 5322 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5592 14368 5825 14396
rect 5592 14356 5598 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 7837 14359 7895 14365
rect 5276 14328 5304 14356
rect 5629 14331 5687 14337
rect 5629 14328 5641 14331
rect 4126 14300 5641 14328
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 2593 14263 2651 14269
rect 2593 14260 2605 14263
rect 2556 14232 2605 14260
rect 2556 14220 2562 14232
rect 2593 14229 2605 14232
rect 2639 14229 2651 14263
rect 3694 14260 3700 14272
rect 3655 14232 3700 14260
rect 2593 14223 2651 14229
rect 3694 14220 3700 14232
rect 3752 14220 3758 14272
rect 3970 14220 3976 14272
rect 4028 14260 4034 14272
rect 4126 14260 4154 14300
rect 5629 14297 5641 14300
rect 5675 14297 5687 14331
rect 5629 14291 5687 14297
rect 4028 14232 4154 14260
rect 7745 14263 7803 14269
rect 4028 14220 4034 14232
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 7852 14260 7880 14359
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 8478 14260 8484 14272
rect 7791 14232 8484 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 1762 14056 1768 14068
rect 1719 14028 1768 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 6512 14028 7849 14056
rect 6512 14016 6518 14028
rect 7837 14025 7849 14028
rect 7883 14056 7895 14059
rect 8386 14056 8392 14068
rect 7883 14028 8392 14056
rect 7883 14025 7895 14028
rect 7837 14019 7895 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 9732 14028 11437 14056
rect 9732 14016 9738 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 11425 14019 11483 14025
rect 9766 13988 9772 14000
rect 9646 13960 9772 13988
rect 2314 13880 2320 13932
rect 2372 13920 2378 13932
rect 2409 13923 2467 13929
rect 2409 13920 2421 13923
rect 2372 13892 2421 13920
rect 2372 13880 2378 13892
rect 2409 13889 2421 13892
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 9646 13920 9674 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 9858 13948 9864 14000
rect 9916 13988 9922 14000
rect 9916 13960 9961 13988
rect 9916 13948 9922 13960
rect 6319 13892 9674 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 3467 13824 4261 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4249 13821 4261 13824
rect 4295 13852 4307 13855
rect 4295 13824 5764 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 2133 13787 2191 13793
rect 2133 13753 2145 13787
rect 2179 13753 2191 13787
rect 2133 13747 2191 13753
rect 2148 13716 2176 13747
rect 2222 13744 2228 13796
rect 2280 13784 2286 13796
rect 3789 13787 3847 13793
rect 2280 13756 2325 13784
rect 2280 13744 2286 13756
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 4157 13787 4215 13793
rect 4157 13784 4169 13787
rect 3835 13756 4169 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 4157 13753 4169 13756
rect 4203 13784 4215 13787
rect 4338 13784 4344 13796
rect 4203 13756 4344 13784
rect 4203 13753 4215 13756
rect 4157 13747 4215 13753
rect 4338 13744 4344 13756
rect 4396 13784 4402 13796
rect 4611 13787 4669 13793
rect 4611 13784 4623 13787
rect 4396 13756 4623 13784
rect 4396 13744 4402 13756
rect 4611 13753 4623 13756
rect 4657 13784 4669 13787
rect 5736 13784 5764 13824
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7392 13861 7420 13892
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6696 13824 6837 13852
rect 6696 13812 6702 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8444 13824 8493 13852
rect 8444 13812 8450 13824
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 9030 13852 9036 13864
rect 8991 13824 9036 13852
rect 8481 13815 8539 13821
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 9309 13855 9367 13861
rect 9309 13821 9321 13855
rect 9355 13852 9367 13855
rect 10321 13855 10379 13861
rect 9355 13824 9389 13852
rect 9355 13821 9367 13824
rect 9309 13815 9367 13821
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 10367 13824 10425 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10413 13821 10425 13824
rect 10459 13852 10471 13855
rect 10870 13852 10876 13864
rect 10459 13824 10732 13852
rect 10831 13824 10876 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 4657 13756 5672 13784
rect 5736 13756 8708 13784
rect 4657 13753 4669 13756
rect 4611 13747 4669 13753
rect 2498 13716 2504 13728
rect 2148 13688 2504 13716
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 5644 13716 5672 13756
rect 5810 13716 5816 13728
rect 5644 13688 5816 13716
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 6638 13716 6644 13728
rect 6599 13688 6644 13716
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 8386 13716 8392 13728
rect 8347 13688 8392 13716
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 8570 13716 8576 13728
rect 8531 13688 8576 13716
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 8680 13716 8708 13756
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9324 13784 9352 13815
rect 10704 13796 10732 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 9180 13756 9352 13784
rect 9180 13744 9186 13756
rect 10686 13744 10692 13796
rect 10744 13744 10750 13796
rect 10505 13719 10563 13725
rect 10505 13716 10517 13719
rect 8680 13688 10517 13716
rect 10505 13685 10517 13688
rect 10551 13685 10563 13719
rect 10505 13679 10563 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1535 13515 1593 13521
rect 1535 13481 1547 13515
rect 1581 13512 1593 13515
rect 1670 13512 1676 13524
rect 1581 13484 1676 13512
rect 1581 13481 1593 13484
rect 1535 13475 1593 13481
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 5592 13484 7665 13512
rect 5592 13472 5598 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10321 13515 10379 13521
rect 10321 13512 10333 13515
rect 9824 13484 10333 13512
rect 9824 13472 9830 13484
rect 10321 13481 10333 13484
rect 10367 13512 10379 13515
rect 10870 13512 10876 13524
rect 10367 13484 10876 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 3326 13404 3332 13456
rect 3384 13444 3390 13456
rect 3786 13444 3792 13456
rect 3384 13416 3792 13444
rect 3384 13404 3390 13416
rect 3786 13404 3792 13416
rect 3844 13444 3850 13456
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 3844 13416 4261 13444
rect 3844 13404 3850 13416
rect 4249 13413 4261 13416
rect 4295 13444 4307 13447
rect 5166 13444 5172 13456
rect 4295 13416 5172 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 5166 13404 5172 13416
rect 5224 13404 5230 13456
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 6175 13447 6233 13453
rect 6175 13444 6187 13447
rect 5868 13416 6187 13444
rect 5868 13404 5874 13416
rect 6175 13413 6187 13416
rect 6221 13444 6233 13447
rect 6546 13444 6552 13456
rect 6221 13416 6552 13444
rect 6221 13413 6233 13416
rect 6175 13407 6233 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 9033 13447 9091 13453
rect 9033 13413 9045 13447
rect 9079 13444 9091 13447
rect 9306 13444 9312 13456
rect 9079 13416 9312 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 9306 13404 9312 13416
rect 9364 13444 9370 13456
rect 10686 13444 10692 13456
rect 9364 13416 10692 13444
rect 9364 13404 9370 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 1464 13379 1522 13385
rect 1464 13345 1476 13379
rect 1510 13376 1522 13379
rect 1578 13376 1584 13388
rect 1510 13348 1584 13376
rect 1510 13345 1522 13348
rect 1464 13339 1522 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2774 13376 2780 13388
rect 2735 13348 2780 13376
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 2406 13308 2412 13320
rect 2367 13280 2412 13308
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13308 4215 13311
rect 4246 13308 4252 13320
rect 4203 13280 4252 13308
rect 4203 13277 4215 13280
rect 4157 13271 4215 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 4430 13308 4436 13320
rect 4391 13280 4436 13308
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 5994 13308 6000 13320
rect 5859 13280 6000 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 7576 13308 7604 13339
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7708 13348 8033 13376
rect 7708 13336 7714 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9858 13376 9864 13388
rect 9723 13348 9864 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9858 13336 9864 13348
rect 9916 13376 9922 13388
rect 11241 13379 11299 13385
rect 11241 13376 11253 13379
rect 9916 13348 11253 13376
rect 9916 13336 9922 13348
rect 11241 13345 11253 13348
rect 11287 13376 11299 13379
rect 11882 13376 11888 13388
rect 11287 13348 11888 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 6696 13280 7972 13308
rect 6696 13268 6702 13280
rect 7944 13252 7972 13280
rect 9416 13280 10057 13308
rect 2133 13243 2191 13249
rect 2133 13209 2145 13243
rect 2179 13240 2191 13243
rect 2222 13240 2228 13252
rect 2179 13212 2228 13240
rect 2179 13209 2191 13212
rect 2133 13203 2191 13209
rect 2222 13200 2228 13212
rect 2280 13240 2286 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 2280 13212 6745 13240
rect 2280 13200 2286 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6733 13203 6791 13209
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 7984 13212 8677 13240
rect 7984 13200 7990 13212
rect 8665 13209 8677 13212
rect 8711 13240 8723 13243
rect 9122 13240 9128 13252
rect 8711 13212 9128 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9416 13184 9444 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 12250 13308 12256 13320
rect 12211 13280 12256 13308
rect 10045 13271 10103 13277
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 11425 13243 11483 13249
rect 11425 13240 11437 13243
rect 9732 13212 11437 13240
rect 9732 13200 9738 13212
rect 11425 13209 11437 13212
rect 11471 13209 11483 13243
rect 11425 13203 11483 13209
rect 3881 13175 3939 13181
rect 3881 13141 3893 13175
rect 3927 13172 3939 13175
rect 4062 13172 4068 13184
rect 3927 13144 4068 13172
rect 3927 13141 3939 13144
rect 3881 13135 3939 13141
rect 4062 13132 4068 13144
rect 4120 13172 4126 13184
rect 6914 13172 6920 13184
rect 4120 13144 6920 13172
rect 4120 13132 4126 13144
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 9398 13172 9404 13184
rect 7064 13144 7109 13172
rect 9359 13144 9404 13172
rect 7064 13132 7070 13144
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 9815 13175 9873 13181
rect 9815 13172 9827 13175
rect 9640 13144 9827 13172
rect 9640 13132 9646 13144
rect 9815 13141 9827 13144
rect 9861 13141 9873 13175
rect 9815 13135 9873 13141
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 10134 13172 10140 13184
rect 9999 13144 10140 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2406 12968 2412 12980
rect 2271 12940 2412 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 3786 12968 3792 12980
rect 3747 12940 3792 12968
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9858 12968 9864 12980
rect 9819 12940 9864 12968
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 5077 12903 5135 12909
rect 5077 12869 5089 12903
rect 5123 12900 5135 12903
rect 5123 12872 8616 12900
rect 5123 12869 5135 12872
rect 5077 12863 5135 12869
rect 1486 12792 1492 12844
rect 1544 12832 1550 12844
rect 2498 12832 2504 12844
rect 1544 12804 2504 12832
rect 1544 12792 1550 12804
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2685 12835 2743 12841
rect 2685 12832 2697 12835
rect 2648 12804 2697 12832
rect 2648 12792 2654 12804
rect 2685 12801 2697 12804
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 3948 12767 4006 12773
rect 3948 12733 3960 12767
rect 3994 12764 4006 12767
rect 4154 12764 4160 12776
rect 3994 12736 4160 12764
rect 3994 12733 4006 12736
rect 3948 12727 4006 12733
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 5184 12773 5212 12872
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 5994 12832 6000 12844
rect 5951 12804 6000 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6052 12804 6561 12832
rect 6052 12792 6058 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 7650 12832 7656 12844
rect 6549 12795 6607 12801
rect 6656 12804 7656 12832
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4212 12736 4353 12764
rect 4212 12724 4218 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5721 12767 5779 12773
rect 5721 12764 5733 12767
rect 5316 12736 5733 12764
rect 5316 12724 5322 12736
rect 5721 12733 5733 12736
rect 5767 12764 5779 12767
rect 6656 12764 6684 12804
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7006 12764 7012 12776
rect 5767 12736 6684 12764
rect 6967 12736 7012 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8444 12736 8493 12764
rect 8444 12724 8450 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8588 12764 8616 12872
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 9088 12804 9413 12832
rect 9088 12792 9094 12804
rect 9401 12801 9413 12804
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9306 12764 9312 12776
rect 8588 12736 9312 12764
rect 8481 12727 8539 12733
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12665 2467 12699
rect 2409 12659 2467 12665
rect 2424 12628 2452 12659
rect 2498 12656 2504 12708
rect 2556 12696 2562 12708
rect 2556 12668 2601 12696
rect 2556 12656 2562 12668
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 6825 12699 6883 12705
rect 6825 12696 6837 12699
rect 4304 12668 6837 12696
rect 4304 12656 4310 12668
rect 6825 12665 6837 12668
rect 6871 12665 6883 12699
rect 6825 12659 6883 12665
rect 3418 12628 3424 12640
rect 2424 12600 3424 12628
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 4019 12631 4077 12637
rect 4019 12628 4031 12631
rect 3844 12600 4031 12628
rect 3844 12588 3850 12600
rect 4019 12597 4031 12600
rect 4065 12597 4077 12631
rect 4019 12591 4077 12597
rect 6273 12631 6331 12637
rect 6273 12597 6285 12631
rect 6319 12628 6331 12631
rect 6546 12628 6552 12640
rect 6319 12600 6552 12628
rect 6319 12597 6331 12600
rect 6273 12591 6331 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12628 8447 12631
rect 8496 12628 8524 12727
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9416 12764 9444 12795
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9548 12804 9597 12832
rect 9548 12792 9554 12804
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 9692 12804 11100 12832
rect 9692 12776 9720 12804
rect 11072 12776 11100 12804
rect 9674 12764 9680 12776
rect 9416 12736 9680 12764
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 10597 12767 10655 12773
rect 10597 12764 10609 12767
rect 10367 12736 10609 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 10597 12733 10609 12736
rect 10643 12733 10655 12767
rect 11054 12764 11060 12776
rect 11015 12736 11060 12764
rect 10597 12727 10655 12733
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 8720 12668 10364 12696
rect 8720 12656 8726 12668
rect 9766 12628 9772 12640
rect 8435 12600 9772 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 10336 12628 10364 12668
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 10336 12600 10517 12628
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10612 12628 10640 12727
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12733 11299 12767
rect 11241 12727 11299 12733
rect 12504 12767 12562 12773
rect 12504 12733 12516 12767
rect 12550 12764 12562 12767
rect 12894 12764 12900 12776
rect 12550 12736 12900 12764
rect 12550 12733 12562 12736
rect 12504 12727 12562 12733
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11256 12696 11284 12727
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 11882 12696 11888 12708
rect 10744 12668 11284 12696
rect 11795 12668 11888 12696
rect 10744 12656 10750 12668
rect 11882 12656 11888 12668
rect 11940 12696 11946 12708
rect 18598 12696 18604 12708
rect 11940 12668 18604 12696
rect 11940 12656 11946 12668
rect 18598 12656 18604 12668
rect 18656 12656 18662 12708
rect 11146 12628 11152 12640
rect 10612 12600 11152 12628
rect 10505 12591 10563 12597
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 12575 12631 12633 12637
rect 12575 12597 12587 12631
rect 12621 12628 12633 12631
rect 12710 12628 12716 12640
rect 12621 12600 12716 12628
rect 12621 12597 12633 12600
rect 12575 12591 12633 12597
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1946 12424 1952 12436
rect 1907 12396 1952 12424
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 6641 12427 6699 12433
rect 6641 12424 6653 12427
rect 6503 12396 6653 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6641 12393 6653 12396
rect 6687 12424 6699 12427
rect 6822 12424 6828 12436
rect 6687 12396 6828 12424
rect 6687 12393 6699 12396
rect 6641 12387 6699 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 11054 12424 11060 12436
rect 7156 12396 10364 12424
rect 11015 12396 11060 12424
rect 7156 12384 7162 12396
rect 2317 12359 2375 12365
rect 2317 12325 2329 12359
rect 2363 12356 2375 12359
rect 2593 12359 2651 12365
rect 2593 12356 2605 12359
rect 2363 12328 2605 12356
rect 2363 12325 2375 12328
rect 2317 12319 2375 12325
rect 2593 12325 2605 12328
rect 2639 12356 2651 12359
rect 2774 12356 2780 12368
rect 2639 12328 2780 12356
rect 2639 12325 2651 12328
rect 2593 12319 2651 12325
rect 2774 12316 2780 12328
rect 2832 12316 2838 12368
rect 4246 12356 4252 12368
rect 4207 12328 4252 12356
rect 4246 12316 4252 12328
rect 4304 12316 4310 12368
rect 4798 12356 4804 12368
rect 4759 12328 4804 12356
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 5629 12359 5687 12365
rect 5629 12325 5641 12359
rect 5675 12356 5687 12359
rect 5994 12356 6000 12368
rect 5675 12328 6000 12356
rect 5675 12325 5687 12328
rect 5629 12319 5687 12325
rect 5994 12316 6000 12328
rect 6052 12356 6058 12368
rect 6914 12356 6920 12368
rect 6052 12328 6920 12356
rect 6052 12316 6058 12328
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 8021 12359 8079 12365
rect 8021 12325 8033 12359
rect 8067 12356 8079 12359
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 8067 12328 8401 12356
rect 8067 12325 8079 12328
rect 8021 12319 8079 12325
rect 8389 12325 8401 12328
rect 8435 12356 8447 12359
rect 9674 12356 9680 12368
rect 8435 12328 9680 12356
rect 8435 12325 8447 12328
rect 8389 12319 8447 12325
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 1464 12291 1522 12297
rect 1464 12257 1476 12291
rect 1510 12288 1522 12291
rect 1578 12288 1584 12300
rect 1510 12260 1584 12288
rect 1510 12257 1522 12260
rect 1464 12251 1522 12257
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 6638 12288 6644 12300
rect 6599 12260 6644 12288
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6788 12260 7021 12288
rect 6788 12248 6794 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7009 12251 7067 12257
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 10336 12297 10364 12396
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 11204 12396 13001 12424
rect 11204 12384 11210 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 10502 12316 10508 12368
rect 10560 12356 10566 12368
rect 11164 12356 11192 12384
rect 10560 12328 11192 12356
rect 10560 12316 10566 12328
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 8168 12260 8493 12288
rect 8168 12248 8174 12260
rect 8481 12257 8493 12260
rect 8527 12288 8539 12291
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 8527 12260 9229 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 9217 12257 9229 12260
rect 9263 12257 9275 12291
rect 9217 12251 9275 12257
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 11698 12288 11704 12300
rect 10367 12260 11468 12288
rect 11659 12260 11704 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2648 12192 2789 12220
rect 2648 12180 2654 12192
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 2924 12192 3924 12220
rect 2924 12180 2930 12192
rect 1762 12112 1768 12164
rect 1820 12152 1826 12164
rect 3421 12155 3479 12161
rect 3421 12152 3433 12155
rect 1820 12124 3433 12152
rect 1820 12112 1826 12124
rect 3421 12121 3433 12124
rect 3467 12152 3479 12155
rect 3786 12152 3792 12164
rect 3467 12124 3792 12152
rect 3467 12121 3479 12124
rect 3421 12115 3479 12121
rect 3786 12112 3792 12124
rect 3844 12112 3850 12164
rect 3896 12152 3924 12192
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 4212 12192 4257 12220
rect 4448 12192 9689 12220
rect 4212 12180 4218 12192
rect 4448 12152 4476 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 9916 12192 11253 12220
rect 9916 12180 9922 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11440 12220 11468 12260
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 11848 12260 12817 12288
rect 11848 12248 11854 12260
rect 12805 12257 12817 12260
rect 12851 12288 12863 12291
rect 13170 12288 13176 12300
rect 12851 12260 13176 12288
rect 12851 12257 12863 12260
rect 12805 12251 12863 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 13872 12260 13917 12288
rect 13872 12248 13878 12260
rect 12342 12220 12348 12232
rect 11440 12192 12348 12220
rect 11241 12183 11299 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 12986 12220 12992 12232
rect 12575 12192 12992 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13955 12223 14013 12229
rect 13955 12220 13967 12223
rect 13504 12192 13967 12220
rect 13504 12180 13510 12192
rect 13955 12189 13967 12192
rect 14001 12189 14013 12223
rect 13955 12183 14013 12189
rect 8018 12152 8024 12164
rect 3896 12124 4476 12152
rect 4816 12124 8024 12152
rect 1535 12087 1593 12093
rect 1535 12053 1547 12087
rect 1581 12084 1593 12087
rect 1854 12084 1860 12096
rect 1581 12056 1860 12084
rect 1581 12053 1593 12056
rect 1535 12047 1593 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4338 12084 4344 12096
rect 3927 12056 4344 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4338 12044 4344 12056
rect 4396 12084 4402 12096
rect 4816 12084 4844 12124
rect 8018 12112 8024 12124
rect 8076 12112 8082 12164
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12152 9183 12155
rect 9217 12155 9275 12161
rect 9217 12152 9229 12155
rect 9171 12124 9229 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9217 12121 9229 12124
rect 9263 12152 9275 12155
rect 9490 12152 9496 12164
rect 9263 12124 9496 12152
rect 9263 12121 9275 12124
rect 9217 12115 9275 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 7650 12084 7656 12096
rect 4396 12056 4844 12084
rect 7611 12056 7656 12084
rect 4396 12044 4402 12056
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 7892 12056 8677 12084
rect 7892 12044 7898 12056
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8665 12047 8723 12053
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 10134 12084 10140 12096
rect 9447 12056 10140 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 10870 12084 10876 12096
rect 10827 12056 10876 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13136 12056 13277 12084
rect 13136 12044 13142 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 3145 11883 3203 11889
rect 3145 11849 3157 11883
rect 3191 11880 3203 11883
rect 3234 11880 3240 11892
rect 3191 11852 3240 11880
rect 3191 11849 3203 11852
rect 3145 11843 3203 11849
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 4246 11880 4252 11892
rect 4207 11852 4252 11880
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6730 11880 6736 11892
rect 5951 11852 6736 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6730 11840 6736 11852
rect 6788 11840 6794 11892
rect 8110 11880 8116 11892
rect 8071 11852 8116 11880
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 9692 11852 13645 11880
rect 2774 11812 2780 11824
rect 2687 11784 2780 11812
rect 2774 11772 2780 11784
rect 2832 11812 2838 11824
rect 7745 11815 7803 11821
rect 7745 11812 7757 11815
rect 2832 11784 7757 11812
rect 2832 11772 2838 11784
rect 7745 11781 7757 11784
rect 7791 11781 7803 11815
rect 7745 11775 7803 11781
rect 1762 11744 1768 11756
rect 1723 11716 1768 11744
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11744 2562 11756
rect 3602 11744 3608 11756
rect 2556 11716 3608 11744
rect 2556 11704 2562 11716
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4948 11716 5181 11744
rect 4948 11704 4954 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 6273 11747 6331 11753
rect 6273 11744 6285 11747
rect 5316 11716 6285 11744
rect 5316 11704 5322 11716
rect 6273 11713 6285 11716
rect 6319 11744 6331 11747
rect 6638 11744 6644 11756
rect 6319 11716 6644 11744
rect 6319 11713 6331 11716
rect 6273 11707 6331 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 9692 11744 9720 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 13814 11880 13820 11892
rect 13780 11852 13820 11880
rect 13780 11840 13786 11852
rect 13814 11840 13820 11852
rect 13872 11880 13878 11892
rect 13872 11852 13965 11880
rect 13872 11840 13878 11852
rect 10042 11772 10048 11824
rect 10100 11812 10106 11824
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10100 11784 10793 11812
rect 10100 11772 10106 11784
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 12253 11815 12311 11821
rect 12253 11781 12265 11815
rect 12299 11812 12311 11815
rect 12713 11815 12771 11821
rect 12713 11812 12725 11815
rect 12299 11784 12725 11812
rect 12299 11781 12311 11784
rect 12253 11775 12311 11781
rect 12713 11781 12725 11784
rect 12759 11812 12771 11815
rect 12894 11812 12900 11824
rect 12759 11784 12900 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13449 11815 13507 11821
rect 13449 11812 13461 11815
rect 13228 11784 13461 11812
rect 13228 11772 13234 11784
rect 13449 11781 13461 11784
rect 13495 11781 13507 11815
rect 13449 11775 13507 11781
rect 7484 11716 9720 11744
rect 9769 11747 9827 11753
rect 7484 11676 7512 11716
rect 9769 11713 9781 11747
rect 9815 11744 9827 11747
rect 10870 11744 10876 11756
rect 9815 11716 10876 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10870 11704 10876 11716
rect 10928 11744 10934 11756
rect 11974 11744 11980 11756
rect 10928 11716 11980 11744
rect 10928 11704 10934 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11744 12127 11747
rect 12584 11747 12642 11753
rect 12584 11744 12596 11747
rect 12115 11716 12596 11744
rect 12115 11713 12127 11716
rect 12069 11707 12127 11713
rect 12584 11713 12596 11716
rect 12630 11713 12642 11747
rect 12584 11707 12642 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 12986 11744 12992 11756
rect 12851 11716 12992 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 7024 11648 7512 11676
rect 8481 11679 8539 11685
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 1946 11608 1952 11620
rect 1903 11580 1952 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 1946 11568 1952 11580
rect 2004 11568 2010 11620
rect 3326 11608 3332 11620
rect 3287 11580 3332 11608
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 3421 11611 3479 11617
rect 3421 11577 3433 11611
rect 3467 11577 3479 11611
rect 4890 11608 4896 11620
rect 4851 11580 4896 11608
rect 3421 11571 3479 11577
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 3436 11540 3464 11571
rect 4890 11568 4896 11580
rect 4948 11568 4954 11620
rect 4985 11611 5043 11617
rect 4985 11577 4997 11611
rect 5031 11608 5043 11611
rect 5994 11608 6000 11620
rect 5031 11580 6000 11608
rect 5031 11577 5043 11580
rect 4985 11571 5043 11577
rect 5994 11568 6000 11580
rect 6052 11568 6058 11620
rect 7024 11608 7052 11648
rect 8481 11645 8493 11679
rect 8527 11676 8539 11679
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8527 11648 8861 11676
rect 8527 11645 8539 11648
rect 8481 11639 8539 11645
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 6104 11580 7052 11608
rect 7146 11611 7204 11617
rect 3292 11512 3464 11540
rect 3292 11500 3298 11512
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4212 11512 4721 11540
rect 4212 11500 4218 11512
rect 4709 11509 4721 11512
rect 4755 11540 4767 11543
rect 6104 11540 6132 11580
rect 7146 11577 7158 11611
rect 7192 11577 7204 11611
rect 8864 11608 8892 11639
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 9180 11648 9413 11676
rect 9180 11636 9186 11648
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9674 11676 9680 11688
rect 9631 11648 9680 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10652 11679 10710 11685
rect 10652 11645 10664 11679
rect 10698 11645 10710 11679
rect 10652 11639 10710 11645
rect 9214 11608 9220 11620
rect 8864 11580 9220 11608
rect 7146 11571 7204 11577
rect 6546 11540 6552 11552
rect 4755 11512 6132 11540
rect 6507 11512 6552 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 6546 11500 6552 11512
rect 6604 11540 6610 11552
rect 7161 11540 7189 11571
rect 9214 11568 9220 11580
rect 9272 11608 9278 11620
rect 10520 11608 10548 11636
rect 9272 11580 10548 11608
rect 9272 11568 9278 11580
rect 6604 11512 7189 11540
rect 6604 11500 6610 11512
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 8536 11512 8677 11540
rect 8536 11500 8542 11512
rect 8665 11509 8677 11512
rect 8711 11509 8723 11543
rect 8665 11503 8723 11509
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9088 11512 9781 11540
rect 9088 11500 9094 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 9769 11503 9827 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10667 11540 10695 11639
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11204 11648 12449 11676
rect 11204 11636 11210 11648
rect 12437 11645 12449 11648
rect 12483 11676 12495 11679
rect 13078 11676 13084 11688
rect 12483 11648 13084 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 14052 11679 14110 11685
rect 14052 11676 14064 11679
rect 13228 11648 14064 11676
rect 13228 11636 13234 11648
rect 14052 11645 14064 11648
rect 14098 11676 14110 11679
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14098 11648 14473 11676
rect 14098 11645 14110 11648
rect 14052 11639 14110 11645
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 11238 11608 11244 11620
rect 11199 11580 11244 11608
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 14139 11611 14197 11617
rect 14139 11608 14151 11611
rect 13320 11580 14151 11608
rect 13320 11568 13326 11580
rect 14139 11577 14151 11580
rect 14185 11577 14197 11611
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14139 11571 14197 11577
rect 14246 11580 15025 11608
rect 11054 11540 11060 11552
rect 10459 11512 11060 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11664 11512 11805 11540
rect 11664 11500 11670 11512
rect 11793 11509 11805 11512
rect 11839 11540 11851 11543
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 11839 11512 12081 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 12069 11503 12127 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13633 11543 13691 11549
rect 13633 11509 13645 11543
rect 13679 11540 13691 11543
rect 14246 11540 14274 11580
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15013 11571 15071 11577
rect 13679 11512 14274 11540
rect 13679 11509 13691 11512
rect 13633 11503 13691 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 3602 11336 3608 11348
rect 3563 11308 3608 11336
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 4126 11308 4721 11336
rect 2038 11268 2044 11280
rect 1999 11240 2044 11268
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11268 2651 11271
rect 2774 11268 2780 11280
rect 2639 11240 2780 11268
rect 2639 11237 2651 11240
rect 2593 11231 2651 11237
rect 2774 11228 2780 11240
rect 2832 11268 2838 11280
rect 4126 11268 4154 11308
rect 4709 11305 4721 11308
rect 4755 11336 4767 11339
rect 4890 11336 4896 11348
rect 4755 11308 4896 11336
rect 4755 11305 4767 11308
rect 4709 11299 4767 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 5994 11336 6000 11348
rect 5767 11308 6000 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 6788 11308 8033 11336
rect 6788 11296 6794 11308
rect 8021 11305 8033 11308
rect 8067 11336 8079 11339
rect 8846 11336 8852 11348
rect 8067 11308 8852 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 10137 11339 10195 11345
rect 10137 11336 10149 11339
rect 9732 11308 10149 11336
rect 9732 11296 9738 11308
rect 10137 11305 10149 11308
rect 10183 11305 10195 11339
rect 10137 11299 10195 11305
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11756 11308 11989 11336
rect 11756 11296 11762 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 12342 11336 12348 11348
rect 12303 11308 12348 11336
rect 11977 11299 12035 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 2832 11240 4154 11268
rect 2832 11228 2838 11240
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6962 11271 7020 11277
rect 6962 11268 6974 11271
rect 6604 11240 6974 11268
rect 6604 11228 6610 11240
rect 6962 11237 6974 11240
rect 7008 11237 7020 11271
rect 6962 11231 7020 11237
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11268 9551 11271
rect 13078 11268 13084 11280
rect 9539 11240 13084 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 3292 11172 7573 11200
rect 3292 11160 3298 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 7561 11163 7619 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9968 11209 9996 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10778 11200 10784 11212
rect 10643 11172 10784 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11514 11200 11520 11212
rect 11475 11172 11520 11200
rect 11241 11163 11299 11169
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 4798 11132 4804 11144
rect 4759 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 8386 11132 8392 11144
rect 8299 11104 8392 11132
rect 6641 11095 6699 11101
rect 6549 11067 6607 11073
rect 6549 11033 6561 11067
rect 6595 11064 6607 11067
rect 6656 11064 6684 11095
rect 8386 11092 8392 11104
rect 8444 11132 8450 11144
rect 8444 11104 8800 11132
rect 8444 11092 8450 11104
rect 8478 11064 8484 11076
rect 6595 11036 8484 11064
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 8772 11073 8800 11104
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 11256 11132 11284 11163
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13630 11200 13636 11212
rect 13219 11172 13636 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14090 11200 14096 11212
rect 14051 11172 14096 11200
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15356 11203 15414 11209
rect 15356 11169 15368 11203
rect 15402 11200 15414 11203
rect 15470 11200 15476 11212
rect 15402 11172 15476 11200
rect 15402 11169 15414 11172
rect 15356 11163 15414 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 11422 11132 11428 11144
rect 9640 11104 11428 11132
rect 9640 11092 9646 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11698 11132 11704 11144
rect 11659 11104 11704 11132
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 11940 11104 12541 11132
rect 11940 11092 11946 11104
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 8757 11067 8815 11073
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 9306 11064 9312 11076
rect 8803 11036 9312 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 10928 11036 12940 11064
rect 10928 11024 10934 11036
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 2869 10999 2927 11005
rect 2869 10996 2881 10999
rect 1912 10968 2881 10996
rect 1912 10956 1918 10968
rect 2869 10965 2881 10968
rect 2915 10965 2927 10999
rect 3326 10996 3332 11008
rect 3287 10968 3332 10996
rect 2869 10959 2927 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 9122 10996 9128 11008
rect 9083 10968 9128 10996
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 12912 10996 12940 11036
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 15427 11067 15485 11073
rect 15427 11064 15439 11067
rect 13596 11036 15439 11064
rect 13596 11024 13602 11036
rect 15427 11033 15439 11036
rect 15473 11033 15485 11067
rect 15427 11027 15485 11033
rect 14231 10999 14289 11005
rect 14231 10996 14243 10999
rect 12912 10968 14243 10996
rect 14231 10965 14243 10968
rect 14277 10965 14289 10999
rect 14231 10959 14289 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1946 10752 1952 10804
rect 2004 10792 2010 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 2004 10764 3433 10792
rect 2004 10752 2010 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 3421 10755 3479 10761
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 7708 10764 10425 10792
rect 7708 10752 7714 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 10413 10755 10471 10761
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11422 10792 11428 10804
rect 11103 10764 11428 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 2222 10684 2228 10736
rect 2280 10724 2286 10736
rect 3145 10727 3203 10733
rect 3145 10724 3157 10727
rect 2280 10696 3157 10724
rect 2280 10684 2286 10696
rect 3145 10693 3157 10696
rect 3191 10724 3203 10727
rect 5994 10724 6000 10736
rect 3191 10696 6000 10724
rect 3191 10693 3203 10696
rect 3145 10687 3203 10693
rect 5994 10684 6000 10696
rect 6052 10684 6058 10736
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 8628 10696 9505 10724
rect 8628 10684 8634 10696
rect 9493 10693 9505 10696
rect 9539 10724 9551 10727
rect 10134 10724 10140 10736
rect 9539 10696 10140 10724
rect 9539 10693 9551 10696
rect 9493 10687 9551 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10778 10724 10784 10736
rect 10284 10696 10784 10724
rect 10284 10684 10290 10696
rect 10778 10684 10784 10696
rect 10836 10684 10842 10736
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 14090 10724 14096 10736
rect 11020 10696 14096 10724
rect 11020 10684 11026 10696
rect 14090 10684 14096 10696
rect 14148 10724 14154 10736
rect 14645 10727 14703 10733
rect 14645 10724 14657 10727
rect 14148 10696 14657 10724
rect 14148 10684 14154 10696
rect 14645 10693 14657 10696
rect 14691 10693 14703 10727
rect 14645 10687 14703 10693
rect 2774 10656 2780 10668
rect 2735 10628 2780 10656
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5868 10628 6285 10656
rect 5868 10616 5874 10628
rect 6273 10625 6285 10628
rect 6319 10656 6331 10659
rect 6319 10628 7420 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 7392 10600 7420 10628
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 9398 10656 9404 10668
rect 7616 10628 9404 10656
rect 7616 10616 7622 10628
rect 9398 10616 9404 10628
rect 9456 10656 9462 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 9456 10628 10333 10656
rect 9456 10616 9462 10628
rect 10321 10625 10333 10628
rect 10367 10656 10379 10659
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10367 10628 11345 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 11333 10625 11345 10628
rect 11379 10656 11391 10659
rect 11379 10628 13814 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 3640 10591 3698 10597
rect 3640 10588 3652 10591
rect 3476 10560 3652 10588
rect 3476 10548 3482 10560
rect 3640 10557 3652 10560
rect 3686 10588 3698 10591
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 3686 10560 4077 10588
rect 3686 10557 3698 10560
rect 3640 10551 3698 10557
rect 4065 10557 4077 10560
rect 4111 10557 4123 10591
rect 4065 10551 4123 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 4571 10560 4997 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4985 10557 4997 10560
rect 5031 10588 5043 10591
rect 7101 10591 7159 10597
rect 5031 10560 6684 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 1302 10480 1308 10532
rect 1360 10520 1366 10532
rect 1854 10520 1860 10532
rect 1360 10492 1860 10520
rect 1360 10480 1366 10492
rect 1854 10480 1860 10492
rect 1912 10520 1918 10532
rect 2133 10523 2191 10529
rect 2133 10520 2145 10523
rect 1912 10492 2145 10520
rect 1912 10480 1918 10492
rect 2133 10489 2145 10492
rect 2179 10489 2191 10523
rect 2133 10483 2191 10489
rect 2222 10480 2228 10532
rect 2280 10520 2286 10532
rect 5166 10520 5172 10532
rect 2280 10492 2325 10520
rect 4816 10492 5172 10520
rect 2280 10480 2286 10492
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 2038 10452 2044 10464
rect 1995 10424 2044 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 2038 10412 2044 10424
rect 2096 10452 2102 10464
rect 2406 10452 2412 10464
rect 2096 10424 2412 10452
rect 2096 10412 2102 10424
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3743 10455 3801 10461
rect 3743 10452 3755 10455
rect 3568 10424 3755 10452
rect 3568 10412 3574 10424
rect 3743 10421 3755 10424
rect 3789 10421 3801 10455
rect 3743 10415 3801 10421
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4816 10461 4844 10492
rect 5166 10480 5172 10492
rect 5224 10520 5230 10532
rect 5306 10523 5364 10529
rect 5306 10520 5318 10523
rect 5224 10492 5318 10520
rect 5224 10480 5230 10492
rect 5306 10489 5318 10492
rect 5352 10520 5364 10523
rect 6546 10520 6552 10532
rect 5352 10492 6552 10520
rect 5352 10489 5364 10492
rect 5306 10483 5364 10489
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 4801 10455 4859 10461
rect 4801 10452 4813 10455
rect 4580 10424 4813 10452
rect 4580 10412 4586 10424
rect 4801 10421 4813 10424
rect 4847 10421 4859 10455
rect 4801 10415 4859 10421
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 5994 10452 6000 10464
rect 5951 10424 6000 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6656 10452 6684 10560
rect 7101 10557 7113 10591
rect 7147 10557 7159 10591
rect 7374 10588 7380 10600
rect 7335 10560 7380 10588
rect 7101 10551 7159 10557
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7116 10520 7144 10551
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 8386 10588 8392 10600
rect 8347 10560 8392 10588
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8846 10588 8852 10600
rect 8807 10560 8852 10588
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 10100 10591 10158 10597
rect 10100 10588 10112 10591
rect 9548 10560 10112 10588
rect 9548 10548 9554 10560
rect 10100 10557 10112 10560
rect 10146 10557 10158 10591
rect 10100 10551 10158 10557
rect 12253 10591 12311 10597
rect 12253 10557 12265 10591
rect 12299 10588 12311 10591
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12299 10560 12725 10588
rect 12299 10557 12311 10560
rect 12253 10551 12311 10557
rect 12713 10557 12725 10560
rect 12759 10588 12771 10591
rect 13354 10588 13360 10600
rect 12759 10560 13360 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13786 10588 13814 10628
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14608 10628 15275 10656
rect 14608 10616 14614 10628
rect 15247 10597 15275 10628
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13786 10560 14197 10588
rect 14185 10557 14197 10560
rect 14231 10588 14243 10591
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14231 10560 15025 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15232 10591 15290 10597
rect 15232 10557 15244 10591
rect 15278 10588 15290 10591
rect 15657 10591 15715 10597
rect 15657 10588 15669 10591
rect 15278 10560 15669 10588
rect 15278 10557 15290 10560
rect 15232 10551 15290 10557
rect 15657 10557 15669 10560
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16244 10591 16302 10597
rect 16244 10588 16256 10591
rect 15896 10560 16256 10588
rect 15896 10548 15902 10560
rect 16244 10557 16256 10560
rect 16290 10588 16302 10591
rect 16669 10591 16727 10597
rect 16669 10588 16681 10591
rect 16290 10560 16681 10588
rect 16290 10557 16302 10560
rect 16244 10551 16302 10557
rect 16669 10557 16681 10560
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 8404 10520 8432 10548
rect 6788 10492 8432 10520
rect 9953 10523 10011 10529
rect 6788 10480 6794 10492
rect 9953 10489 9965 10523
rect 9999 10520 10011 10523
rect 10686 10520 10692 10532
rect 9999 10492 10692 10520
rect 9999 10489 10011 10492
rect 9953 10483 10011 10489
rect 10686 10480 10692 10492
rect 10744 10520 10750 10532
rect 11790 10520 11796 10532
rect 10744 10492 11796 10520
rect 10744 10480 10750 10492
rect 11790 10480 11796 10492
rect 11848 10480 11854 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12032 10492 14095 10520
rect 12032 10480 12038 10492
rect 6917 10455 6975 10461
rect 6917 10452 6929 10455
rect 6656 10424 6929 10452
rect 6917 10421 6929 10424
rect 6963 10421 6975 10455
rect 6917 10415 6975 10421
rect 7834 10412 7840 10464
rect 7892 10452 7898 10464
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7892 10424 8033 10452
rect 7892 10412 7898 10424
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 8021 10415 8079 10421
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11572 10424 11713 10452
rect 11572 10412 11578 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 11701 10415 11759 10421
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 14067 10452 14095 10492
rect 14734 10480 14740 10532
rect 14792 10520 14798 10532
rect 15470 10520 15476 10532
rect 14792 10492 15476 10520
rect 14792 10480 14798 10492
rect 15470 10480 15476 10492
rect 15528 10520 15534 10532
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 15528 10492 16037 10520
rect 15528 10480 15534 10492
rect 16025 10489 16037 10492
rect 16071 10489 16083 10523
rect 16025 10483 16083 10489
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14067 10424 14381 10452
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14369 10415 14427 10421
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15335 10455 15393 10461
rect 15335 10452 15347 10455
rect 14516 10424 15347 10452
rect 14516 10412 14522 10424
rect 15335 10421 15347 10424
rect 15381 10421 15393 10455
rect 15335 10415 15393 10421
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16347 10455 16405 10461
rect 16347 10452 16359 10455
rect 15712 10424 16359 10452
rect 15712 10412 15718 10424
rect 16347 10421 16359 10424
rect 16393 10421 16405 10455
rect 16347 10415 16405 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3510 10248 3516 10260
rect 2731 10220 3516 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 1670 10140 1676 10192
rect 1728 10180 1734 10192
rect 1765 10183 1823 10189
rect 1765 10180 1777 10183
rect 1728 10152 1777 10180
rect 1728 10140 1734 10152
rect 1765 10149 1777 10152
rect 1811 10149 1823 10183
rect 1765 10143 1823 10149
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 2700 10044 2728 10211
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4203 10251 4261 10257
rect 4203 10248 4215 10251
rect 3936 10220 4215 10248
rect 3936 10208 3942 10220
rect 4203 10217 4215 10220
rect 4249 10217 4261 10251
rect 4203 10211 4261 10217
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4798 10248 4804 10260
rect 4755 10220 4804 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4798 10208 4804 10220
rect 4856 10248 4862 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4856 10220 5365 10248
rect 4856 10208 4862 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 6730 10248 6736 10260
rect 6691 10220 6736 10248
rect 5353 10211 5411 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8444 10220 9137 10248
rect 8444 10208 8450 10220
rect 9125 10217 9137 10220
rect 9171 10248 9183 10251
rect 9306 10248 9312 10260
rect 9171 10220 9312 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9306 10208 9312 10220
rect 9364 10248 9370 10260
rect 10686 10248 10692 10260
rect 9364 10220 10692 10248
rect 9364 10208 9370 10220
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11146 10248 11152 10260
rect 11107 10220 11152 10248
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 13630 10248 13636 10260
rect 11256 10220 13636 10248
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 8846 10180 8852 10192
rect 8803 10152 8852 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 11256 10180 11284 10220
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 8996 10152 11284 10180
rect 8996 10140 9002 10152
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 11572 10152 13308 10180
rect 11572 10140 11578 10152
rect 3881 10115 3939 10121
rect 3881 10081 3893 10115
rect 3927 10112 3939 10115
rect 4111 10115 4169 10121
rect 4111 10112 4123 10115
rect 3927 10084 4123 10112
rect 3927 10081 3939 10084
rect 3881 10075 3939 10081
rect 4111 10081 4123 10084
rect 4157 10112 4169 10115
rect 5074 10112 5080 10124
rect 4157 10084 5080 10112
rect 4157 10081 4169 10084
rect 4111 10075 4169 10081
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5258 10112 5264 10124
rect 5219 10084 5264 10112
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5810 10112 5816 10124
rect 5408 10084 5816 10112
rect 5408 10072 5414 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7984 10084 8033 10112
rect 7984 10072 7990 10084
rect 8021 10081 8033 10084
rect 8067 10112 8079 10115
rect 9398 10112 9404 10124
rect 8067 10084 9404 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 9398 10072 9404 10084
rect 9456 10112 9462 10124
rect 9950 10112 9956 10124
rect 9456 10084 9956 10112
rect 9456 10072 9462 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10134 10112 10140 10124
rect 10095 10084 10140 10112
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11422 10112 11428 10124
rect 11383 10084 11428 10112
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 12250 10112 12256 10124
rect 11839 10084 12256 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 13078 10112 13084 10124
rect 13039 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13280 10121 13308 10152
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13630 10112 13636 10124
rect 13311 10084 13636 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 16368 10115 16426 10121
rect 16368 10081 16380 10115
rect 16414 10112 16426 10115
rect 16482 10112 16488 10124
rect 16414 10084 16488 10112
rect 16414 10081 16426 10084
rect 16368 10075 16426 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 6822 10044 6828 10056
rect 1719 10016 2728 10044
rect 6783 10016 6828 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7708 10016 7849 10044
rect 7708 10004 7714 10016
rect 7837 10013 7849 10016
rect 7883 10044 7895 10047
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 7883 10016 8401 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 8389 10013 8401 10016
rect 8435 10044 8447 10047
rect 9030 10044 9036 10056
rect 8435 10016 9036 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 11974 10044 11980 10056
rect 11935 10016 11980 10044
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 13538 10044 13544 10056
rect 13499 10016 13544 10044
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15378 10044 15384 10056
rect 15335 10016 15384 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 2314 9976 2320 9988
rect 2271 9948 2320 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 2314 9936 2320 9948
rect 2372 9976 2378 9988
rect 2961 9979 3019 9985
rect 2961 9976 2973 9979
rect 2372 9948 2973 9976
rect 2372 9936 2378 9948
rect 2961 9945 2973 9948
rect 3007 9945 3019 9979
rect 2961 9939 3019 9945
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 11882 9976 11888 9988
rect 5500 9948 11888 9976
rect 5500 9936 5506 9948
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4580 9880 4997 9908
rect 4580 9868 4586 9880
rect 4985 9877 4997 9880
rect 5031 9877 5043 9911
rect 4985 9871 5043 9877
rect 7561 9911 7619 9917
rect 7561 9877 7573 9911
rect 7607 9908 7619 9911
rect 7834 9908 7840 9920
rect 7607 9880 7840 9908
rect 7607 9877 7619 9880
rect 7561 9871 7619 9877
rect 7834 9868 7840 9880
rect 7892 9908 7898 9920
rect 8159 9911 8217 9917
rect 8159 9908 8171 9911
rect 7892 9880 8171 9908
rect 7892 9868 7898 9880
rect 8159 9877 8171 9880
rect 8205 9877 8217 9911
rect 8159 9871 8217 9877
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8662 9908 8668 9920
rect 8343 9880 8668 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 9490 9908 9496 9920
rect 9451 9880 9496 9908
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 10778 9908 10784 9920
rect 10691 9880 10784 9908
rect 10778 9868 10784 9880
rect 10836 9908 10842 9920
rect 11790 9908 11796 9920
rect 10836 9880 11796 9908
rect 10836 9868 10842 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 16439 9911 16497 9917
rect 16439 9877 16451 9911
rect 16485 9908 16497 9911
rect 16574 9908 16580 9920
rect 16485 9880 16580 9908
rect 16485 9877 16497 9880
rect 16439 9871 16497 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5077 9707 5135 9713
rect 5077 9673 5089 9707
rect 5123 9704 5135 9707
rect 5258 9704 5264 9716
rect 5123 9676 5264 9704
rect 5123 9673 5135 9676
rect 5077 9667 5135 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 8849 9707 8907 9713
rect 8849 9704 8861 9707
rect 7432 9676 8861 9704
rect 7432 9664 7438 9676
rect 8849 9673 8861 9676
rect 8895 9673 8907 9707
rect 8849 9667 8907 9673
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 9548 9676 10609 9704
rect 9548 9664 9554 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 10597 9667 10655 9673
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11609 9707 11667 9713
rect 11609 9704 11621 9707
rect 11480 9676 11621 9704
rect 11480 9664 11486 9676
rect 11609 9673 11621 9676
rect 11655 9704 11667 9707
rect 12158 9704 12164 9716
rect 11655 9676 12164 9704
rect 11655 9673 11667 9676
rect 11609 9667 11667 9673
rect 12158 9664 12164 9676
rect 12216 9704 12222 9716
rect 13078 9704 13084 9716
rect 12216 9676 13084 9704
rect 12216 9664 12222 9676
rect 13078 9664 13084 9676
rect 13136 9704 13142 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 13136 9676 13277 9704
rect 13136 9664 13142 9676
rect 13265 9673 13277 9676
rect 13311 9673 13323 9707
rect 13265 9667 13323 9673
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2148 9608 3157 9636
rect 2148 9577 2176 9608
rect 3145 9605 3157 9608
rect 3191 9636 3203 9639
rect 6822 9636 6828 9648
rect 3191 9608 6828 9636
rect 3191 9605 3203 9608
rect 3145 9599 3203 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7834 9596 7840 9648
rect 7892 9636 7898 9648
rect 8527 9639 8585 9645
rect 8527 9636 8539 9639
rect 7892 9608 8539 9636
rect 7892 9596 7898 9608
rect 8527 9605 8539 9608
rect 8573 9605 8585 9639
rect 8662 9636 8668 9648
rect 8623 9608 8668 9636
rect 8527 9599 8585 9605
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13688 9608 13829 9636
rect 13688 9596 13694 9608
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 2222 9528 2228 9580
rect 2280 9568 2286 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2280 9540 2421 9568
rect 2280 9528 2286 9540
rect 2409 9537 2421 9540
rect 2455 9568 2467 9571
rect 2590 9568 2596 9580
rect 2455 9540 2596 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8680 9568 8708 9596
rect 8159 9540 8708 9568
rect 8757 9571 8815 9577
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9030 9568 9036 9580
rect 8803 9540 9036 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10459 9540 11284 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3476 9472 3617 9500
rect 3476 9460 3482 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4709 9503 4767 9509
rect 4212 9472 4257 9500
rect 4212 9460 4218 9472
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 4755 9472 5825 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 5813 9469 5825 9472
rect 5859 9500 5871 9503
rect 5994 9500 6000 9512
rect 5859 9472 6000 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7466 9500 7472 9512
rect 6687 9472 7472 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8386 9500 8392 9512
rect 8347 9472 8392 9500
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 11256 9509 11284 9540
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 12676 9540 14013 9568
rect 12676 9528 12682 9540
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 10781 9503 10839 9509
rect 10781 9469 10793 9503
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11606 9500 11612 9512
rect 11287 9472 11612 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 2130 9392 2136 9444
rect 2188 9432 2194 9444
rect 2225 9435 2283 9441
rect 2225 9432 2237 9435
rect 2188 9404 2237 9432
rect 2188 9392 2194 9404
rect 2225 9401 2237 9404
rect 2271 9401 2283 9435
rect 2225 9395 2283 9401
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 5169 9435 5227 9441
rect 5169 9432 5181 9435
rect 2464 9404 5181 9432
rect 2464 9392 2470 9404
rect 5169 9401 5181 9404
rect 5215 9401 5227 9435
rect 10796 9432 10824 9463
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12584 9472 12909 9500
rect 12584 9460 12590 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 15470 9500 15476 9512
rect 15383 9472 15476 9500
rect 14093 9463 14151 9469
rect 11146 9432 11152 9444
rect 10796 9404 11152 9432
rect 5169 9395 5227 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 13170 9432 13176 9444
rect 13131 9404 13176 9432
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14108 9432 14136 9463
rect 15470 9460 15476 9472
rect 15528 9500 15534 9512
rect 15657 9503 15715 9509
rect 15657 9500 15669 9503
rect 15528 9472 15669 9500
rect 15528 9460 15534 9472
rect 15657 9469 15669 9472
rect 15703 9469 15715 9503
rect 15657 9463 15715 9469
rect 15562 9432 15568 9444
rect 14056 9404 14136 9432
rect 15523 9404 15568 9432
rect 14056 9392 14062 9404
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 18230 9432 18236 9444
rect 16408 9404 18236 9432
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3878 9364 3884 9376
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9364 9827 9367
rect 10134 9364 10140 9376
rect 9815 9336 10140 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12250 9364 12256 9376
rect 12023 9336 12256 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13311 9336 13553 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13541 9333 13553 9336
rect 13587 9364 13599 9367
rect 16408 9364 16436 9404
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 13587 9336 16436 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16577 9367 16635 9373
rect 16577 9364 16589 9367
rect 16540 9336 16589 9364
rect 16540 9324 16546 9336
rect 16577 9333 16589 9336
rect 16623 9333 16635 9367
rect 16577 9327 16635 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 5350 9160 5356 9172
rect 5311 9132 5356 9160
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 7561 9163 7619 9169
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 7650 9160 7656 9172
rect 7607 9132 7656 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 7926 9160 7932 9172
rect 7887 9132 7932 9160
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8849 9163 8907 9169
rect 8849 9129 8861 9163
rect 8895 9160 8907 9163
rect 9125 9163 9183 9169
rect 9125 9160 9137 9163
rect 8895 9132 9137 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 9125 9129 9137 9132
rect 9171 9160 9183 9163
rect 10781 9163 10839 9169
rect 9171 9132 9996 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2498 9092 2504 9104
rect 2455 9064 2504 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 4427 9095 4485 9101
rect 4427 9061 4439 9095
rect 4473 9092 4485 9095
rect 4522 9092 4528 9104
rect 4473 9064 4528 9092
rect 4473 9061 4485 9064
rect 4427 9055 4485 9061
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 5997 9095 6055 9101
rect 5997 9061 6009 9095
rect 6043 9092 6055 9095
rect 6270 9092 6276 9104
rect 6043 9064 6276 9092
rect 6043 9061 6055 9064
rect 5997 9055 6055 9061
rect 6270 9052 6276 9064
rect 6328 9092 6334 9104
rect 9858 9092 9864 9104
rect 6328 9064 9864 9092
rect 6328 9052 6334 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 9968 9092 9996 9132
rect 10781 9129 10793 9163
rect 10827 9160 10839 9163
rect 11330 9160 11336 9172
rect 10827 9132 11336 9160
rect 10827 9129 10839 9132
rect 10781 9123 10839 9129
rect 11330 9120 11336 9132
rect 11388 9160 11394 9172
rect 12526 9160 12532 9172
rect 11388 9132 12532 9160
rect 11388 9120 11394 9132
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12802 9160 12808 9172
rect 12636 9132 12808 9160
rect 12636 9092 12664 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 13872 9132 16896 9160
rect 13872 9120 13878 9132
rect 12894 9092 12900 9104
rect 9968 9064 12664 9092
rect 12855 9064 12900 9092
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13906 9092 13912 9104
rect 13044 9064 13912 9092
rect 13044 9052 13050 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 15470 9092 15476 9104
rect 15431 9064 15476 9092
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3936 8996 4077 9024
rect 3936 8984 3942 8996
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 8662 9024 8668 9036
rect 8575 8996 8668 9024
rect 4065 8987 4123 8993
rect 8662 8984 8668 8996
rect 8720 9024 8726 9036
rect 8849 9027 8907 9033
rect 8849 9024 8861 9027
rect 8720 8996 8861 9024
rect 8720 8984 8726 8996
rect 8849 8993 8861 8996
rect 8895 8993 8907 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 8849 8987 8907 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 11422 9024 11428 9036
rect 11383 8996 11428 9024
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 16868 9033 16896 9132
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 9024 16911 9027
rect 16942 9024 16948 9036
rect 16899 8996 16948 9024
rect 16899 8993 16911 8996
rect 16853 8987 16911 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17932 9027 17990 9033
rect 17932 8993 17944 9027
rect 17978 9024 17990 9027
rect 18414 9024 18420 9036
rect 17978 8996 18420 9024
rect 17978 8993 17990 8996
rect 17932 8987 17990 8993
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18912 9027 18970 9033
rect 18912 8993 18924 9027
rect 18958 8993 18970 9027
rect 18912 8987 18970 8993
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5629 8959 5687 8965
rect 5629 8956 5641 8959
rect 5316 8928 5641 8956
rect 5316 8916 5322 8928
rect 5629 8925 5641 8928
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6546 8956 6552 8968
rect 5951 8928 6552 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 8803 8928 11836 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 11808 8900 11836 8928
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12492 8928 12817 8956
rect 12492 8916 12498 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13630 8956 13636 8968
rect 13495 8928 13636 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 13630 8916 13636 8928
rect 13688 8956 13694 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 13688 8928 15393 8956
rect 13688 8916 13694 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 15381 8919 15439 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 17494 8916 17500 8968
rect 17552 8956 17558 8968
rect 18927 8956 18955 8987
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 17552 8928 19349 8956
rect 17552 8916 17558 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 2958 8848 2964 8900
rect 3016 8888 3022 8900
rect 3697 8891 3755 8897
rect 3697 8888 3709 8891
rect 3016 8860 3709 8888
rect 3016 8848 3022 8860
rect 3697 8857 3709 8860
rect 3743 8888 3755 8891
rect 4154 8888 4160 8900
rect 3743 8860 4160 8888
rect 3743 8857 3755 8860
rect 3697 8851 3755 8857
rect 4154 8848 4160 8860
rect 4212 8888 4218 8900
rect 4890 8888 4896 8900
rect 4212 8860 4896 8888
rect 4212 8848 4218 8860
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 5132 8860 6469 8888
rect 5132 8848 5138 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 9122 8848 9128 8900
rect 9180 8888 9186 8900
rect 9861 8891 9919 8897
rect 9861 8888 9873 8891
rect 9180 8860 9873 8888
rect 9180 8848 9186 8860
rect 9861 8857 9873 8860
rect 9907 8857 9919 8891
rect 11146 8888 11152 8900
rect 11107 8860 11152 8888
rect 9861 8851 9919 8857
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 11790 8848 11796 8900
rect 11848 8888 11854 8900
rect 13814 8888 13820 8900
rect 11848 8860 13820 8888
rect 11848 8848 11854 8860
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 13924 8860 14228 8888
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 1946 8820 1952 8832
rect 1811 8792 1952 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2130 8820 2136 8832
rect 2091 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3200 8792 3249 8820
rect 3200 8780 3206 8792
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 4982 8820 4988 8832
rect 4943 8792 4988 8820
rect 3237 8783 3295 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 12342 8820 12348 8832
rect 5224 8792 12348 8820
rect 5224 8780 5230 8792
rect 12342 8780 12348 8792
rect 12400 8820 12406 8832
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 12400 8792 12449 8820
rect 12400 8780 12406 8792
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13924 8820 13952 8860
rect 12584 8792 13952 8820
rect 12584 8780 12590 8792
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14200 8820 14228 8860
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 14056 8792 14101 8820
rect 14200 8792 17049 8820
rect 14056 8780 14062 8792
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17037 8783 17095 8789
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 18003 8823 18061 8829
rect 18003 8820 18015 8823
rect 17184 8792 18015 8820
rect 17184 8780 17190 8792
rect 18003 8789 18015 8792
rect 18049 8789 18061 8823
rect 18003 8783 18061 8789
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19015 8823 19073 8829
rect 19015 8820 19027 8823
rect 18932 8792 19027 8820
rect 18932 8780 18938 8792
rect 19015 8789 19027 8792
rect 19061 8789 19073 8823
rect 19015 8783 19073 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 4982 8616 4988 8628
rect 2556 8588 4988 8616
rect 2556 8576 2562 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 6270 8616 6276 8628
rect 6231 8588 6276 8616
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6546 8616 6552 8628
rect 6507 8588 6552 8616
rect 6546 8576 6552 8588
rect 6604 8616 6610 8628
rect 8113 8619 8171 8625
rect 6604 8588 6868 8616
rect 6604 8576 6610 8588
rect 2314 8548 2320 8560
rect 2275 8520 2320 8548
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 4948 8520 5948 8548
rect 4948 8508 4954 8520
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5132 8452 5549 8480
rect 5132 8440 5138 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 3200 8384 3249 8412
rect 3200 8372 3206 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 5920 8412 5948 8520
rect 6840 8489 6868 8588
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8662 8616 8668 8628
rect 8159 8588 8668 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9398 8616 9404 8628
rect 9359 8588 9404 8616
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9824 8588 10057 8616
rect 9824 8576 9830 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 12526 8616 12532 8628
rect 11204 8588 12532 8616
rect 11204 8576 11210 8588
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 15105 8619 15163 8625
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15470 8616 15476 8628
rect 15151 8588 15476 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 18230 8616 18236 8628
rect 18191 8588 18236 8616
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18509 8619 18567 8625
rect 18509 8616 18521 8619
rect 18472 8588 18521 8616
rect 18472 8576 18478 8588
rect 18509 8585 18521 8588
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 7558 8508 7564 8560
rect 7616 8548 7622 8560
rect 7834 8548 7840 8560
rect 7616 8520 7840 8548
rect 7616 8508 7622 8520
rect 7834 8508 7840 8520
rect 7892 8548 7898 8560
rect 8435 8551 8493 8557
rect 8435 8548 8447 8551
rect 7892 8520 8447 8548
rect 7892 8508 7898 8520
rect 8435 8517 8447 8520
rect 8481 8517 8493 8551
rect 8435 8511 8493 8517
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 8846 8548 8852 8560
rect 8619 8520 8852 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 8846 8508 8852 8520
rect 8904 8548 8910 8560
rect 9950 8548 9956 8560
rect 8904 8520 9956 8548
rect 8904 8508 8910 8520
rect 9950 8508 9956 8520
rect 10008 8548 10014 8560
rect 11164 8548 11192 8576
rect 10008 8520 11192 8548
rect 10008 8508 10014 8520
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 19199 8551 19257 8557
rect 19199 8548 19211 8551
rect 12492 8520 19211 8548
rect 12492 8508 12498 8520
rect 19199 8517 19211 8520
rect 19245 8517 19257 8551
rect 19199 8511 19257 8517
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 7524 8452 7757 8480
rect 7524 8440 7530 8452
rect 7745 8449 7757 8452
rect 7791 8480 7803 8483
rect 8662 8480 8668 8492
rect 7791 8452 8668 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 8772 8412 8800 8443
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9732 8452 9781 8480
rect 9732 8440 9738 8452
rect 9769 8449 9781 8452
rect 9815 8480 9827 8483
rect 12986 8480 12992 8492
rect 9815 8452 12992 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13228 8452 13814 8480
rect 13228 8440 13234 8452
rect 5920 8384 8800 8412
rect 3237 8375 3295 8381
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10100 8384 10793 8412
rect 10100 8372 10106 8384
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 11330 8412 11336 8424
rect 11291 8384 11336 8412
rect 10781 8375 10839 8381
rect 1762 8344 1768 8356
rect 1723 8316 1768 8344
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 1946 8344 1952 8356
rect 1903 8316 1952 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 1946 8304 1952 8316
rect 2004 8344 2010 8356
rect 3053 8347 3111 8353
rect 2004 8316 2820 8344
rect 2004 8304 2010 8316
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2685 8279 2743 8285
rect 2685 8276 2697 8279
rect 2648 8248 2697 8276
rect 2648 8236 2654 8248
rect 2685 8245 2697 8248
rect 2731 8245 2743 8279
rect 2792 8276 2820 8316
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3599 8347 3657 8353
rect 3599 8344 3611 8347
rect 3099 8316 3611 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3599 8313 3611 8316
rect 3645 8344 3657 8347
rect 5258 8344 5264 8356
rect 3645 8316 4568 8344
rect 5219 8316 5264 8344
rect 3645 8313 3657 8316
rect 3599 8307 3657 8313
rect 4540 8288 4568 8316
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 6638 8344 6644 8356
rect 5399 8316 6644 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 4157 8279 4215 8285
rect 4157 8276 4169 8279
rect 2792 8248 4169 8276
rect 2685 8239 2743 8245
rect 4157 8245 4169 8248
rect 4203 8245 4215 8279
rect 4522 8276 4528 8288
rect 4483 8248 4528 8276
rect 4157 8239 4215 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5368 8276 5396 8307
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 7926 8304 7932 8356
rect 7984 8344 7990 8356
rect 8294 8344 8300 8356
rect 7984 8316 8300 8344
rect 7984 8304 7990 8316
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 10796 8344 10824 8375
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 11563 8384 12449 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 12437 8381 12449 8384
rect 12483 8412 12495 8415
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 12483 8384 13645 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 13786 8412 13814 8452
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 14792 8452 19150 8480
rect 14792 8440 14798 8452
rect 14182 8412 14188 8424
rect 13786 8384 14188 8412
rect 13633 8375 13691 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 15841 8415 15899 8421
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 15887 8384 16037 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 16025 8381 16037 8384
rect 16071 8412 16083 8415
rect 16206 8412 16212 8424
rect 16071 8384 16212 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 19122 8421 19150 8452
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18877 8415 18935 8421
rect 18877 8412 18889 8415
rect 18095 8384 18889 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18877 8381 18889 8384
rect 18923 8381 18935 8415
rect 18877 8375 18935 8381
rect 19107 8415 19165 8421
rect 19107 8381 19119 8415
rect 19153 8412 19165 8415
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19153 8384 19533 8412
rect 19153 8381 19165 8384
rect 19107 8375 19165 8381
rect 19521 8381 19533 8384
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 10796 8316 11805 8344
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 11793 8307 11851 8313
rect 12253 8347 12311 8353
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 12299 8316 12770 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12758 8313 12770 8316
rect 12804 8344 12816 8347
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 12804 8316 14105 8344
rect 12804 8313 12816 8316
rect 12758 8307 12816 8313
rect 14093 8313 14105 8316
rect 14139 8344 14151 8347
rect 14274 8344 14280 8356
rect 14139 8316 14280 8344
rect 14139 8313 14151 8316
rect 14093 8307 14151 8313
rect 5123 8248 5396 8276
rect 7377 8279 7435 8285
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 7377 8245 7389 8279
rect 7423 8276 7435 8279
rect 8846 8276 8852 8288
rect 7423 8248 8852 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 11422 8276 11428 8288
rect 10735 8248 11428 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 11808 8276 11836 8307
rect 14274 8304 14280 8316
rect 14332 8344 14338 8356
rect 14506 8347 14564 8353
rect 14506 8344 14518 8347
rect 14332 8316 14518 8344
rect 14332 8304 14338 8316
rect 14506 8313 14518 8316
rect 14552 8313 14564 8347
rect 14506 8307 14564 8313
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 15933 8347 15991 8353
rect 15933 8344 15945 8347
rect 15528 8316 15945 8344
rect 15528 8304 15534 8316
rect 15933 8313 15945 8316
rect 15979 8313 15991 8347
rect 15933 8307 15991 8313
rect 13170 8276 13176 8288
rect 11808 8248 13176 8276
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 14366 8236 14372 8288
rect 14424 8276 14430 8288
rect 18064 8276 18092 8375
rect 14424 8248 18092 8276
rect 14424 8236 14430 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4157 8075 4215 8081
rect 4157 8072 4169 8075
rect 4120 8044 4169 8072
rect 4120 8032 4126 8044
rect 4157 8041 4169 8044
rect 4203 8041 4215 8075
rect 4157 8035 4215 8041
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5350 8072 5356 8084
rect 5307 8044 5356 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5350 8032 5356 8044
rect 5408 8072 5414 8084
rect 8386 8072 8392 8084
rect 5408 8044 8392 8072
rect 5408 8032 5414 8044
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 11514 8072 11520 8084
rect 8711 8044 11520 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12434 8072 12440 8084
rect 12395 8044 12440 8072
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 12894 8072 12900 8084
rect 12851 8044 12900 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13909 8075 13967 8081
rect 13909 8072 13921 8075
rect 13228 8044 13921 8072
rect 13228 8032 13234 8044
rect 13909 8041 13921 8044
rect 13955 8041 13967 8075
rect 13909 8035 13967 8041
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 19107 8075 19165 8081
rect 19107 8072 19119 8075
rect 14700 8044 19119 8072
rect 14700 8032 14706 8044
rect 19107 8041 19119 8044
rect 19153 8041 19165 8075
rect 19107 8035 19165 8041
rect 3142 8004 3148 8016
rect 3103 7976 3148 8004
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 6083 8007 6141 8013
rect 6083 8004 6095 8007
rect 4580 7976 6095 8004
rect 4580 7964 4586 7976
rect 6083 7973 6095 7976
rect 6129 8004 6141 8007
rect 6178 8004 6184 8016
rect 6129 7976 6184 8004
rect 6129 7973 6141 7976
rect 6083 7967 6141 7973
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 10597 8007 10655 8013
rect 9088 7976 10272 8004
rect 9088 7964 9094 7976
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2682 7936 2688 7948
rect 2643 7908 2688 7936
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7905 4399 7939
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4341 7899 4399 7905
rect 1535 7871 1593 7877
rect 1535 7837 1547 7871
rect 1581 7868 1593 7871
rect 1762 7868 1768 7880
rect 1581 7840 1768 7868
rect 1581 7837 1593 7840
rect 1535 7831 1593 7837
rect 1762 7828 1768 7840
rect 1820 7868 1826 7880
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 1820 7840 3433 7868
rect 1820 7828 1826 7840
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 4356 7868 4384 7899
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 7006 7936 7012 7948
rect 6919 7908 7012 7936
rect 7006 7896 7012 7908
rect 7064 7936 7070 7948
rect 8938 7936 8944 7948
rect 7064 7908 8944 7936
rect 7064 7896 7070 7908
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7936 9183 7939
rect 9398 7936 9404 7948
rect 9171 7908 9404 7936
rect 9171 7905 9183 7908
rect 9125 7899 9183 7905
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 9766 7936 9772 7948
rect 9539 7908 9772 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 4706 7868 4712 7880
rect 4356 7840 4712 7868
rect 3421 7831 3479 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 2038 7692 2044 7744
rect 2096 7732 2102 7744
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 2096 7704 2237 7732
rect 2096 7692 2102 7704
rect 2225 7701 2237 7704
rect 2271 7701 2283 7735
rect 5534 7732 5540 7744
rect 5495 7704 5540 7732
rect 2225 7695 2283 7701
rect 5534 7692 5540 7704
rect 5592 7732 5598 7744
rect 5736 7732 5764 7831
rect 6638 7800 6644 7812
rect 6599 7772 6644 7800
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 7944 7800 7972 7831
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8168 7840 8401 7868
rect 8168 7828 8174 7840
rect 8389 7837 8401 7840
rect 8435 7868 8447 7871
rect 9030 7868 9036 7880
rect 8435 7840 9036 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9508 7800 9536 7899
rect 9766 7896 9772 7908
rect 9824 7936 9830 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9824 7908 9873 7936
rect 9824 7896 9830 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10244 7877 10272 7976
rect 10597 7973 10609 8007
rect 10643 8004 10655 8007
rect 11330 8004 11336 8016
rect 10643 7976 11336 8004
rect 10643 7973 10655 7976
rect 10597 7967 10655 7973
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 12066 8004 12072 8016
rect 11480 7976 12072 8004
rect 11480 7964 11486 7976
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 13081 8007 13139 8013
rect 13081 7973 13093 8007
rect 13127 8004 13139 8007
rect 13354 8004 13360 8016
rect 13127 7976 13360 8004
rect 13127 7973 13139 7976
rect 13081 7967 13139 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 13630 8004 13636 8016
rect 13591 7976 13636 8004
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 15378 8004 15384 8016
rect 15339 7976 15384 8004
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 15473 8007 15531 8013
rect 15473 7973 15485 8007
rect 15519 8004 15531 8007
rect 15562 8004 15568 8016
rect 15519 7976 15568 8004
rect 15519 7973 15531 7976
rect 15473 7967 15531 7973
rect 15562 7964 15568 7976
rect 15620 7964 15626 8016
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7936 10839 7939
rect 10965 7939 11023 7945
rect 10965 7936 10977 7939
rect 10827 7908 10977 7936
rect 10827 7905 10839 7908
rect 10781 7899 10839 7905
rect 10965 7905 10977 7908
rect 11011 7936 11023 7939
rect 11146 7936 11152 7948
rect 11011 7908 11152 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11146 7896 11152 7908
rect 11204 7936 11210 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 11204 7908 11253 7936
rect 11204 7896 11210 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 11606 7936 11612 7948
rect 11567 7908 11612 7936
rect 11241 7899 11299 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 10008 7871 10066 7877
rect 10008 7837 10020 7871
rect 10054 7868 10066 7871
rect 10229 7871 10287 7877
rect 10054 7840 10180 7868
rect 10054 7837 10066 7840
rect 10008 7831 10066 7837
rect 7944 7772 9536 7800
rect 10152 7800 10180 7840
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 11882 7868 11888 7880
rect 10275 7840 11888 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13262 7868 13268 7880
rect 13035 7840 13268 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 11054 7800 11060 7812
rect 10152 7772 11060 7800
rect 11054 7760 11060 7772
rect 11112 7800 11118 7812
rect 11992 7800 12020 7831
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13648 7868 13676 7964
rect 17954 7936 17960 7948
rect 17915 7908 17960 7936
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 19004 7939 19062 7945
rect 19004 7936 19016 7939
rect 18748 7908 19016 7936
rect 18748 7896 18754 7908
rect 19004 7905 19016 7908
rect 19050 7905 19062 7939
rect 19004 7899 19062 7905
rect 23636 7939 23694 7945
rect 23636 7905 23648 7939
rect 23682 7936 23694 7939
rect 23842 7936 23848 7948
rect 23682 7908 23848 7936
rect 23682 7905 23694 7908
rect 23636 7899 23694 7905
rect 23842 7896 23848 7908
rect 23900 7896 23906 7948
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 13648 7840 15025 7868
rect 15013 7837 15025 7840
rect 15059 7837 15071 7871
rect 16022 7868 16028 7880
rect 15983 7840 16028 7868
rect 15013 7831 15071 7837
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 18138 7868 18144 7880
rect 18099 7840 18144 7868
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 11112 7772 15884 7800
rect 11112 7760 11118 7772
rect 7558 7732 7564 7744
rect 5592 7704 5764 7732
rect 7519 7704 7564 7732
rect 5592 7692 5598 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 8159 7735 8217 7741
rect 8159 7732 8171 7735
rect 7984 7704 8171 7732
rect 7984 7692 7990 7704
rect 8159 7701 8171 7704
rect 8205 7701 8217 7735
rect 8159 7695 8217 7701
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8662 7732 8668 7744
rect 8343 7704 8668 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10226 7732 10232 7744
rect 10183 7704 10232 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10226 7692 10232 7704
rect 10284 7732 10290 7744
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10284 7704 10793 7732
rect 10284 7692 10290 7704
rect 10781 7701 10793 7704
rect 10827 7701 10839 7735
rect 10781 7695 10839 7701
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 13722 7732 13728 7744
rect 11848 7704 13728 7732
rect 11848 7692 11854 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15856 7732 15884 7772
rect 16942 7732 16948 7744
rect 15856 7704 16948 7732
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 23707 7735 23765 7741
rect 23707 7701 23719 7735
rect 23753 7732 23765 7735
rect 24210 7732 24216 7744
rect 23753 7704 24216 7732
rect 23753 7701 23765 7704
rect 23707 7695 23765 7701
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2958 7528 2964 7540
rect 2919 7500 2964 7528
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4706 7528 4712 7540
rect 4126 7500 4712 7528
rect 2682 7460 2688 7472
rect 2595 7432 2688 7460
rect 2682 7420 2688 7432
rect 2740 7460 2746 7472
rect 4126 7460 4154 7500
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5077 7531 5135 7537
rect 5077 7497 5089 7531
rect 5123 7528 5135 7531
rect 5442 7528 5448 7540
rect 5123 7500 5448 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7558 7528 7564 7540
rect 6687 7500 7564 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 10118 7531 10176 7537
rect 7975 7500 8708 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8680 7472 8708 7500
rect 10118 7497 10130 7531
rect 10164 7528 10176 7531
rect 10778 7528 10784 7540
rect 10164 7500 10784 7528
rect 10164 7497 10176 7500
rect 10118 7491 10176 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11940 7500 12173 7528
rect 11940 7488 11946 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 13354 7528 13360 7540
rect 12759 7500 13360 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15562 7528 15568 7540
rect 15335 7500 15568 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 5166 7460 5172 7472
rect 2740 7432 4154 7460
rect 4264 7432 5172 7460
rect 2740 7420 2746 7432
rect 1578 7392 1584 7404
rect 1539 7364 1584 7392
rect 1578 7352 1584 7364
rect 1636 7352 1642 7404
rect 4264 7392 4292 7432
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 5316 7432 5948 7460
rect 5316 7420 5322 7432
rect 3620 7364 4292 7392
rect 4341 7395 4399 7401
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 3620 7333 3648 7364
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 5534 7392 5540 7404
rect 4387 7364 5540 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5920 7401 5948 7432
rect 8662 7420 8668 7472
rect 8720 7460 8726 7472
rect 9217 7463 9275 7469
rect 9217 7460 9229 7463
rect 8720 7432 9229 7460
rect 8720 7420 8726 7432
rect 9217 7429 9229 7432
rect 9263 7429 9275 7463
rect 10226 7460 10232 7472
rect 10187 7432 10232 7460
rect 9217 7423 9275 7429
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 11296 7432 13645 7460
rect 11296 7420 11302 7432
rect 13633 7429 13645 7432
rect 13679 7460 13691 7463
rect 13679 7432 14412 7460
rect 13679 7429 13691 7432
rect 13633 7423 13691 7429
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 5951 7364 7205 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8343 7364 8769 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8757 7361 8769 7364
rect 8803 7392 8815 7395
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 8803 7364 10333 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 3436 7296 3617 7324
rect 3436 7200 3464 7296
rect 3605 7293 3617 7296
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7324 4215 7327
rect 4246 7324 4252 7336
rect 4203 7296 4252 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 4246 7284 4252 7296
rect 4304 7324 4310 7336
rect 8536 7327 8594 7333
rect 4304 7296 5120 7324
rect 4304 7284 4310 7296
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 5092 7188 5120 7296
rect 8536 7293 8548 7327
rect 8582 7324 8594 7327
rect 8662 7324 8668 7336
rect 8582 7296 8668 7324
rect 8582 7293 8594 7296
rect 8536 7287 8594 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9824 7296 9965 7324
rect 9824 7284 9830 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 5258 7256 5264 7268
rect 5219 7228 5264 7256
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 5442 7256 5448 7268
rect 5399 7228 5448 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 6917 7259 6975 7265
rect 6917 7225 6929 7259
rect 6963 7225 6975 7259
rect 6917 7219 6975 7225
rect 5994 7188 6000 7200
rect 5092 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 6932 7188 6960 7219
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 7064 7228 7109 7256
rect 7064 7216 7070 7228
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 8352 7228 8401 7256
rect 8352 7216 8358 7228
rect 8389 7225 8401 7228
rect 8435 7225 8447 7259
rect 8389 7219 8447 7225
rect 10060 7200 10088 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 14384 7392 14412 7432
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 16761 7463 16819 7469
rect 16761 7460 16773 7463
rect 15436 7432 16773 7460
rect 15436 7420 15442 7432
rect 16761 7429 16773 7432
rect 16807 7429 16819 7463
rect 16761 7423 16819 7429
rect 13228 7364 13860 7392
rect 13228 7352 13234 7364
rect 10134 7284 10140 7336
rect 10192 7324 10198 7336
rect 13832 7333 13860 7364
rect 14384 7364 15976 7392
rect 14384 7333 14412 7364
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 10192 7296 12817 7324
rect 10192 7284 10198 7296
rect 12805 7293 12817 7296
rect 12851 7324 12863 7327
rect 13817 7327 13875 7333
rect 12851 7296 13400 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 10686 7256 10692 7268
rect 10647 7228 10692 7256
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11517 7259 11575 7265
rect 11517 7225 11529 7259
rect 11563 7256 11575 7259
rect 11606 7256 11612 7268
rect 11563 7228 11612 7256
rect 11563 7225 11575 7228
rect 11517 7219 11575 7225
rect 11606 7216 11612 7228
rect 11664 7256 11670 7268
rect 12526 7256 12532 7268
rect 11664 7228 12532 7256
rect 11664 7216 11670 7228
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 9030 7188 9036 7200
rect 6880 7160 6960 7188
rect 8991 7160 9036 7188
rect 6880 7148 6886 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7188 9275 7191
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 9263 7160 9505 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9493 7157 9505 7160
rect 9539 7188 9551 7191
rect 9674 7188 9680 7200
rect 9539 7160 9680 7188
rect 9539 7157 9551 7160
rect 9493 7151 9551 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10042 7188 10048 7200
rect 9907 7160 10048 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 11885 7191 11943 7197
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 12066 7188 12072 7200
rect 11931 7160 12072 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 13170 7188 13176 7200
rect 13035 7160 13176 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13372 7197 13400 7296
rect 13817 7293 13829 7327
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 15948 7333 15976 7364
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 14884 7296 15393 7324
rect 14884 7284 14890 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7324 15991 7327
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 15979 7296 16405 7324
rect 15979 7293 15991 7296
rect 15933 7287 15991 7293
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16393 7287 16451 7293
rect 16942 7284 16948 7296
rect 17000 7324 17006 7336
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17000 7296 17417 7324
rect 17000 7284 17006 7296
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 18141 7327 18199 7333
rect 18141 7293 18153 7327
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 14553 7259 14611 7265
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 16114 7256 16120 7268
rect 14599 7228 15332 7256
rect 16075 7228 16120 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 15304 7200 15332 7228
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 18046 7256 18052 7268
rect 18007 7228 18052 7256
rect 18046 7216 18052 7228
rect 18104 7216 18110 7268
rect 13357 7191 13415 7197
rect 13357 7157 13369 7191
rect 13403 7188 13415 7191
rect 14090 7188 14096 7200
rect 13403 7160 14096 7188
rect 13403 7157 13415 7160
rect 13357 7151 13415 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14826 7188 14832 7200
rect 14787 7160 14832 7188
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 15286 7148 15292 7200
rect 15344 7148 15350 7200
rect 17126 7188 17132 7200
rect 17087 7160 17132 7188
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 17862 7188 17868 7200
rect 17823 7160 17868 7188
rect 17862 7148 17868 7160
rect 17920 7188 17926 7200
rect 18156 7188 18184 7287
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 19648 7327 19706 7333
rect 19648 7324 19660 7327
rect 18288 7296 19660 7324
rect 18288 7284 18294 7296
rect 19648 7293 19660 7296
rect 19694 7324 19706 7327
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19694 7296 20085 7324
rect 19694 7293 19706 7296
rect 19648 7287 19706 7293
rect 20073 7293 20085 7296
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 20676 7327 20734 7333
rect 20676 7293 20688 7327
rect 20722 7324 20734 7327
rect 20722 7293 20735 7324
rect 20676 7287 20735 7293
rect 17920 7160 18184 7188
rect 17920 7148 17926 7160
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18748 7160 19073 7188
rect 18748 7148 18754 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19150 7148 19156 7200
rect 19208 7188 19214 7200
rect 19751 7191 19809 7197
rect 19751 7188 19763 7191
rect 19208 7160 19763 7188
rect 19208 7148 19214 7160
rect 19751 7157 19763 7160
rect 19797 7157 19809 7191
rect 20707 7188 20735 7287
rect 20898 7284 20904 7336
rect 20956 7324 20962 7336
rect 21704 7327 21762 7333
rect 21704 7324 21716 7327
rect 20956 7296 21716 7324
rect 20956 7284 20962 7296
rect 21704 7293 21716 7296
rect 21750 7324 21762 7327
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 21750 7296 22109 7324
rect 21750 7293 21762 7296
rect 21704 7287 21762 7293
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 20763 7259 20821 7265
rect 20763 7225 20775 7259
rect 20809 7256 20821 7259
rect 20809 7228 21680 7256
rect 20809 7225 20821 7228
rect 20763 7219 20821 7225
rect 21652 7200 21680 7228
rect 21082 7188 21088 7200
rect 20707 7160 21088 7188
rect 19751 7151 19809 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 21634 7148 21640 7200
rect 21692 7148 21698 7200
rect 21775 7191 21833 7197
rect 21775 7157 21787 7191
rect 21821 7188 21833 7191
rect 22002 7188 22008 7200
rect 21821 7160 22008 7188
rect 21821 7157 21833 7160
rect 21775 7151 21833 7157
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 23842 7188 23848 7200
rect 23803 7160 23848 7188
rect 23842 7148 23848 7160
rect 23900 7148 23906 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 2148 6956 3065 6984
rect 2038 6916 2044 6928
rect 1999 6888 2044 6916
rect 2038 6876 2044 6888
rect 2096 6876 2102 6928
rect 2148 6925 2176 6956
rect 3053 6953 3065 6956
rect 3099 6984 3111 6987
rect 5534 6984 5540 6996
rect 3099 6956 5540 6984
rect 3099 6953 3111 6956
rect 3053 6947 3111 6953
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 6365 6987 6423 6993
rect 6365 6953 6377 6987
rect 6411 6984 6423 6987
rect 7006 6984 7012 6996
rect 6411 6956 7012 6984
rect 6411 6953 6423 6956
rect 6365 6947 6423 6953
rect 7006 6944 7012 6956
rect 7064 6944 7070 6996
rect 7561 6987 7619 6993
rect 7561 6953 7573 6987
rect 7607 6984 7619 6987
rect 8110 6984 8116 6996
rect 7607 6956 8116 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9214 6984 9220 6996
rect 9171 6956 9220 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9364 6956 9413 6984
rect 9364 6944 9370 6956
rect 9401 6953 9413 6956
rect 9447 6984 9459 6987
rect 10321 6987 10379 6993
rect 9447 6956 10272 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 2133 6919 2191 6925
rect 2133 6885 2145 6919
rect 2179 6885 2191 6919
rect 2133 6879 2191 6885
rect 5807 6919 5865 6925
rect 5807 6885 5819 6919
rect 5853 6916 5865 6919
rect 6178 6916 6184 6928
rect 5853 6888 6184 6916
rect 5853 6885 5865 6888
rect 5807 6879 5865 6885
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 8021 6919 8079 6925
rect 8021 6916 8033 6919
rect 7432 6888 8033 6916
rect 7432 6876 7438 6888
rect 8021 6885 8033 6888
rect 8067 6916 8079 6919
rect 9324 6916 9352 6944
rect 9692 6925 9720 6956
rect 8067 6888 9352 6916
rect 9677 6919 9735 6925
rect 8067 6885 8079 6888
rect 8021 6879 8079 6885
rect 9677 6885 9689 6919
rect 9723 6885 9735 6919
rect 10244 6916 10272 6956
rect 10321 6953 10333 6987
rect 10367 6984 10379 6987
rect 12710 6984 12716 6996
rect 10367 6956 12572 6984
rect 12671 6956 12716 6984
rect 10367 6953 10379 6956
rect 10321 6947 10379 6953
rect 11146 6916 11152 6928
rect 10244 6888 11152 6916
rect 9677 6879 9735 6885
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 12544 6916 12572 6956
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 13081 6987 13139 6993
rect 13081 6953 13093 6987
rect 13127 6984 13139 6987
rect 13262 6984 13268 6996
rect 13127 6956 13268 6984
rect 13127 6953 13139 6956
rect 13081 6947 13139 6953
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 16206 6984 16212 6996
rect 16167 6956 16212 6984
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17954 6984 17960 6996
rect 17915 6956 17960 6984
rect 17954 6944 17960 6956
rect 18012 6984 18018 6996
rect 18233 6987 18291 6993
rect 18233 6984 18245 6987
rect 18012 6956 18245 6984
rect 18012 6944 18018 6956
rect 18233 6953 18245 6956
rect 18279 6953 18291 6987
rect 18233 6947 18291 6953
rect 13446 6916 13452 6928
rect 12544 6888 13452 6916
rect 13446 6876 13452 6888
rect 13504 6916 13510 6928
rect 13504 6888 14136 6916
rect 13504 6876 13510 6888
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 3050 6848 3056 6860
rect 2731 6820 3056 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4100 6851 4158 6857
rect 4100 6848 4112 6851
rect 3844 6820 4112 6848
rect 3844 6808 3850 6820
rect 4100 6817 4112 6820
rect 4146 6817 4158 6851
rect 4100 6811 4158 6817
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7558 6848 7564 6860
rect 7239 6820 7564 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7558 6808 7564 6820
rect 7616 6848 7622 6860
rect 8168 6851 8226 6857
rect 8168 6848 8180 6851
rect 7616 6820 8180 6848
rect 7616 6808 7622 6820
rect 8168 6817 8180 6820
rect 8214 6848 8226 6851
rect 8662 6848 8668 6860
rect 8214 6820 8668 6848
rect 8214 6817 8226 6820
rect 8168 6811 8226 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 9916 6820 11069 6848
rect 9916 6808 9922 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11238 6848 11244 6860
rect 11199 6820 11244 6848
rect 11057 6811 11115 6817
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 11440 6820 12357 6848
rect 4246 6780 4252 6792
rect 4126 6752 4252 6780
rect 3697 6715 3755 6721
rect 3697 6681 3709 6715
rect 3743 6712 3755 6715
rect 4126 6712 4154 6752
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8570 6780 8576 6792
rect 8435 6752 8576 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 10042 6780 10048 6792
rect 9646 6752 9867 6780
rect 10003 6752 10048 6780
rect 4614 6712 4620 6724
rect 3743 6684 4154 6712
rect 4527 6684 4620 6712
rect 3743 6681 3755 6684
rect 3697 6675 3755 6681
rect 4614 6672 4620 6684
rect 4672 6712 4678 6724
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 4672 6684 8493 6712
rect 4672 6672 4678 6684
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 9646 6712 9674 6752
rect 8720 6684 9674 6712
rect 9839 6721 9867 6752
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11440 6780 11468 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 14108 6857 14136 6888
rect 14274 6876 14280 6928
rect 14332 6916 14338 6928
rect 15610 6919 15668 6925
rect 15610 6916 15622 6919
rect 14332 6888 15622 6916
rect 14332 6876 14338 6888
rect 15610 6885 15622 6888
rect 15656 6885 15668 6919
rect 15610 6879 15668 6885
rect 18138 6876 18144 6928
rect 18196 6916 18202 6928
rect 18969 6919 19027 6925
rect 18969 6916 18981 6919
rect 18196 6888 18981 6916
rect 18196 6876 18202 6888
rect 18969 6885 18981 6888
rect 19015 6916 19027 6919
rect 19058 6916 19064 6928
rect 19015 6888 19064 6916
rect 19015 6885 19027 6888
rect 18969 6879 19027 6885
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13228 6820 13645 6848
rect 13228 6808 13234 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 14093 6851 14151 6857
rect 14093 6817 14105 6851
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 16114 6808 16120 6860
rect 16172 6848 16178 6860
rect 16758 6848 16764 6860
rect 16172 6820 16764 6848
rect 16172 6808 16178 6820
rect 16758 6808 16764 6820
rect 16816 6848 16822 6860
rect 17037 6851 17095 6857
rect 17037 6848 17049 6851
rect 16816 6820 17049 6848
rect 16816 6808 16822 6820
rect 17037 6817 17049 6820
rect 17083 6817 17095 6851
rect 20806 6848 20812 6860
rect 20767 6820 20812 6848
rect 17037 6811 17095 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 21818 6808 21824 6860
rect 21876 6848 21882 6860
rect 21948 6851 22006 6857
rect 21948 6848 21960 6851
rect 21876 6820 21960 6848
rect 21876 6808 21882 6820
rect 21948 6817 21960 6820
rect 21994 6817 22006 6851
rect 21948 6811 22006 6817
rect 24210 6808 24216 6860
rect 24268 6848 24274 6860
rect 24581 6851 24639 6857
rect 24581 6848 24593 6851
rect 24268 6820 24593 6848
rect 24268 6808 24274 6820
rect 24581 6817 24593 6820
rect 24627 6817 24639 6851
rect 24581 6811 24639 6817
rect 11606 6780 11612 6792
rect 10612 6752 11468 6780
rect 11519 6752 11612 6780
rect 9839 6715 9900 6721
rect 9839 6684 9854 6715
rect 8720 6672 8726 6684
rect 9842 6681 9854 6684
rect 9888 6712 9900 6715
rect 10612 6712 10640 6752
rect 11606 6740 11612 6752
rect 11664 6780 11670 6792
rect 11882 6780 11888 6792
rect 11664 6752 11888 6780
rect 11664 6740 11670 6752
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12250 6780 12256 6792
rect 12023 6752 12256 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 15286 6780 15292 6792
rect 15247 6752 15292 6780
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 17000 6752 18889 6780
rect 17000 6740 17006 6752
rect 18877 6749 18889 6752
rect 18923 6780 18935 6783
rect 19334 6780 19340 6792
rect 18923 6752 19340 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 21039 6783 21097 6789
rect 21039 6749 21051 6783
rect 21085 6780 21097 6783
rect 23842 6780 23848 6792
rect 21085 6752 23848 6780
rect 21085 6749 21097 6752
rect 21039 6743 21097 6749
rect 23842 6740 23848 6752
rect 23900 6740 23906 6792
rect 11379 6715 11437 6721
rect 11379 6712 11391 6715
rect 9888 6684 10640 6712
rect 10796 6684 11391 6712
rect 9888 6681 9900 6684
rect 9842 6675 9900 6681
rect 10796 6656 10824 6684
rect 11379 6681 11391 6684
rect 11425 6681 11437 6715
rect 11379 6675 11437 6681
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12400 6684 13124 6712
rect 12400 6672 12406 6684
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1452 6616 1593 6644
rect 1452 6604 1458 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 4203 6647 4261 6653
rect 4203 6613 4215 6647
rect 4249 6644 4261 6647
rect 4430 6644 4436 6656
rect 4249 6616 4436 6644
rect 4249 6613 4261 6616
rect 4203 6607 4261 6613
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 4890 6644 4896 6656
rect 4851 6616 4896 6644
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7926 6644 7932 6656
rect 7887 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8846 6644 8852 6656
rect 8343 6616 8852 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10134 6644 10140 6656
rect 9999 6616 10140 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10778 6644 10784 6656
rect 10739 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11514 6644 11520 6656
rect 11475 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 13096 6644 13124 6684
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 17126 6712 17132 6724
rect 13228 6684 17132 6712
rect 13228 6672 13234 6684
rect 17126 6672 17132 6684
rect 17184 6672 17190 6724
rect 18782 6672 18788 6724
rect 18840 6712 18846 6724
rect 19429 6715 19487 6721
rect 19429 6712 19441 6715
rect 18840 6684 19441 6712
rect 18840 6672 18846 6684
rect 19429 6681 19441 6684
rect 19475 6712 19487 6715
rect 24118 6712 24124 6724
rect 19475 6684 24124 6712
rect 19475 6681 19487 6684
rect 19429 6675 19487 6681
rect 24118 6672 24124 6684
rect 24176 6672 24182 6724
rect 19150 6644 19156 6656
rect 13096 6616 19156 6644
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 22051 6647 22109 6653
rect 22051 6644 22063 6647
rect 19300 6616 22063 6644
rect 19300 6604 19306 6616
rect 22051 6613 22063 6616
rect 22097 6613 22109 6647
rect 22051 6607 22109 6613
rect 24765 6647 24823 6653
rect 24765 6613 24777 6647
rect 24811 6644 24823 6647
rect 26786 6644 26792 6656
rect 24811 6616 26792 6644
rect 24811 6613 24823 6616
rect 24765 6607 24823 6613
rect 26786 6604 26792 6616
rect 26844 6604 26850 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2455 6412 2697 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2685 6409 2697 6412
rect 2731 6440 2743 6443
rect 2866 6440 2872 6452
rect 2731 6412 2872 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 3844 6412 4353 6440
rect 3844 6400 3850 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5592 6412 5825 6440
rect 5592 6400 5598 6412
rect 5813 6409 5825 6412
rect 5859 6440 5871 6443
rect 7098 6440 7104 6452
rect 5859 6412 7104 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7374 6440 7380 6452
rect 7335 6412 7380 6440
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8462 6443 8520 6449
rect 8462 6440 8474 6443
rect 7984 6412 8474 6440
rect 7984 6400 7990 6412
rect 8462 6409 8474 6412
rect 8508 6440 8520 6443
rect 9490 6440 9496 6452
rect 8508 6412 9496 6440
rect 8508 6409 8520 6412
rect 8462 6403 8520 6409
rect 9490 6400 9496 6412
rect 9548 6440 9554 6452
rect 10026 6443 10084 6449
rect 10026 6440 10038 6443
rect 9548 6412 10038 6440
rect 9548 6400 9554 6412
rect 10026 6409 10038 6412
rect 10072 6440 10084 6443
rect 10778 6440 10784 6452
rect 10072 6412 10784 6440
rect 10072 6409 10084 6412
rect 10026 6403 10084 6409
rect 10778 6400 10784 6412
rect 10836 6440 10842 6452
rect 11330 6440 11336 6452
rect 10836 6412 11336 6440
rect 10836 6400 10842 6412
rect 11330 6400 11336 6412
rect 11388 6440 11394 6452
rect 11701 6443 11759 6449
rect 11701 6440 11713 6443
rect 11388 6412 11713 6440
rect 11388 6400 11394 6412
rect 11701 6409 11713 6412
rect 11747 6440 11759 6443
rect 13170 6440 13176 6452
rect 11747 6412 13176 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 13320 6412 13461 6440
rect 13320 6400 13326 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 14826 6440 14832 6452
rect 14231 6412 14832 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15344 6412 16221 6440
rect 15344 6400 15350 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16758 6440 16764 6452
rect 16719 6412 16764 6440
rect 16209 6403 16267 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 17954 6440 17960 6452
rect 17911 6412 17960 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19392 6412 19441 6440
rect 19392 6400 19398 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 21818 6400 21824 6452
rect 21876 6440 21882 6452
rect 22005 6443 22063 6449
rect 22005 6440 22017 6443
rect 21876 6412 22017 6440
rect 21876 6400 21882 6412
rect 22005 6409 22017 6412
rect 22051 6409 22063 6443
rect 22005 6403 22063 6409
rect 24210 6400 24216 6452
rect 24268 6440 24274 6452
rect 24581 6443 24639 6449
rect 24581 6440 24593 6443
rect 24268 6412 24593 6440
rect 24268 6400 24274 6412
rect 24581 6409 24593 6412
rect 24627 6409 24639 6443
rect 24581 6403 24639 6409
rect 2225 6375 2283 6381
rect 2225 6341 2237 6375
rect 2271 6372 2283 6375
rect 3050 6372 3056 6384
rect 2271 6344 3056 6372
rect 2271 6341 2283 6344
rect 2225 6335 2283 6341
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6372 7803 6375
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 7791 6344 8585 6372
rect 7791 6341 7803 6344
rect 7745 6335 7803 6341
rect 8573 6341 8585 6344
rect 8619 6372 8631 6375
rect 9674 6372 9680 6384
rect 8619 6344 9680 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 9674 6332 9680 6344
rect 9732 6372 9738 6384
rect 10134 6372 10140 6384
rect 9732 6344 10140 6372
rect 9732 6332 9738 6344
rect 10134 6332 10140 6344
rect 10192 6372 10198 6384
rect 10192 6344 11008 6372
rect 10192 6332 10198 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 2498 6304 2504 6316
rect 1719 6276 2504 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3234 6304 3240 6316
rect 3191 6276 3240 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3234 6264 3240 6276
rect 3292 6304 3298 6316
rect 4062 6304 4068 6316
rect 3292 6276 4068 6304
rect 3292 6264 3298 6276
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 8662 6304 8668 6316
rect 8575 6276 8668 6304
rect 8662 6264 8668 6276
rect 8720 6304 8726 6316
rect 10229 6307 10287 6313
rect 8720 6276 9444 6304
rect 8720 6264 8726 6276
rect 4890 6236 4896 6248
rect 4851 6208 4896 6236
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 8570 6236 8576 6248
rect 8159 6208 8576 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9416 6245 9444 6276
rect 10229 6273 10241 6307
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6236 9459 6239
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9447 6208 9781 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 9769 6205 9781 6208
rect 9815 6236 9827 6239
rect 10042 6236 10048 6248
rect 9815 6208 10048 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10042 6196 10048 6208
rect 10100 6236 10106 6248
rect 10244 6236 10272 6267
rect 10100 6208 10272 6236
rect 10100 6196 10106 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2409 6171 2467 6177
rect 2409 6168 2421 6171
rect 1811 6140 2421 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2409 6137 2421 6140
rect 2455 6137 2467 6171
rect 2409 6131 2467 6137
rect 3053 6171 3111 6177
rect 3053 6137 3065 6171
rect 3099 6168 3111 6171
rect 3507 6171 3565 6177
rect 3507 6168 3519 6171
rect 3099 6140 3519 6168
rect 3099 6137 3111 6140
rect 3053 6131 3111 6137
rect 3507 6137 3519 6140
rect 3553 6168 3565 6171
rect 5255 6171 5313 6177
rect 3553 6140 4844 6168
rect 3553 6137 3565 6140
rect 3507 6131 3565 6137
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 4816 6109 4844 6140
rect 5255 6137 5267 6171
rect 5301 6137 5313 6171
rect 5255 6131 5313 6137
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3200 6072 4077 6100
rect 3200 6060 3206 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5270 6100 5298 6131
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 6457 6171 6515 6177
rect 6457 6168 6469 6171
rect 5500 6140 6469 6168
rect 5500 6128 5506 6140
rect 6457 6137 6469 6140
rect 6503 6137 6515 6171
rect 6457 6131 6515 6137
rect 8297 6171 8355 6177
rect 8297 6137 8309 6171
rect 8343 6168 8355 6171
rect 9214 6168 9220 6180
rect 8343 6140 9220 6168
rect 8343 6137 8355 6140
rect 8297 6131 8355 6137
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 9858 6168 9864 6180
rect 9819 6140 9864 6168
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 6178 6100 6184 6112
rect 4847 6072 6184 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8168 6072 8953 6100
rect 8168 6060 8174 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 8941 6063 8999 6069
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10980 6109 11008 6344
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 14734 6372 14740 6384
rect 12032 6344 14740 6372
rect 12032 6332 12038 6344
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 19242 6372 19248 6384
rect 15304 6344 19248 6372
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12710 6304 12716 6316
rect 12575 6276 12716 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13044 6276 13921 6304
rect 13044 6264 13050 6276
rect 13909 6273 13921 6276
rect 13955 6304 13967 6307
rect 14366 6304 14372 6316
rect 13955 6276 14372 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14016 6245 14044 6276
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15304 6313 15332 6344
rect 19242 6332 19248 6344
rect 19300 6332 19306 6384
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15160 6276 15301 6304
rect 15160 6264 15166 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 16942 6304 16948 6316
rect 16903 6276 16948 6304
rect 15289 6267 15347 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 18782 6304 18788 6316
rect 18743 6276 18788 6304
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19484 6276 21991 6304
rect 19484 6264 19490 6276
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13979 6208 14013 6236
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 14826 6236 14832 6248
rect 14240 6208 14832 6236
rect 14240 6196 14246 6208
rect 14826 6196 14832 6208
rect 14884 6236 14890 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 14884 6208 15025 6236
rect 14884 6196 14890 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 15013 6199 15071 6205
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 21244 6239 21302 6245
rect 21244 6205 21256 6239
rect 21290 6236 21302 6239
rect 21542 6236 21548 6248
rect 21290 6208 21548 6236
rect 21290 6205 21302 6208
rect 21244 6199 21302 6205
rect 21542 6196 21548 6208
rect 21600 6236 21606 6248
rect 21637 6239 21695 6245
rect 21637 6236 21649 6239
rect 21600 6208 21649 6236
rect 21600 6196 21606 6208
rect 21637 6205 21649 6208
rect 21683 6205 21695 6239
rect 21963 6236 21991 6276
rect 22224 6239 22282 6245
rect 22224 6236 22236 6239
rect 21963 6208 22236 6236
rect 21637 6199 21695 6205
rect 22224 6205 22236 6208
rect 22270 6236 22282 6239
rect 22649 6239 22707 6245
rect 22649 6236 22661 6239
rect 22270 6208 22661 6236
rect 22270 6205 22282 6208
rect 22224 6199 22282 6205
rect 22649 6205 22661 6208
rect 22695 6205 22707 6239
rect 22649 6199 22707 6205
rect 23728 6239 23786 6245
rect 23728 6205 23740 6239
rect 23774 6236 23786 6239
rect 24118 6236 24124 6248
rect 23774 6208 24124 6236
rect 23774 6205 23786 6208
rect 23728 6199 23786 6205
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 12618 6168 12624 6180
rect 12299 6140 12624 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 13170 6168 13176 6180
rect 13131 6140 13176 6168
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 14642 6168 14648 6180
rect 13786 6140 14648 6168
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 9824 6072 10517 6100
rect 9824 6060 9830 6072
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 10505 6063 10563 6069
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 11011 6072 11345 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11333 6069 11345 6072
rect 11379 6100 11391 6103
rect 11422 6100 11428 6112
rect 11379 6072 11428 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 13786 6100 13814 6140
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 14737 6171 14795 6177
rect 14737 6137 14749 6171
rect 14783 6168 14795 6171
rect 15381 6171 15439 6177
rect 14783 6140 15240 6168
rect 14783 6137 14795 6140
rect 14737 6131 14795 6137
rect 11940 6072 13814 6100
rect 15212 6100 15240 6140
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 15470 6168 15476 6180
rect 15427 6140 15476 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 15396 6100 15424 6131
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 15930 6168 15936 6180
rect 15891 6140 15936 6168
rect 15930 6128 15936 6140
rect 15988 6168 15994 6180
rect 18138 6168 18144 6180
rect 15988 6140 18144 6168
rect 15988 6128 15994 6140
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6137 18291 6171
rect 18233 6131 18291 6137
rect 15212 6072 15424 6100
rect 11940 6060 11946 6072
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 17402 6100 17408 6112
rect 16908 6072 17408 6100
rect 16908 6060 16914 6072
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17954 6060 17960 6112
rect 18012 6100 18018 6112
rect 18248 6100 18276 6131
rect 18966 6128 18972 6180
rect 19024 6168 19030 6180
rect 19613 6171 19671 6177
rect 19613 6168 19625 6171
rect 19024 6140 19625 6168
rect 19024 6128 19030 6140
rect 19613 6137 19625 6140
rect 19659 6137 19671 6171
rect 19613 6131 19671 6137
rect 21450 6128 21456 6180
rect 21508 6168 21514 6180
rect 22327 6171 22385 6177
rect 22327 6168 22339 6171
rect 21508 6140 22339 6168
rect 21508 6128 21514 6140
rect 22327 6137 22339 6140
rect 22373 6137 22385 6171
rect 22327 6131 22385 6137
rect 18012 6072 18276 6100
rect 18012 6060 18018 6072
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 20806 6100 20812 6112
rect 20496 6072 20812 6100
rect 20496 6060 20502 6072
rect 20806 6060 20812 6072
rect 20864 6100 20870 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20864 6072 20913 6100
rect 20864 6060 20870 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 20901 6063 20959 6069
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 21315 6103 21373 6109
rect 21315 6100 21327 6103
rect 21140 6072 21327 6100
rect 21140 6060 21146 6072
rect 21315 6069 21327 6072
rect 21361 6069 21373 6103
rect 21315 6063 21373 6069
rect 23799 6103 23857 6109
rect 23799 6069 23811 6103
rect 23845 6100 23857 6103
rect 23934 6100 23940 6112
rect 23845 6072 23940 6100
rect 23845 6069 23857 6072
rect 23799 6063 23857 6069
rect 23934 6060 23940 6072
rect 23992 6060 23998 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2498 5896 2504 5908
rect 2459 5868 2504 5896
rect 2498 5856 2504 5868
rect 2556 5896 2562 5908
rect 2774 5896 2780 5908
rect 2556 5868 2780 5896
rect 2556 5856 2562 5868
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 4430 5896 4436 5908
rect 2884 5868 4436 5896
rect 1670 5828 1676 5840
rect 1631 5800 1676 5828
rect 1670 5788 1676 5800
rect 1728 5788 1734 5840
rect 2038 5788 2044 5840
rect 2096 5828 2102 5840
rect 2225 5831 2283 5837
rect 2225 5828 2237 5831
rect 2096 5800 2237 5828
rect 2096 5788 2102 5800
rect 2225 5797 2237 5800
rect 2271 5797 2283 5831
rect 2225 5791 2283 5797
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2884 5692 2912 5868
rect 4430 5856 4436 5868
rect 4488 5896 4494 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4488 5868 4537 5896
rect 4488 5856 4494 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 5442 5896 5448 5908
rect 5403 5868 5448 5896
rect 4525 5859 4583 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6696 5868 7021 5896
rect 6696 5856 6702 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 8662 5896 8668 5908
rect 8435 5868 8668 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 10781 5899 10839 5905
rect 10781 5865 10793 5899
rect 10827 5896 10839 5899
rect 11422 5896 11428 5908
rect 10827 5868 11428 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 11606 5896 11612 5908
rect 11567 5868 11612 5896
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 13446 5896 13452 5908
rect 13407 5868 13452 5896
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 15102 5896 15108 5908
rect 15063 5868 15108 5896
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16206 5896 16212 5908
rect 15887 5868 16212 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17405 5899 17463 5905
rect 17405 5865 17417 5899
rect 17451 5865 17463 5899
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 17405 5859 17463 5865
rect 3234 5828 3240 5840
rect 3195 5800 3240 5828
rect 3234 5788 3240 5800
rect 3292 5788 3298 5840
rect 5994 5828 6000 5840
rect 5907 5800 6000 5828
rect 4154 5769 4160 5772
rect 4132 5763 4160 5769
rect 4132 5729 4144 5763
rect 4132 5723 4160 5729
rect 4154 5720 4160 5723
rect 4212 5720 4218 5772
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 5350 5760 5356 5772
rect 4764 5732 5356 5760
rect 4764 5720 4770 5732
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5920 5769 5948 5800
rect 5994 5788 6000 5800
rect 6052 5828 6058 5840
rect 9030 5828 9036 5840
rect 6052 5800 9036 5828
rect 6052 5788 6058 5800
rect 9030 5788 9036 5800
rect 9088 5788 9094 5840
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 9677 5831 9735 5837
rect 9677 5828 9689 5831
rect 9272 5800 9689 5828
rect 9272 5788 9278 5800
rect 9677 5797 9689 5800
rect 9723 5828 9735 5831
rect 11238 5828 11244 5840
rect 9723 5800 11244 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 11238 5788 11244 5800
rect 11296 5788 11302 5840
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 12114 5831 12172 5837
rect 12114 5828 12126 5831
rect 12032 5800 12126 5828
rect 12032 5788 12038 5800
rect 12114 5797 12126 5800
rect 12160 5797 12172 5831
rect 12114 5791 12172 5797
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 17420 5828 17448 5859
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 19705 5899 19763 5905
rect 19705 5865 19717 5899
rect 19751 5896 19763 5899
rect 19978 5896 19984 5908
rect 19751 5868 19984 5896
rect 19751 5865 19763 5868
rect 19705 5859 19763 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 17862 5828 17868 5840
rect 13228 5800 16712 5828
rect 17420 5800 17868 5828
rect 13228 5788 13234 5800
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 5905 5723 5963 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7466 5760 7472 5772
rect 7427 5732 7472 5760
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 11793 5763 11851 5769
rect 11793 5760 11805 5763
rect 11756 5732 11805 5760
rect 11756 5720 11762 5732
rect 11793 5729 11805 5732
rect 11839 5729 11851 5763
rect 11793 5723 11851 5729
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12584 5732 13093 5760
rect 12584 5720 12590 5732
rect 13081 5729 13093 5732
rect 13127 5760 13139 5763
rect 13354 5760 13360 5772
rect 13127 5732 13360 5760
rect 13127 5729 13139 5732
rect 13081 5723 13139 5729
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 13630 5760 13636 5772
rect 13591 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 14093 5723 14151 5729
rect 1627 5664 2912 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2958 5652 2964 5704
rect 3016 5692 3022 5704
rect 6822 5692 6828 5704
rect 3016 5664 6828 5692
rect 3016 5652 3022 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 8478 5692 8484 5704
rect 8439 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5692 9091 5695
rect 9508 5692 9536 5720
rect 9824 5695 9882 5701
rect 9824 5692 9836 5695
rect 9079 5664 9836 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9824 5661 9836 5664
rect 9870 5661 9882 5695
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 9824 5655 9882 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 14108 5692 14136 5723
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 14366 5692 14372 5704
rect 13504 5664 14136 5692
rect 14327 5664 14372 5692
rect 13504 5652 13510 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 16482 5692 16488 5704
rect 14936 5664 16488 5692
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 3513 5627 3571 5633
rect 3513 5624 3525 5627
rect 1912 5596 3525 5624
rect 1912 5584 1918 5596
rect 3513 5593 3525 5596
rect 3559 5624 3571 5627
rect 4203 5627 4261 5633
rect 4203 5624 4215 5627
rect 3559 5596 4215 5624
rect 3559 5593 3571 5596
rect 3513 5587 3571 5593
rect 4203 5593 4215 5596
rect 4249 5593 4261 5627
rect 4203 5587 4261 5593
rect 12618 5584 12624 5636
rect 12676 5624 12682 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12676 5596 12725 5624
rect 12676 5584 12682 5596
rect 12713 5593 12725 5596
rect 12759 5624 12771 5627
rect 13998 5624 14004 5636
rect 12759 5596 14004 5624
rect 12759 5593 12771 5596
rect 12713 5587 12771 5593
rect 13998 5584 14004 5596
rect 14056 5584 14062 5636
rect 5258 5556 5264 5568
rect 5219 5528 5264 5556
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5556 8079 5559
rect 8846 5556 8852 5568
rect 8067 5528 8852 5556
rect 8067 5525 8079 5528
rect 8021 5519 8079 5525
rect 8846 5516 8852 5528
rect 8904 5556 8910 5568
rect 9953 5559 10011 5565
rect 9953 5556 9965 5559
rect 8904 5528 9965 5556
rect 8904 5516 8910 5528
rect 9953 5525 9965 5528
rect 9999 5525 10011 5559
rect 10134 5556 10140 5568
rect 10095 5528 10140 5556
rect 9953 5519 10011 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14936 5556 14964 5664
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 16684 5692 16712 5800
rect 17862 5788 17868 5800
rect 17920 5828 17926 5840
rect 18417 5831 18475 5837
rect 18417 5828 18429 5831
rect 17920 5800 18429 5828
rect 17920 5788 17926 5800
rect 18417 5797 18429 5800
rect 18463 5828 18475 5831
rect 19058 5828 19064 5840
rect 18463 5800 19064 5828
rect 18463 5797 18475 5800
rect 18417 5791 18475 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 19518 5788 19524 5840
rect 19576 5828 19582 5840
rect 23615 5831 23673 5837
rect 23615 5828 23627 5831
rect 19576 5800 23627 5828
rect 19576 5788 19582 5800
rect 23615 5797 23627 5800
rect 23661 5797 23673 5831
rect 23615 5791 23673 5797
rect 18969 5763 19027 5769
rect 18969 5729 18981 5763
rect 19015 5760 19027 5763
rect 19150 5760 19156 5772
rect 19015 5732 19156 5760
rect 19015 5729 19027 5732
rect 18969 5723 19027 5729
rect 19150 5720 19156 5732
rect 19208 5760 19214 5772
rect 20898 5760 20904 5772
rect 19208 5732 20904 5760
rect 19208 5720 19214 5732
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 22462 5760 22468 5772
rect 21048 5732 21093 5760
rect 22423 5732 22468 5760
rect 21048 5720 21054 5732
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 23290 5720 23296 5772
rect 23348 5760 23354 5772
rect 23512 5763 23570 5769
rect 23512 5760 23524 5763
rect 23348 5732 23524 5760
rect 23348 5720 23354 5732
rect 23512 5729 23524 5732
rect 23558 5729 23570 5763
rect 23512 5723 23570 5729
rect 18325 5695 18383 5701
rect 18325 5692 18337 5695
rect 16684 5664 18337 5692
rect 18325 5661 18337 5664
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18340 5624 18368 5655
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 19797 5695 19855 5701
rect 19797 5692 19809 5695
rect 18472 5664 19809 5692
rect 18472 5652 18478 5664
rect 19797 5661 19809 5664
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 18506 5624 18512 5636
rect 18340 5596 18512 5624
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 15470 5556 15476 5568
rect 13596 5528 14964 5556
rect 15431 5528 15476 5556
rect 13596 5516 13602 5528
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 16356 5528 21189 5556
rect 16356 5516 16362 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 22603 5559 22661 5565
rect 22603 5525 22615 5559
rect 22649 5556 22661 5559
rect 23382 5556 23388 5568
rect 22649 5528 23388 5556
rect 22649 5525 22661 5528
rect 22603 5519 22661 5525
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 7466 5352 7472 5364
rect 5592 5324 7472 5352
rect 5592 5312 5598 5324
rect 7466 5312 7472 5324
rect 7524 5352 7530 5364
rect 7929 5355 7987 5361
rect 7929 5352 7941 5355
rect 7524 5324 7941 5352
rect 7524 5312 7530 5324
rect 7929 5321 7941 5324
rect 7975 5352 7987 5355
rect 9766 5352 9772 5364
rect 7975 5324 9772 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10042 5352 10048 5364
rect 9907 5324 10048 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10042 5312 10048 5324
rect 10100 5352 10106 5364
rect 15470 5352 15476 5364
rect 10100 5324 15476 5352
rect 10100 5312 10106 5324
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 17865 5355 17923 5361
rect 17865 5321 17877 5355
rect 17911 5352 17923 5355
rect 18046 5352 18052 5364
rect 17911 5324 18052 5352
rect 17911 5321 17923 5324
rect 17865 5315 17923 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 19168 5324 20729 5352
rect 658 5244 664 5296
rect 716 5284 722 5296
rect 4154 5284 4160 5296
rect 716 5256 4160 5284
rect 716 5244 722 5256
rect 4154 5244 4160 5256
rect 4212 5284 4218 5296
rect 4433 5287 4491 5293
rect 4433 5284 4445 5287
rect 4212 5256 4445 5284
rect 4212 5244 4218 5256
rect 4433 5253 4445 5256
rect 4479 5253 4491 5287
rect 4433 5247 4491 5253
rect 5077 5287 5135 5293
rect 5077 5253 5089 5287
rect 5123 5284 5135 5287
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 5123 5256 6653 5284
rect 5123 5253 5135 5256
rect 5077 5247 5135 5253
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1854 5216 1860 5228
rect 1719 5188 1860 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 3142 5148 3148 5160
rect 2424 5120 3148 5148
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 2038 5080 2044 5092
rect 1811 5052 2044 5080
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 2038 5040 2044 5052
rect 2096 5080 2102 5092
rect 2424 5080 2452 5120
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3418 5148 3424 5160
rect 3375 5120 3424 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 3878 5148 3884 5160
rect 3839 5120 3884 5148
rect 3878 5108 3884 5120
rect 3936 5148 3942 5160
rect 4614 5148 4620 5160
rect 3936 5120 4620 5148
rect 3936 5108 3942 5120
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5184 5157 5212 5256
rect 6641 5253 6653 5256
rect 6687 5284 6699 5287
rect 7190 5284 7196 5296
rect 6687 5256 7196 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 7190 5244 7196 5256
rect 7248 5284 7254 5296
rect 11330 5284 11336 5296
rect 7248 5256 8708 5284
rect 11291 5256 11336 5284
rect 7248 5244 7254 5256
rect 8680 5225 8708 5256
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 13630 5284 13636 5296
rect 13591 5256 13636 5284
rect 13630 5244 13636 5256
rect 13688 5244 13694 5296
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 13964 5256 15117 5284
rect 13964 5244 13970 5256
rect 15105 5253 15117 5256
rect 15151 5284 15163 5287
rect 15194 5284 15200 5296
rect 15151 5256 15200 5284
rect 15151 5253 15163 5256
rect 15105 5247 15163 5253
rect 15194 5244 15200 5256
rect 15252 5284 15258 5296
rect 15252 5256 16344 5284
rect 15252 5244 15258 5256
rect 6273 5219 6331 5225
rect 6273 5185 6285 5219
rect 6319 5216 6331 5219
rect 8665 5219 8723 5225
rect 6319 5188 7420 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5117 5227 5151
rect 5169 5111 5227 5117
rect 5258 5108 5264 5160
rect 5316 5148 5322 5160
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 5316 5120 5733 5148
rect 5316 5108 5322 5120
rect 5721 5117 5733 5120
rect 5767 5148 5779 5151
rect 6288 5148 6316 5179
rect 7098 5148 7104 5160
rect 5767 5120 6316 5148
rect 7059 5120 7104 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7392 5157 7420 5188
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 8711 5188 10241 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 8110 5148 8116 5160
rect 7423 5120 8116 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 9048 5157 9076 5188
rect 10229 5185 10241 5188
rect 10275 5216 10287 5219
rect 12158 5216 12164 5228
rect 10275 5188 12164 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 10134 5148 10140 5160
rect 9355 5120 10140 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 2682 5080 2688 5092
rect 2096 5052 2452 5080
rect 2643 5052 2688 5080
rect 2096 5040 2102 5052
rect 2682 5040 2688 5052
rect 2740 5040 2746 5092
rect 4157 5083 4215 5089
rect 4157 5049 4169 5083
rect 4203 5080 4215 5083
rect 4890 5080 4896 5092
rect 4203 5052 4896 5080
rect 4203 5049 4215 5052
rect 4157 5043 4215 5049
rect 4890 5040 4896 5052
rect 4948 5040 4954 5092
rect 8294 5080 8300 5092
rect 8207 5052 8300 5080
rect 8294 5040 8300 5052
rect 8352 5080 8358 5092
rect 9324 5080 9352 5111
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 10612 5157 10640 5188
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12526 5216 12532 5228
rect 12487 5188 12532 5216
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 13170 5216 13176 5228
rect 13131 5188 13176 5216
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15378 5216 15384 5228
rect 15335 5188 15384 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16316 5216 16344 5256
rect 16390 5244 16396 5296
rect 16448 5284 16454 5296
rect 19168 5284 19196 5324
rect 20717 5321 20729 5324
rect 20763 5352 20775 5355
rect 20990 5352 20996 5364
rect 20763 5324 20996 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 16448 5256 19196 5284
rect 24121 5287 24179 5293
rect 16448 5244 16454 5256
rect 24121 5253 24133 5287
rect 24167 5284 24179 5287
rect 25590 5284 25596 5296
rect 24167 5256 25596 5284
rect 24167 5253 24179 5256
rect 24121 5247 24179 5253
rect 25590 5244 25596 5256
rect 25648 5244 25654 5296
rect 17678 5216 17684 5228
rect 16316 5188 17684 5216
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18414 5216 18420 5228
rect 18187 5188 18420 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 19150 5216 19156 5228
rect 18831 5188 19156 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 21177 5219 21235 5225
rect 21177 5216 21189 5219
rect 19392 5188 21189 5216
rect 19392 5176 19398 5188
rect 21177 5185 21189 5188
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 10781 5151 10839 5157
rect 10781 5148 10793 5151
rect 10744 5120 10793 5148
rect 10744 5108 10750 5120
rect 10781 5117 10793 5120
rect 10827 5117 10839 5151
rect 10781 5111 10839 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14090 5148 14096 5160
rect 14047 5120 14096 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14090 5108 14096 5120
rect 14148 5148 14154 5160
rect 16945 5151 17003 5157
rect 14148 5120 14596 5148
rect 14148 5108 14154 5120
rect 9490 5080 9496 5092
rect 8352 5052 9352 5080
rect 9451 5052 9496 5080
rect 8352 5040 8358 5052
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 11057 5083 11115 5089
rect 11057 5049 11069 5083
rect 11103 5080 11115 5083
rect 12158 5080 12164 5092
rect 11103 5052 12164 5080
rect 11103 5049 11115 5052
rect 11057 5043 11115 5049
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 12618 5040 12624 5092
rect 12676 5080 12682 5092
rect 14568 5089 14596 5120
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17770 5148 17776 5160
rect 16991 5120 17776 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5117 19763 5151
rect 19705 5111 19763 5117
rect 14553 5083 14611 5089
rect 12676 5052 12721 5080
rect 12676 5040 12682 5052
rect 14553 5049 14565 5083
rect 14599 5080 14611 5083
rect 15381 5083 15439 5089
rect 14599 5052 15332 5080
rect 14599 5049 14611 5052
rect 14553 5043 14611 5049
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 3326 5012 3332 5024
rect 1912 4984 3332 5012
rect 1912 4972 1918 4984
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 5258 5012 5264 5024
rect 5219 4984 5264 5012
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6914 5012 6920 5024
rect 6875 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 11974 5012 11980 5024
rect 11931 4984 11980 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12636 5012 12664 5040
rect 14182 5012 14188 5024
rect 12299 4984 12664 5012
rect 14143 4984 14188 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 15304 5012 15332 5052
rect 15381 5049 15393 5083
rect 15427 5080 15439 5083
rect 16206 5080 16212 5092
rect 15427 5052 16212 5080
rect 15427 5049 15439 5052
rect 15381 5043 15439 5049
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 18233 5083 18291 5089
rect 18233 5049 18245 5083
rect 18279 5049 18291 5083
rect 19613 5083 19671 5089
rect 19613 5080 19625 5083
rect 18233 5043 18291 5049
rect 18984 5052 19625 5080
rect 15746 5012 15752 5024
rect 15304 4984 15752 5012
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 16172 4984 16497 5012
rect 16172 4972 16178 4984
rect 16485 4981 16497 4984
rect 16531 5012 16543 5015
rect 16850 5012 16856 5024
rect 16531 4984 16856 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16850 4972 16856 4984
rect 16908 5012 16914 5024
rect 17586 5012 17592 5024
rect 16908 4984 17592 5012
rect 16908 4972 16914 4984
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18248 5012 18276 5043
rect 18104 4984 18276 5012
rect 18104 4972 18110 4984
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 18984 5012 19012 5052
rect 19613 5049 19625 5052
rect 19659 5049 19671 5083
rect 19613 5043 19671 5049
rect 18380 4984 19012 5012
rect 18380 4972 18386 4984
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 19300 4984 19441 5012
rect 19300 4972 19306 4984
rect 19429 4981 19441 4984
rect 19475 5012 19487 5015
rect 19720 5012 19748 5111
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20772 5120 21097 5148
rect 20772 5108 20778 5120
rect 21085 5117 21097 5120
rect 21131 5148 21143 5151
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 21131 5120 21281 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 23934 5148 23940 5160
rect 23895 5120 23940 5148
rect 21269 5111 21327 5117
rect 23934 5108 23940 5120
rect 23992 5148 23998 5160
rect 24489 5151 24547 5157
rect 24489 5148 24501 5151
rect 23992 5120 24501 5148
rect 23992 5108 23998 5120
rect 24489 5117 24501 5120
rect 24535 5117 24547 5151
rect 24489 5111 24547 5117
rect 25108 5151 25166 5157
rect 25108 5117 25120 5151
rect 25154 5148 25166 5151
rect 25154 5120 25452 5148
rect 25154 5117 25166 5120
rect 25108 5111 25166 5117
rect 22186 5040 22192 5092
rect 22244 5080 22250 5092
rect 23290 5080 23296 5092
rect 22244 5052 23296 5080
rect 22244 5040 22250 5052
rect 23290 5040 23296 5052
rect 23348 5080 23354 5092
rect 23385 5083 23443 5089
rect 23385 5080 23397 5083
rect 23348 5052 23397 5080
rect 23348 5040 23354 5052
rect 23385 5049 23397 5052
rect 23431 5049 23443 5083
rect 23385 5043 23443 5049
rect 25424 5024 25452 5120
rect 19475 4984 19748 5012
rect 19475 4981 19487 4984
rect 19429 4975 19487 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 22462 5012 22468 5024
rect 20588 4984 22468 5012
rect 20588 4972 20594 4984
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 25179 5015 25237 5021
rect 25179 5012 25191 5015
rect 23532 4984 25191 5012
rect 23532 4972 23538 4984
rect 25179 4981 25191 4984
rect 25225 4981 25237 5015
rect 25179 4975 25237 4981
rect 25406 4972 25412 5024
rect 25464 5012 25470 5024
rect 25501 5015 25559 5021
rect 25501 5012 25513 5015
rect 25464 4984 25513 5012
rect 25464 4972 25470 4984
rect 25501 4981 25513 4984
rect 25547 4981 25559 5015
rect 25501 4975 25559 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3878 4808 3884 4820
rect 3559 4780 3884 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 5350 4808 5356 4820
rect 5311 4780 5356 4808
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 5994 4808 6000 4820
rect 5859 4780 6000 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 7926 4808 7932 4820
rect 7883 4780 7932 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8904 4780 9045 4808
rect 8904 4768 8910 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9272 4780 9413 4808
rect 9272 4768 9278 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 10686 4808 10692 4820
rect 9401 4771 9459 4777
rect 9784 4780 10272 4808
rect 10647 4780 10692 4808
rect 2130 4740 2136 4752
rect 2091 4712 2136 4740
rect 2130 4700 2136 4712
rect 2188 4700 2194 4752
rect 4427 4743 4485 4749
rect 4427 4709 4439 4743
rect 4473 4740 4485 4743
rect 4522 4740 4528 4752
rect 4473 4712 4528 4740
rect 4473 4709 4485 4712
rect 4427 4703 4485 4709
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 9784 4749 9812 4780
rect 6318 4743 6376 4749
rect 6318 4740 6330 4743
rect 6236 4712 6330 4740
rect 6236 4700 6242 4712
rect 6318 4709 6330 4712
rect 6364 4709 6376 4743
rect 6318 4703 6376 4709
rect 9769 4743 9827 4749
rect 9769 4709 9781 4743
rect 9815 4709 9827 4743
rect 9769 4703 9827 4709
rect 9861 4743 9919 4749
rect 9861 4709 9873 4743
rect 9907 4740 9919 4743
rect 10134 4740 10140 4752
rect 9907 4712 10140 4740
rect 9907 4709 9919 4712
rect 9861 4703 9919 4709
rect 10134 4700 10140 4712
rect 10192 4700 10198 4752
rect 10244 4740 10272 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11756 4780 11805 4808
rect 11756 4768 11762 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12434 4808 12440 4820
rect 12299 4780 12440 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12434 4768 12440 4780
rect 12492 4808 12498 4820
rect 18693 4811 18751 4817
rect 18693 4808 18705 4811
rect 12492 4780 18705 4808
rect 12492 4768 12498 4780
rect 18693 4777 18705 4780
rect 18739 4777 18751 4811
rect 18693 4771 18751 4777
rect 11149 4743 11207 4749
rect 11149 4740 11161 4743
rect 10244 4712 11161 4740
rect 11149 4709 11161 4712
rect 11195 4740 11207 4743
rect 11882 4740 11888 4752
rect 11195 4712 11888 4740
rect 11195 4709 11207 4712
rect 11149 4703 11207 4709
rect 11882 4700 11888 4712
rect 11940 4700 11946 4752
rect 12529 4743 12587 4749
rect 12529 4709 12541 4743
rect 12575 4740 12587 4743
rect 12618 4740 12624 4752
rect 12575 4712 12624 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 12894 4700 12900 4752
rect 12952 4740 12958 4752
rect 12952 4712 13124 4740
rect 12952 4700 12958 4712
rect 2774 4672 2780 4684
rect 2735 4644 2780 4672
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3844 4644 4077 4672
rect 3844 4632 3850 4644
rect 4065 4641 4077 4644
rect 4111 4672 4123 4675
rect 5258 4672 5264 4684
rect 4111 4644 5264 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6638 4672 6644 4684
rect 6043 4644 6644 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 7156 4644 7297 4672
rect 7156 4632 7162 4644
rect 7285 4641 7297 4644
rect 7331 4672 7343 4675
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7331 4644 8033 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8021 4635 8079 4641
rect 8036 4604 8064 4635
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 13096 4672 13124 4712
rect 13446 4700 13452 4752
rect 13504 4740 13510 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 13504 4712 13645 4740
rect 13504 4700 13510 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 14826 4700 14832 4752
rect 14884 4740 14890 4752
rect 15610 4743 15668 4749
rect 15610 4740 15622 4743
rect 14884 4712 15622 4740
rect 14884 4700 14890 4712
rect 15610 4709 15622 4712
rect 15656 4740 15668 4743
rect 15930 4740 15936 4752
rect 15656 4712 15936 4740
rect 15656 4709 15668 4712
rect 15610 4703 15668 4709
rect 15930 4700 15936 4712
rect 15988 4740 15994 4752
rect 16114 4740 16120 4752
rect 15988 4712 16120 4740
rect 15988 4700 15994 4712
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 16482 4740 16488 4752
rect 16443 4712 16488 4740
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 18141 4743 18199 4749
rect 18141 4709 18153 4743
rect 18187 4740 18199 4743
rect 18414 4740 18420 4752
rect 18187 4712 18420 4740
rect 18187 4709 18199 4712
rect 18141 4703 18199 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 18506 4700 18512 4752
rect 18564 4740 18570 4752
rect 18564 4712 18609 4740
rect 18564 4700 18570 4712
rect 23290 4700 23296 4752
rect 23348 4740 23354 4752
rect 23348 4712 24751 4740
rect 23348 4700 23354 4712
rect 13909 4675 13967 4681
rect 13909 4672 13921 4675
rect 13096 4644 13921 4672
rect 13909 4641 13921 4644
rect 13955 4672 13967 4675
rect 13998 4672 14004 4684
rect 13955 4644 14004 4672
rect 13955 4641 13967 4644
rect 13909 4635 13967 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 14792 4644 15301 4672
rect 14792 4632 14798 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 16206 4672 16212 4684
rect 16119 4644 16212 4672
rect 15289 4635 15347 4641
rect 16206 4632 16212 4644
rect 16264 4672 16270 4684
rect 16390 4672 16396 4684
rect 16264 4644 16396 4672
rect 16264 4632 16270 4644
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 17092 4644 17141 4672
rect 17092 4632 17098 4644
rect 17129 4641 17141 4644
rect 17175 4641 17187 4675
rect 17129 4635 17187 4641
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4641 18659 4675
rect 19058 4672 19064 4684
rect 19019 4644 19064 4672
rect 18601 4635 18659 4641
rect 8662 4604 8668 4616
rect 8036 4576 8668 4604
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 10008 4576 10057 4604
rect 10008 4564 10014 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11330 4604 11336 4616
rect 11287 4576 11336 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4604 12495 4607
rect 14090 4604 14096 4616
rect 12483 4576 14096 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 18616 4604 18644 4635
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20864 4644 21005 4672
rect 20864 4632 20870 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 22002 4632 22008 4684
rect 22060 4672 22066 4684
rect 22554 4672 22560 4684
rect 22060 4644 22560 4672
rect 22060 4632 22066 4644
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 23014 4632 23020 4684
rect 23072 4672 23078 4684
rect 24723 4681 24751 4712
rect 23696 4675 23754 4681
rect 23696 4672 23708 4675
rect 23072 4644 23708 4672
rect 23072 4632 23078 4644
rect 23696 4641 23708 4644
rect 23742 4641 23754 4675
rect 23696 4635 23754 4641
rect 24708 4675 24766 4681
rect 24708 4641 24720 4675
rect 24754 4672 24766 4675
rect 25498 4672 25504 4684
rect 24754 4644 25504 4672
rect 24754 4641 24766 4644
rect 24708 4635 24766 4641
rect 25498 4632 25504 4644
rect 25556 4632 25562 4684
rect 18690 4604 18696 4616
rect 14240 4576 18696 4604
rect 14240 4564 14246 4576
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20312 4576 20913 4604
rect 20312 4564 20318 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 21726 4564 21732 4616
rect 21784 4604 21790 4616
rect 24811 4607 24869 4613
rect 24811 4604 24823 4607
rect 21784 4576 24823 4604
rect 21784 4564 21790 4576
rect 24811 4573 24823 4576
rect 24857 4573 24869 4607
rect 24811 4567 24869 4573
rect 12989 4539 13047 4545
rect 12989 4505 13001 4539
rect 13035 4536 13047 4539
rect 13446 4536 13452 4548
rect 13035 4508 13452 4536
rect 13035 4505 13047 4508
rect 12989 4499 13047 4505
rect 13446 4496 13452 4508
rect 13504 4496 13510 4548
rect 14550 4496 14556 4548
rect 14608 4536 14614 4548
rect 19242 4536 19248 4548
rect 14608 4508 19248 4536
rect 14608 4496 14614 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 22741 4539 22799 4545
rect 22741 4505 22753 4539
rect 22787 4536 22799 4539
rect 24946 4536 24952 4548
rect 22787 4508 24952 4536
rect 22787 4505 22799 4508
rect 22741 4499 22799 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4304 4440 4997 4468
rect 4304 4428 4310 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7190 4468 7196 4480
rect 6963 4440 7196 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 11480 4440 14105 4468
rect 11480 4428 11486 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 15105 4471 15163 4477
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 15378 4468 15384 4480
rect 15151 4440 15384 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 17310 4468 17316 4480
rect 17271 4440 17316 4468
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 23799 4471 23857 4477
rect 23799 4437 23811 4471
rect 23845 4468 23857 4471
rect 24670 4468 24676 4480
rect 23845 4440 24676 4468
rect 23845 4437 23857 4440
rect 23799 4431 23857 4437
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1728 4236 1777 4264
rect 1728 4224 1734 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 6638 4264 6644 4276
rect 6599 4236 6644 4264
rect 1765 4227 1823 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 8294 4264 8300 4276
rect 7147 4236 8300 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 8294 4224 8300 4236
rect 8352 4224 8358 4276
rect 8662 4264 8668 4276
rect 8575 4236 8668 4264
rect 8662 4224 8668 4236
rect 8720 4264 8726 4276
rect 9582 4264 9588 4276
rect 8720 4236 9588 4264
rect 8720 4224 8726 4236
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 17310 4264 17316 4276
rect 10980 4236 17316 4264
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2823 4100 3249 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3237 4097 3249 4100
rect 3283 4128 3295 4131
rect 6914 4128 6920 4140
rect 3283 4100 6920 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 8680 4128 8708 4224
rect 10686 4196 10692 4208
rect 9416 4168 10692 4196
rect 9416 4128 9444 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 10873 4199 10931 4205
rect 10873 4165 10885 4199
rect 10919 4196 10931 4199
rect 10980 4196 11008 4236
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 17420 4236 18276 4264
rect 10919 4168 11008 4196
rect 10919 4165 10931 4168
rect 10873 4159 10931 4165
rect 7852 4100 8708 4128
rect 9232 4100 9444 4128
rect 2038 4060 2044 4072
rect 1999 4032 2044 4060
rect 2038 4020 2044 4032
rect 2096 4020 2102 4072
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4029 5503 4063
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 5445 4023 5503 4029
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3599 3995 3657 4001
rect 3599 3992 3611 3995
rect 3191 3964 3611 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 3599 3961 3611 3964
rect 3645 3992 3657 3995
rect 5077 3995 5135 4001
rect 3645 3964 4568 3992
rect 3645 3961 3657 3964
rect 3599 3955 3657 3961
rect 4540 3936 4568 3964
rect 5077 3961 5089 3995
rect 5123 3992 5135 3995
rect 5460 3992 5488 4023
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 7852 4069 7880 4100
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 5736 4032 7481 4060
rect 5736 3992 5764 4032
rect 7469 4029 7481 4032
rect 7515 4060 7527 4063
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7515 4032 7849 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 9122 4060 9128 4072
rect 8343 4032 9128 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 5902 3992 5908 4004
rect 5123 3964 5764 3992
rect 5863 3964 5908 3992
rect 5123 3961 5135 3964
rect 5077 3955 5135 3961
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8128 3992 8156 4023
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9232 3992 9260 4100
rect 10980 4069 11008 4168
rect 14090 4156 14096 4208
rect 14148 4196 14154 4208
rect 14277 4199 14335 4205
rect 14277 4196 14289 4199
rect 14148 4168 14289 4196
rect 14148 4156 14154 4168
rect 14277 4165 14289 4168
rect 14323 4196 14335 4199
rect 17420 4196 17448 4236
rect 14323 4168 17448 4196
rect 14323 4165 14335 4168
rect 14277 4159 14335 4165
rect 17586 4156 17592 4208
rect 17644 4196 17650 4208
rect 17773 4199 17831 4205
rect 17773 4196 17785 4199
rect 17644 4168 17785 4196
rect 17644 4156 17650 4168
rect 17773 4165 17785 4168
rect 17819 4196 17831 4199
rect 17954 4196 17960 4208
rect 17819 4168 17960 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 18248 4196 18276 4236
rect 18598 4224 18604 4276
rect 18656 4264 18662 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18656 4236 18981 4264
rect 18656 4224 18662 4236
rect 18969 4233 18981 4236
rect 19015 4264 19027 4267
rect 19978 4264 19984 4276
rect 19015 4236 19984 4264
rect 19015 4233 19027 4236
rect 18969 4227 19027 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 22554 4264 22560 4276
rect 22515 4236 22560 4264
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24811 4267 24869 4273
rect 24811 4264 24823 4267
rect 24176 4236 24823 4264
rect 24176 4224 24182 4236
rect 24811 4233 24823 4236
rect 24857 4233 24869 4267
rect 25498 4264 25504 4276
rect 25459 4236 25504 4264
rect 24811 4227 24869 4233
rect 25498 4224 25504 4236
rect 25556 4224 25562 4276
rect 21082 4196 21088 4208
rect 18248 4168 21088 4196
rect 21082 4156 21088 4168
rect 21140 4156 21146 4208
rect 11054 4088 11060 4140
rect 11112 4128 11118 4140
rect 11425 4131 11483 4137
rect 11425 4128 11437 4131
rect 11112 4100 11437 4128
rect 11112 4088 11118 4100
rect 11425 4097 11437 4100
rect 11471 4097 11483 4131
rect 12434 4128 12440 4140
rect 12395 4100 12440 4128
rect 11425 4091 11483 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 14424 4100 15485 4128
rect 14424 4088 14430 4100
rect 15473 4097 15485 4100
rect 15519 4128 15531 4131
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 15519 4100 16681 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 19245 4131 19303 4137
rect 19245 4128 19257 4131
rect 18748 4100 19257 4128
rect 18748 4088 18754 4100
rect 19245 4097 19257 4100
rect 19291 4097 19303 4131
rect 19245 4091 19303 4097
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 23624 4100 24751 4128
rect 23624 4088 23630 4100
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 7708 3964 9260 3992
rect 9487 3995 9545 4001
rect 7708 3952 7714 3964
rect 9487 3961 9499 3995
rect 9533 3992 9545 3995
rect 9766 3992 9772 4004
rect 9533 3964 9772 3992
rect 9533 3961 9545 3964
rect 9487 3955 9545 3961
rect 3418 3884 3424 3936
rect 3476 3924 3482 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 3476 3896 4169 3924
rect 3476 3884 3482 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4522 3924 4528 3936
rect 4435 3896 4528 3924
rect 4157 3887 4215 3893
rect 4522 3884 4528 3896
rect 4580 3924 4586 3936
rect 6178 3924 6184 3936
rect 4580 3896 6184 3924
rect 4580 3884 4586 3896
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 9030 3924 9036 3936
rect 8943 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3924 9094 3936
rect 9502 3924 9530 3955
rect 9766 3952 9772 3964
rect 9824 3992 9830 4004
rect 11164 3992 11192 4023
rect 12158 4020 12164 4072
rect 12216 4060 12222 4072
rect 18046 4060 18052 4072
rect 12216 4032 18052 4060
rect 12216 4020 12222 4032
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 19797 4063 19855 4069
rect 19797 4060 19809 4063
rect 18196 4032 19809 4060
rect 18196 4020 18202 4032
rect 19797 4029 19809 4032
rect 19843 4029 19855 4063
rect 19797 4023 19855 4029
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4029 19947 4063
rect 19889 4023 19947 4029
rect 21453 4063 21511 4069
rect 21453 4029 21465 4063
rect 21499 4029 21511 4063
rect 21453 4023 21511 4029
rect 23728 4063 23786 4069
rect 23728 4029 23740 4063
rect 23774 4060 23786 4063
rect 24118 4060 24124 4072
rect 23774 4032 24124 4060
rect 23774 4029 23786 4032
rect 23728 4023 23786 4029
rect 11882 3992 11888 4004
rect 9824 3964 10456 3992
rect 11164 3964 11888 3992
rect 9824 3952 9830 3964
rect 10042 3924 10048 3936
rect 9088 3896 9530 3924
rect 10003 3896 10048 3924
rect 9088 3884 9094 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10192 3896 10333 3924
rect 10192 3884 10198 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10428 3924 10456 3964
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 12253 3995 12311 4001
rect 12253 3992 12265 3995
rect 12032 3964 12265 3992
rect 12032 3952 12038 3964
rect 12253 3961 12265 3964
rect 12299 3992 12311 3995
rect 12799 3995 12857 4001
rect 12799 3992 12811 3995
rect 12299 3964 12811 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12799 3961 12811 3964
rect 12845 3992 12857 3995
rect 14182 3992 14188 4004
rect 12845 3964 14188 3992
rect 12845 3961 12857 3964
rect 12799 3955 12857 3961
rect 14182 3952 14188 3964
rect 14240 3992 14246 4004
rect 15013 3995 15071 4001
rect 15013 3992 15025 3995
rect 14240 3964 15025 3992
rect 14240 3952 14246 3964
rect 15013 3961 15025 3964
rect 15059 3992 15071 3995
rect 15381 3995 15439 4001
rect 15381 3992 15393 3995
rect 15059 3964 15393 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 15381 3961 15393 3964
rect 15427 3992 15439 3995
rect 15835 3995 15893 4001
rect 15835 3992 15847 3995
rect 15427 3964 15847 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 15835 3961 15847 3964
rect 15881 3992 15893 3995
rect 15930 3992 15936 4004
rect 15881 3964 15936 3992
rect 15881 3961 15893 3964
rect 15835 3955 15893 3961
rect 15930 3952 15936 3964
rect 15988 3952 15994 4004
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18370 3995 18428 4001
rect 18370 3992 18382 3995
rect 18012 3964 18382 3992
rect 18012 3952 18018 3964
rect 18370 3961 18382 3964
rect 18416 3961 18428 3995
rect 18370 3955 18428 3961
rect 18506 3952 18512 4004
rect 18564 3992 18570 4004
rect 19613 3995 19671 4001
rect 19613 3992 19625 3995
rect 18564 3964 19625 3992
rect 18564 3952 18570 3964
rect 19613 3961 19625 3964
rect 19659 3992 19671 3995
rect 19904 3992 19932 4023
rect 21358 3992 21364 4004
rect 19659 3964 19932 3992
rect 21319 3964 21364 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 21358 3952 21364 3964
rect 21416 3952 21422 4004
rect 11992 3924 12020 3952
rect 13354 3924 13360 3936
rect 10428 3896 12020 3924
rect 13315 3896 13360 3924
rect 10321 3887 10379 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13998 3924 14004 3936
rect 13959 3896 14004 3924
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14458 3924 14464 3936
rect 14419 3896 14464 3924
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16942 3924 16948 3936
rect 16439 3896 16948 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 17402 3924 17408 3936
rect 17092 3896 17137 3924
rect 17363 3896 17408 3924
rect 17092 3884 17098 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19426 3924 19432 3936
rect 18932 3896 19432 3924
rect 18932 3884 18938 3896
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 20806 3924 20812 3936
rect 20680 3896 20812 3924
rect 20680 3884 20686 3896
rect 20806 3884 20812 3896
rect 20864 3884 20870 3936
rect 21082 3884 21088 3936
rect 21140 3924 21146 3936
rect 21177 3927 21235 3933
rect 21177 3924 21189 3927
rect 21140 3896 21189 3924
rect 21140 3884 21146 3896
rect 21177 3893 21189 3896
rect 21223 3924 21235 3927
rect 21468 3924 21496 4023
rect 24118 4020 24124 4032
rect 24176 4020 24182 4072
rect 24723 4069 24751 4100
rect 24708 4063 24766 4069
rect 24708 4029 24720 4063
rect 24754 4060 24766 4063
rect 25133 4063 25191 4069
rect 25133 4060 25145 4063
rect 24754 4032 25145 4060
rect 24754 4029 24766 4032
rect 24708 4023 24766 4029
rect 25133 4029 25145 4032
rect 25179 4029 25191 4063
rect 25133 4023 25191 4029
rect 23014 3952 23020 4004
rect 23072 3992 23078 4004
rect 24489 3995 24547 4001
rect 24489 3992 24501 3995
rect 23072 3964 24501 3992
rect 23072 3952 23078 3964
rect 24489 3961 24501 3964
rect 24535 3961 24547 3995
rect 24489 3955 24547 3961
rect 21223 3896 21496 3924
rect 21223 3893 21235 3896
rect 21177 3887 21235 3893
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 23799 3927 23857 3933
rect 23799 3924 23811 3927
rect 21600 3896 23811 3924
rect 21600 3884 21606 3896
rect 23799 3893 23811 3896
rect 23845 3893 23857 3927
rect 23799 3887 23857 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1535 3723 1593 3729
rect 1535 3689 1547 3723
rect 1581 3720 1593 3723
rect 1854 3720 1860 3732
rect 1581 3692 1860 3720
rect 1581 3689 1593 3692
rect 1535 3683 1593 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2038 3720 2044 3732
rect 1995 3692 2044 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2774 3720 2780 3732
rect 2363 3692 2780 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3510 3720 3516 3732
rect 3471 3692 3516 3720
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 3786 3720 3792 3732
rect 3747 3692 3792 3720
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5626 3720 5632 3732
rect 5307 3692 5632 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 7650 3720 7656 3732
rect 7611 3692 7656 3720
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 9784 3692 11161 3720
rect 2593 3655 2651 3661
rect 2593 3621 2605 3655
rect 2639 3652 2651 3655
rect 3418 3652 3424 3664
rect 2639 3624 3424 3652
rect 2639 3621 2651 3624
rect 2593 3615 2651 3621
rect 3418 3612 3424 3624
rect 3476 3612 3482 3664
rect 3878 3652 3884 3664
rect 3614 3624 3884 3652
rect 1464 3587 1522 3593
rect 1464 3553 1476 3587
rect 1510 3584 1522 3587
rect 1670 3584 1676 3596
rect 1510 3556 1676 3584
rect 1510 3553 1522 3556
rect 1464 3547 1522 3553
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 3510 3516 3516 3528
rect 2547 3488 3516 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3050 3448 3056 3460
rect 3011 3420 3056 3448
rect 3050 3408 3056 3420
rect 3108 3448 3114 3460
rect 3614 3448 3642 3624
rect 3878 3612 3884 3624
rect 3936 3652 3942 3664
rect 4157 3655 4215 3661
rect 4157 3652 4169 3655
rect 3936 3624 4169 3652
rect 3936 3612 3942 3624
rect 4157 3621 4169 3624
rect 4203 3621 4215 3655
rect 4157 3615 4215 3621
rect 4246 3612 4252 3664
rect 4304 3652 4310 3664
rect 4798 3652 4804 3664
rect 4304 3624 4349 3652
rect 4759 3624 4804 3652
rect 4304 3612 4310 3624
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 5991 3655 6049 3661
rect 5991 3621 6003 3655
rect 6037 3652 6049 3655
rect 6178 3652 6184 3664
rect 6037 3624 6184 3652
rect 6037 3621 6049 3624
rect 5991 3615 6049 3621
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8199 3655 8257 3661
rect 8199 3652 8211 3655
rect 8076 3624 8211 3652
rect 8076 3612 8082 3624
rect 8199 3621 8211 3624
rect 8245 3652 8257 3655
rect 9030 3652 9036 3664
rect 8245 3624 9036 3652
rect 8245 3621 8257 3624
rect 8199 3615 8257 3621
rect 9030 3612 9036 3624
rect 9088 3612 9094 3664
rect 9784 3661 9812 3692
rect 11149 3689 11161 3692
rect 11195 3720 11207 3723
rect 12342 3720 12348 3732
rect 11195 3692 12348 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 14274 3720 14280 3732
rect 12483 3692 14136 3720
rect 14235 3692 14280 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 9769 3655 9827 3661
rect 9769 3621 9781 3655
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 9861 3655 9919 3661
rect 9861 3621 9873 3655
rect 9907 3652 9919 3655
rect 10042 3652 10048 3664
rect 9907 3624 10048 3652
rect 9907 3621 9919 3624
rect 9861 3615 9919 3621
rect 10042 3612 10048 3624
rect 10100 3652 10106 3664
rect 11238 3652 11244 3664
rect 10100 3624 11244 3652
rect 10100 3612 10106 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 11664 3624 11713 3652
rect 11664 3612 11670 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 13170 3652 13176 3664
rect 13131 3624 13176 3652
rect 11701 3615 11759 3621
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 13265 3655 13323 3661
rect 13265 3621 13277 3655
rect 13311 3652 13323 3655
rect 13354 3652 13360 3664
rect 13311 3624 13360 3652
rect 13311 3621 13323 3624
rect 13265 3615 13323 3621
rect 13354 3612 13360 3624
rect 13412 3652 13418 3664
rect 13814 3652 13820 3664
rect 13412 3624 13820 3652
rect 13412 3612 13418 3624
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 14108 3652 14136 3692
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15013 3723 15071 3729
rect 15013 3720 15025 3723
rect 14792 3692 15025 3720
rect 14792 3680 14798 3692
rect 15013 3689 15025 3692
rect 15059 3689 15071 3723
rect 17402 3720 17408 3732
rect 15013 3683 15071 3689
rect 15212 3692 17408 3720
rect 15212 3652 15240 3692
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 18046 3720 18052 3732
rect 18007 3692 18052 3720
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19150 3720 19156 3732
rect 18739 3692 19156 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 14108 3624 15240 3652
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 15657 3655 15715 3661
rect 15657 3652 15669 3655
rect 15344 3624 15669 3652
rect 15344 3612 15350 3624
rect 15657 3621 15669 3624
rect 15703 3652 15715 3655
rect 16206 3652 16212 3664
rect 15703 3624 16212 3652
rect 15703 3621 15715 3624
rect 15657 3615 15715 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 17218 3652 17224 3664
rect 17179 3624 17224 3652
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 18966 3652 18972 3664
rect 18879 3624 18972 3652
rect 18966 3612 18972 3624
rect 19024 3652 19030 3664
rect 19242 3652 19248 3664
rect 19024 3624 19248 3652
rect 19024 3612 19030 3624
rect 19242 3612 19248 3624
rect 19300 3612 19306 3664
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 20864 3556 21005 3584
rect 20864 3544 20870 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 22278 3544 22284 3596
rect 22336 3584 22342 3596
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 22336 3556 22569 3584
rect 22336 3544 22342 3556
rect 22557 3553 22569 3556
rect 22603 3553 22615 3587
rect 24210 3584 24216 3596
rect 24171 3556 24216 3584
rect 22557 3547 22615 3553
rect 24210 3544 24216 3556
rect 24268 3544 24274 3596
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 5902 3516 5908 3528
rect 5675 3488 5908 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 5902 3476 5908 3488
rect 5960 3516 5966 3528
rect 6270 3516 6276 3528
rect 5960 3488 6276 3516
rect 5960 3476 5966 3488
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 7926 3516 7932 3528
rect 7883 3488 7932 3516
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 11882 3516 11888 3528
rect 11655 3488 11888 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12986 3516 12992 3528
rect 12299 3488 12992 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 13446 3476 13452 3488
rect 13504 3516 13510 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 13504 3488 14749 3516
rect 13504 3476 13510 3488
rect 14737 3485 14749 3488
rect 14783 3516 14795 3519
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 14783 3488 15577 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 15565 3485 15577 3488
rect 15611 3485 15623 3519
rect 15565 3479 15623 3485
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3516 16267 3519
rect 16390 3516 16396 3528
rect 16255 3488 16396 3516
rect 16255 3485 16267 3488
rect 16209 3479 16267 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 17126 3516 17132 3528
rect 16540 3488 17132 3516
rect 16540 3476 16546 3488
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 3108 3420 3642 3448
rect 3108 3408 3114 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7285 3451 7343 3457
rect 7285 3448 7297 3451
rect 6972 3420 7297 3448
rect 6972 3408 6978 3420
rect 7285 3417 7297 3420
rect 7331 3448 7343 3451
rect 9674 3448 9680 3460
rect 7331 3420 9680 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 10321 3451 10379 3457
rect 10321 3448 10333 3451
rect 10008 3420 10333 3448
rect 10008 3408 10014 3420
rect 10321 3417 10333 3420
rect 10367 3448 10379 3451
rect 12437 3451 12495 3457
rect 12437 3448 12449 3451
rect 10367 3420 12449 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 12437 3417 12449 3420
rect 12483 3417 12495 3451
rect 12437 3411 12495 3417
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 17034 3448 17040 3460
rect 14884 3420 17040 3448
rect 14884 3408 14890 3420
rect 17034 3408 17040 3420
rect 17092 3408 17098 3460
rect 6549 3383 6607 3389
rect 6549 3349 6561 3383
rect 6595 3380 6607 3383
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6595 3352 6837 3380
rect 6595 3349 6607 3352
rect 6549 3343 6607 3349
rect 6825 3349 6837 3352
rect 6871 3380 6883 3383
rect 7006 3380 7012 3392
rect 6871 3352 7012 3380
rect 6871 3349 6883 3352
rect 6825 3343 6883 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 8757 3383 8815 3389
rect 8757 3380 8769 3383
rect 8628 3352 8769 3380
rect 8628 3340 8634 3352
rect 8757 3349 8769 3352
rect 8803 3349 8815 3383
rect 8757 3343 8815 3349
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10689 3383 10747 3389
rect 10689 3380 10701 3383
rect 9456 3352 10701 3380
rect 9456 3340 9462 3352
rect 10689 3349 10701 3352
rect 10735 3380 10747 3383
rect 10870 3380 10876 3392
rect 10735 3352 10876 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12894 3380 12900 3392
rect 12855 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 17420 3380 17448 3479
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18874 3516 18880 3528
rect 17828 3488 18880 3516
rect 17828 3476 17834 3488
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19150 3516 19156 3528
rect 19111 3488 19156 3516
rect 19150 3476 19156 3488
rect 19208 3516 19214 3528
rect 20530 3516 20536 3528
rect 19208 3488 20536 3516
rect 19208 3476 19214 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20898 3516 20904 3528
rect 20859 3488 20904 3516
rect 20898 3476 20904 3488
rect 20956 3476 20962 3528
rect 22462 3516 22468 3528
rect 22423 3488 22468 3516
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 24026 3516 24032 3528
rect 23987 3488 24032 3516
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 17954 3408 17960 3460
rect 18012 3448 18018 3460
rect 20070 3448 20076 3460
rect 18012 3420 20076 3448
rect 18012 3408 18018 3420
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 18414 3380 18420 3392
rect 13504 3352 18420 3380
rect 13504 3340 13510 3352
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 19794 3380 19800 3392
rect 19755 3352 19800 3380
rect 19794 3340 19800 3352
rect 19852 3340 19858 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1673 3179 1731 3185
rect 1673 3176 1685 3179
rect 1636 3148 1685 3176
rect 1636 3136 1642 3148
rect 1673 3145 1685 3148
rect 1719 3145 1731 3179
rect 1673 3139 1731 3145
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 4295 3179 4353 3185
rect 4295 3176 4307 3179
rect 3752 3148 4307 3176
rect 3752 3136 3758 3148
rect 4295 3145 4307 3148
rect 4341 3145 4353 3179
rect 6641 3179 6699 3185
rect 6641 3176 6653 3179
rect 4295 3139 4353 3145
rect 5276 3148 6653 3176
rect 3050 3108 3056 3120
rect 3011 3080 3056 3108
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3476 3080 3801 3108
rect 3476 3068 3482 3080
rect 3789 3077 3801 3080
rect 3835 3077 3847 3111
rect 3789 3071 3847 3077
rect 2222 3000 2228 3052
rect 2280 3040 2286 3052
rect 5276 3049 5304 3148
rect 6641 3145 6653 3148
rect 6687 3176 6699 3179
rect 8478 3176 8484 3188
rect 6687 3148 8484 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9490 3176 9496 3188
rect 9451 3148 9496 3176
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 15565 3179 15623 3185
rect 15565 3176 15577 3179
rect 14516 3148 15577 3176
rect 14516 3136 14522 3148
rect 15565 3145 15577 3148
rect 15611 3176 15623 3179
rect 15611 3148 16252 3176
rect 15611 3145 15623 3148
rect 15565 3139 15623 3145
rect 7929 3111 7987 3117
rect 7929 3108 7941 3111
rect 6748 3080 7941 3108
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2280 3012 2513 3040
rect 2280 3000 2286 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 6236 3012 6285 3040
rect 6236 3000 6242 3012
rect 6273 3009 6285 3012
rect 6319 3040 6331 3043
rect 6748 3040 6776 3080
rect 7929 3077 7941 3080
rect 7975 3108 7987 3111
rect 8018 3108 8024 3120
rect 7975 3080 8024 3108
rect 7975 3077 7987 3080
rect 7929 3071 7987 3077
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 8297 3111 8355 3117
rect 8297 3077 8309 3111
rect 8343 3108 8355 3111
rect 8570 3108 8576 3120
rect 8343 3080 8576 3108
rect 8343 3077 8355 3080
rect 8297 3071 8355 3077
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 6914 3040 6920 3052
rect 6319 3012 6776 3040
rect 6875 3012 6920 3040
rect 6319 3009 6331 3012
rect 6273 3003 6331 3009
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 9398 3040 9404 3052
rect 8527 3012 9404 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9508 3040 9536 3136
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 12802 3108 12808 3120
rect 9640 3080 12808 3108
rect 9640 3068 9646 3080
rect 12802 3068 12808 3080
rect 12860 3068 12866 3120
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9508 3012 9965 3040
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 11238 3040 11244 3052
rect 11199 3012 11244 3040
rect 9953 3003 10011 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 16224 3049 16252 3148
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 17092 3148 19073 3176
rect 17092 3136 17098 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 19242 3176 19248 3188
rect 19203 3148 19248 3176
rect 19061 3139 19119 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 20806 3176 20812 3188
rect 20767 3148 20812 3176
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 24210 3176 24216 3188
rect 24171 3148 24216 3176
rect 24210 3136 24216 3148
rect 24268 3136 24274 3188
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 24903 3179 24961 3185
rect 24903 3176 24915 3179
rect 24820 3148 24915 3176
rect 24820 3136 24826 3148
rect 24903 3145 24915 3148
rect 24949 3145 24961 3179
rect 24903 3139 24961 3145
rect 17218 3108 17224 3120
rect 17131 3080 17224 3108
rect 17218 3068 17224 3080
rect 17276 3108 17282 3120
rect 18690 3108 18696 3120
rect 17276 3080 18696 3108
rect 17276 3068 17282 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 18782 3068 18788 3120
rect 18840 3108 18846 3120
rect 19889 3111 19947 3117
rect 19889 3108 19901 3111
rect 18840 3080 19901 3108
rect 18840 3068 18846 3080
rect 19889 3077 19901 3080
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3009 16267 3043
rect 16209 3003 16267 3009
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16485 3043 16543 3049
rect 16485 3040 16497 3043
rect 16448 3012 16497 3040
rect 16448 3000 16454 3012
rect 16485 3009 16497 3012
rect 16531 3009 16543 3043
rect 16485 3003 16543 3009
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17460 3012 18337 3040
rect 17460 3000 17466 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3040 19027 3043
rect 19150 3040 19156 3052
rect 19015 3012 19156 3040
rect 19015 3009 19027 3012
rect 18969 3003 19027 3009
rect 19150 3000 19156 3012
rect 19208 3000 19214 3052
rect 19242 3000 19248 3052
rect 19300 3040 19306 3052
rect 22186 3040 22192 3052
rect 19300 3012 22192 3040
rect 19300 3000 19306 3012
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 1464 2975 1522 2981
rect 1464 2941 1476 2975
rect 1510 2972 1522 2975
rect 4224 2975 4282 2981
rect 1510 2944 1624 2972
rect 1510 2941 1522 2944
rect 1464 2935 1522 2941
rect 1596 2836 1624 2944
rect 4224 2941 4236 2975
rect 4270 2972 4282 2975
rect 5905 2975 5963 2981
rect 4270 2944 4752 2972
rect 4270 2941 4282 2944
rect 4224 2935 4282 2941
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 1949 2907 2007 2913
rect 1949 2904 1961 2907
rect 1728 2876 1961 2904
rect 1728 2864 1734 2876
rect 1949 2873 1961 2876
rect 1995 2904 2007 2907
rect 2498 2904 2504 2916
rect 1995 2876 2504 2904
rect 1995 2873 2007 2876
rect 1949 2867 2007 2873
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 2639 2876 3556 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1596 2808 2329 2836
rect 2317 2805 2329 2808
rect 2363 2836 2375 2839
rect 3142 2836 3148 2848
rect 2363 2808 3148 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 3528 2845 3556 2876
rect 3513 2839 3571 2845
rect 3513 2805 3525 2839
rect 3559 2836 3571 2839
rect 3602 2836 3608 2848
rect 3559 2808 3608 2836
rect 3559 2805 3571 2808
rect 3513 2799 3571 2805
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 4724 2845 4752 2944
rect 5905 2941 5917 2975
rect 5951 2972 5963 2975
rect 5951 2944 6776 2972
rect 5951 2941 5963 2944
rect 5905 2935 5963 2941
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5350 2904 5356 2916
rect 5123 2876 5356 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 4798 2836 4804 2848
rect 4755 2808 4804 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 6748 2836 6776 2944
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 9824 2944 10358 2972
rect 9824 2932 9830 2944
rect 7006 2904 7012 2916
rect 6967 2876 7012 2904
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7098 2864 7104 2916
rect 7156 2904 7162 2916
rect 7561 2907 7619 2913
rect 7561 2904 7573 2907
rect 7156 2876 7573 2904
rect 7156 2864 7162 2876
rect 7561 2873 7573 2876
rect 7607 2904 7619 2907
rect 7607 2876 8064 2904
rect 7607 2873 7619 2876
rect 7561 2867 7619 2873
rect 7650 2836 7656 2848
rect 6748 2808 7656 2836
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 8036 2836 8064 2876
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 9125 2907 9183 2913
rect 8628 2876 8673 2904
rect 8628 2864 8634 2876
rect 9125 2873 9137 2907
rect 9171 2904 9183 2907
rect 10134 2904 10140 2916
rect 9171 2876 10140 2904
rect 9171 2873 9183 2876
rect 9125 2867 9183 2873
rect 10134 2864 10140 2876
rect 10192 2864 10198 2916
rect 10330 2913 10358 2944
rect 13786 2944 15209 2972
rect 10315 2907 10373 2913
rect 10315 2873 10327 2907
rect 10361 2873 10373 2907
rect 12802 2904 12808 2916
rect 12763 2876 12808 2904
rect 10315 2867 10373 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 12894 2864 12900 2916
rect 12952 2904 12958 2916
rect 13786 2904 13814 2944
rect 15197 2941 15209 2944
rect 15243 2972 15255 2975
rect 16022 2972 16028 2984
rect 15243 2944 16028 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2972 19119 2975
rect 19794 2972 19800 2984
rect 19107 2944 19800 2972
rect 19107 2941 19119 2944
rect 19061 2935 19119 2941
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2941 21511 2975
rect 23382 2972 23388 2984
rect 23295 2944 23388 2972
rect 21453 2935 21511 2941
rect 12952 2876 13814 2904
rect 12952 2864 12958 2876
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14598 2907 14656 2913
rect 14598 2904 14610 2907
rect 14240 2876 14610 2904
rect 14240 2864 14246 2876
rect 14598 2873 14610 2876
rect 14644 2873 14656 2907
rect 14598 2867 14656 2873
rect 16298 2864 16304 2916
rect 16356 2904 16362 2916
rect 18417 2907 18475 2913
rect 16356 2876 16401 2904
rect 16356 2864 16362 2876
rect 18417 2873 18429 2907
rect 18463 2904 18475 2907
rect 18598 2904 18604 2916
rect 18463 2876 18604 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 8754 2836 8760 2848
rect 8036 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 16025 2839 16083 2845
rect 13872 2808 13917 2836
rect 13872 2796 13878 2808
rect 16025 2805 16037 2839
rect 16071 2836 16083 2839
rect 16316 2836 16344 2864
rect 16071 2808 16344 2836
rect 17865 2839 17923 2845
rect 16071 2805 16083 2808
rect 16025 2799 16083 2805
rect 17865 2805 17877 2839
rect 17911 2836 17923 2839
rect 18432 2836 18460 2867
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19613 2907 19671 2913
rect 19613 2904 19625 2907
rect 19392 2876 19625 2904
rect 19392 2864 19398 2876
rect 19613 2873 19625 2876
rect 19659 2904 19671 2907
rect 20364 2904 20392 2935
rect 21358 2904 21364 2916
rect 19659 2876 20392 2904
rect 21319 2876 21364 2904
rect 19659 2873 19671 2876
rect 19613 2867 19671 2873
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 21174 2836 21180 2848
rect 17911 2808 18460 2836
rect 21135 2808 21180 2836
rect 17911 2805 17923 2808
rect 17865 2799 17923 2805
rect 21174 2796 21180 2808
rect 21232 2836 21238 2848
rect 21468 2836 21496 2935
rect 23382 2932 23388 2944
rect 23440 2972 23446 2984
rect 24854 2981 24860 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23440 2944 23673 2972
rect 23440 2932 23446 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 24832 2975 24860 2981
rect 24832 2972 24844 2975
rect 24767 2944 24844 2972
rect 23661 2935 23719 2941
rect 24832 2941 24844 2944
rect 24912 2972 24918 2984
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 24912 2944 25237 2972
rect 24832 2935 24860 2941
rect 24854 2932 24860 2935
rect 24912 2932 24918 2944
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 22336 2876 22477 2904
rect 22336 2864 22342 2876
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22465 2867 22523 2873
rect 23842 2836 23848 2848
rect 21232 2808 21496 2836
rect 23803 2808 23848 2836
rect 21232 2796 21238 2808
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1302 2592 1308 2644
rect 1360 2632 1366 2644
rect 1535 2635 1593 2641
rect 1535 2632 1547 2635
rect 1360 2604 1547 2632
rect 1360 2592 1366 2604
rect 1535 2601 1547 2604
rect 1581 2601 1593 2635
rect 1535 2595 1593 2601
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4387 2635 4445 2641
rect 4387 2632 4399 2635
rect 4028 2604 4399 2632
rect 4028 2592 4034 2604
rect 4387 2601 4399 2604
rect 4433 2601 4445 2635
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 4387 2595 4445 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 7926 2632 7932 2644
rect 7887 2604 7932 2632
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8619 2635 8677 2641
rect 8619 2632 8631 2635
rect 8352 2604 8631 2632
rect 8352 2592 8358 2604
rect 8619 2601 8631 2604
rect 8665 2601 8677 2635
rect 8619 2595 8677 2601
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 10781 2635 10839 2641
rect 10781 2632 10793 2635
rect 8812 2604 10793 2632
rect 8812 2592 8818 2604
rect 10781 2601 10793 2604
rect 10827 2601 10839 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10781 2595 10839 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11882 2632 11888 2644
rect 11379 2604 11888 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 14001 2635 14059 2641
rect 14001 2632 14013 2635
rect 13228 2604 14013 2632
rect 13228 2592 13234 2604
rect 14001 2601 14013 2604
rect 14047 2601 14059 2635
rect 15286 2632 15292 2644
rect 15247 2604 15292 2632
rect 14001 2595 14059 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 17126 2592 17132 2644
rect 17184 2632 17190 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17184 2604 17693 2632
rect 17184 2592 17190 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 18874 2592 18880 2644
rect 18932 2632 18938 2644
rect 19337 2635 19395 2641
rect 19337 2632 19349 2635
rect 18932 2604 19349 2632
rect 18932 2592 18938 2604
rect 19337 2601 19349 2604
rect 19383 2601 19395 2635
rect 19337 2595 19395 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2590 2564 2596 2576
rect 2363 2536 2596 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2590 2524 2596 2536
rect 2648 2524 2654 2576
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 4706 2564 4712 2576
rect 3191 2536 4712 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5169 2567 5227 2573
rect 5169 2533 5181 2567
rect 5215 2564 5227 2567
rect 5442 2564 5448 2576
rect 5215 2536 5448 2564
rect 5215 2533 5227 2536
rect 5169 2527 5227 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 6730 2564 6736 2576
rect 6691 2536 6736 2564
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 7190 2564 7196 2576
rect 7147 2536 7196 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 9950 2564 9956 2576
rect 9631 2536 9956 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 10870 2524 10876 2576
rect 10928 2564 10934 2576
rect 12345 2567 12403 2573
rect 12345 2564 12357 2567
rect 10928 2536 12357 2564
rect 10928 2524 10934 2536
rect 12345 2533 12357 2536
rect 12391 2564 12403 2567
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12391 2536 12817 2564
rect 12391 2533 12403 2536
rect 12345 2527 12403 2533
rect 12805 2533 12817 2536
rect 12851 2564 12863 2567
rect 16482 2564 16488 2576
rect 12851 2536 16488 2564
rect 12851 2533 12863 2536
rect 12805 2527 12863 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 16577 2567 16635 2573
rect 16577 2533 16589 2567
rect 16623 2564 16635 2567
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16623 2536 16865 2564
rect 16623 2533 16635 2536
rect 16577 2527 16635 2533
rect 16853 2533 16865 2536
rect 16899 2564 16911 2567
rect 18138 2564 18144 2576
rect 16899 2536 18144 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18506 2564 18512 2576
rect 18248 2536 18512 2564
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1854 2496 1860 2508
rect 1510 2468 1860 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 3878 2496 3884 2508
rect 3839 2468 3884 2496
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4316 2499 4374 2505
rect 4316 2465 4328 2499
rect 4362 2496 4374 2499
rect 5997 2499 6055 2505
rect 4362 2468 4844 2496
rect 4362 2465 4374 2468
rect 4316 2459 4374 2465
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3510 2428 3516 2440
rect 2547 2400 3516 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4816 2369 4844 2468
rect 5997 2465 6009 2499
rect 6043 2496 6055 2499
rect 8548 2499 8606 2505
rect 6043 2468 6868 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2428 5411 2431
rect 6840 2428 6868 2468
rect 8548 2465 8560 2499
rect 8594 2496 8606 2499
rect 8938 2496 8944 2508
rect 8594 2468 8944 2496
rect 8594 2465 8606 2468
rect 8548 2459 8606 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 14921 2499 14979 2505
rect 14921 2465 14933 2499
rect 14967 2496 14979 2499
rect 15562 2496 15568 2508
rect 14967 2468 15568 2496
rect 14967 2465 14979 2468
rect 14921 2459 14979 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 17460 2468 17505 2496
rect 17460 2456 17466 2468
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 5399 2400 6361 2428
rect 6840 2400 7021 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 4801 2363 4859 2369
rect 4801 2329 4813 2363
rect 4847 2360 4859 2363
rect 5534 2360 5540 2372
rect 4847 2332 5540 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 1854 2292 1860 2304
rect 1815 2264 1860 2292
rect 1854 2252 1860 2264
rect 1912 2252 1918 2304
rect 6333 2292 6361 2400
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7098 2428 7104 2440
rect 7055 2400 7104 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7650 2428 7656 2440
rect 7563 2400 7656 2428
rect 7650 2388 7656 2400
rect 7708 2428 7714 2440
rect 9582 2428 9588 2440
rect 7708 2400 9588 2428
rect 7708 2388 7714 2400
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 9861 2391 9919 2397
rect 9876 2360 9904 2391
rect 10134 2388 10140 2400
rect 10192 2428 10198 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 10192 2400 12725 2428
rect 10192 2388 10198 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12713 2391 12771 2397
rect 11146 2360 11152 2372
rect 9876 2332 11152 2360
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 12728 2360 12756 2391
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 14415 2400 16129 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 16117 2397 16129 2400
rect 16163 2428 16175 2431
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16163 2400 16773 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17000 2400 18061 2428
rect 17000 2388 17006 2400
rect 18049 2397 18061 2400
rect 18095 2428 18107 2431
rect 18248 2428 18276 2536
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 18690 2524 18696 2576
rect 18748 2564 18754 2576
rect 21177 2567 21235 2573
rect 21177 2564 21189 2567
rect 18748 2536 21189 2564
rect 18748 2524 18754 2536
rect 21177 2533 21189 2536
rect 21223 2533 21235 2567
rect 21177 2527 21235 2533
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2496 19119 2499
rect 19242 2496 19248 2508
rect 19107 2468 19248 2496
rect 19107 2465 19119 2468
rect 19061 2459 19119 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19484 2468 19901 2496
rect 19484 2456 19490 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20441 2459 20499 2465
rect 20916 2468 21281 2496
rect 18414 2428 18420 2440
rect 18095 2400 18276 2428
rect 18375 2400 18420 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 20916 2437 20944 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 21692 2468 22753 2496
rect 21692 2456 21698 2468
rect 22741 2465 22753 2468
rect 22787 2496 22799 2499
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22787 2468 23305 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 23992 2468 24041 2496
rect 23992 2456 23998 2468
rect 24029 2465 24041 2468
rect 24075 2496 24087 2499
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24075 2468 24593 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 24670 2456 24676 2508
rect 24728 2496 24734 2508
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24728 2468 25145 2496
rect 24728 2456 24734 2468
rect 25133 2465 25145 2468
rect 25179 2496 25191 2499
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25179 2468 25697 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 18524 2400 20913 2428
rect 13633 2363 13691 2369
rect 13633 2360 13645 2363
rect 12728 2332 13645 2360
rect 13633 2329 13645 2332
rect 13679 2329 13691 2363
rect 13633 2323 13691 2329
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 18524 2360 18552 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 16080 2332 18552 2360
rect 20073 2363 20131 2369
rect 16080 2320 16086 2332
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 20806 2360 20812 2372
rect 20119 2332 20812 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 20806 2320 20812 2332
rect 20864 2320 20870 2372
rect 22646 2320 22652 2372
rect 22704 2360 22710 2372
rect 24213 2363 24271 2369
rect 24213 2360 24225 2363
rect 22704 2332 24225 2360
rect 22704 2320 22710 2332
rect 24213 2329 24225 2332
rect 24259 2329 24271 2363
rect 24213 2323 24271 2329
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 6333 2264 8309 2292
rect 8297 2261 8309 2264
rect 8343 2292 8355 2295
rect 8846 2292 8852 2304
rect 8343 2264 8852 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 12069 2295 12127 2301
rect 12069 2261 12081 2295
rect 12115 2292 12127 2295
rect 12802 2292 12808 2304
rect 12115 2264 12808 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 15749 2295 15807 2301
rect 15749 2261 15761 2295
rect 15795 2292 15807 2295
rect 16390 2292 16396 2304
rect 15795 2264 16396 2292
rect 15795 2261 15807 2264
rect 15749 2255 15807 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 18414 2252 18420 2304
rect 18472 2292 18478 2304
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 18472 2264 19717 2292
rect 18472 2252 18478 2264
rect 19705 2261 19717 2264
rect 19751 2261 19763 2295
rect 19705 2255 19763 2261
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 22060 2264 22937 2292
rect 22060 2252 22066 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 24728 2264 25329 2292
rect 24728 2252 24734 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 3418 2048 3424 2100
rect 3476 2088 3482 2100
rect 6638 2088 6644 2100
rect 3476 2060 6644 2088
rect 3476 2048 3482 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 12710 2048 12716 2100
rect 12768 2088 12774 2100
rect 18414 2088 18420 2100
rect 12768 2060 18420 2088
rect 12768 2048 12774 2060
rect 18414 2048 18420 2060
rect 18472 2048 18478 2100
rect 4614 1980 4620 2032
rect 4672 2020 4678 2032
rect 8938 2020 8944 2032
rect 4672 1992 8944 2020
rect 4672 1980 4678 1992
rect 8938 1980 8944 1992
rect 8996 1980 9002 2032
rect 13998 1980 14004 2032
rect 14056 2020 14062 2032
rect 16850 2020 16856 2032
rect 14056 1992 16856 2020
rect 14056 1980 14062 1992
rect 16850 1980 16856 1992
rect 16908 1980 16914 2032
rect 14734 1912 14740 1964
rect 14792 1952 14798 1964
rect 21726 1952 21732 1964
rect 14792 1924 21732 1952
rect 14792 1912 14798 1924
rect 21726 1912 21732 1924
rect 21784 1912 21790 1964
rect 13998 184 14004 196
rect 6748 156 14004 184
rect 6748 128 6776 156
rect 13998 144 14004 156
rect 14056 144 14062 196
rect 6730 76 6736 128
rect 6788 76 6794 128
rect 9950 76 9956 128
rect 10008 116 10014 128
rect 18230 116 18236 128
rect 10008 88 18236 116
rect 10008 76 10014 88
rect 18230 76 18236 88
rect 18288 76 18294 128
rect 9122 8 9128 60
rect 9180 48 9186 60
rect 10962 48 10968 60
rect 9180 20 10968 48
rect 9180 8 9186 20
rect 10962 8 10968 20
rect 11020 8 11026 60
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1584 24395 1636 24404
rect 1584 24361 1593 24395
rect 1593 24361 1627 24395
rect 1627 24361 1636 24395
rect 1584 24352 1636 24361
rect 1492 24216 1544 24268
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1124 23808 1176 23860
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 1492 23672 1544 23724
rect 3424 23672 3476 23724
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 4896 23468 4948 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1400 22924 1452 22976
rect 1952 22924 2004 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2044 21335 2096 21344
rect 2044 21301 2053 21335
rect 2053 21301 2087 21335
rect 2087 21301 2096 21335
rect 2044 21292 2096 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1492 21088 1544 21140
rect 2044 21088 2096 21140
rect 2228 20952 2280 21004
rect 2596 20952 2648 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 1400 20204 1452 20256
rect 1860 20247 1912 20256
rect 1860 20213 1869 20247
rect 1869 20213 1903 20247
rect 1903 20213 1912 20247
rect 1860 20204 1912 20213
rect 2596 20247 2648 20256
rect 2596 20213 2605 20247
rect 2605 20213 2639 20247
rect 2639 20213 2648 20247
rect 2596 20204 2648 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 2228 20000 2280 20052
rect 2320 19864 2372 19916
rect 3332 19864 3384 19916
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 3332 19499 3384 19508
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 2136 19252 2188 19304
rect 3332 19184 3384 19236
rect 4804 19184 4856 19236
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 3516 19159 3568 19168
rect 3516 19125 3525 19159
rect 3525 19125 3559 19159
rect 3559 19125 3568 19159
rect 3516 19116 3568 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 112 18912 164 18964
rect 2044 18912 2096 18964
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 3976 18819 4028 18828
rect 3976 18785 3985 18819
rect 3985 18785 4019 18819
rect 4019 18785 4028 18819
rect 3976 18776 4028 18785
rect 20 18640 72 18692
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3424 18368 3476 18420
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 6000 18164 6052 18216
rect 2964 18139 3016 18148
rect 2964 18105 2973 18139
rect 2973 18105 3007 18139
rect 3007 18105 3016 18139
rect 2964 18096 3016 18105
rect 2688 18028 2740 18080
rect 3056 18028 3108 18080
rect 3976 18028 4028 18080
rect 5264 18028 5316 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 3516 17824 3568 17876
rect 4896 17824 4948 17876
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 4988 17688 5040 17740
rect 5540 17688 5592 17740
rect 3424 17620 3476 17672
rect 5172 17620 5224 17672
rect 1768 17484 1820 17536
rect 2504 17484 2556 17536
rect 3884 17484 3936 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1952 17280 2004 17332
rect 3240 17212 3292 17264
rect 3516 17144 3568 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 5540 17212 5592 17264
rect 5264 17187 5316 17196
rect 3608 17144 3660 17153
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 7564 17076 7616 17128
rect 3424 17051 3476 17060
rect 3424 17017 3433 17051
rect 3433 17017 3467 17051
rect 3467 17017 3476 17051
rect 3424 17008 3476 17017
rect 5356 17051 5408 17060
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 6000 17008 6052 17060
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 2872 16940 2924 16992
rect 4988 16940 5040 16992
rect 8116 16940 8168 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 2872 16736 2924 16788
rect 5264 16779 5316 16788
rect 5264 16745 5273 16779
rect 5273 16745 5307 16779
rect 5307 16745 5316 16779
rect 5264 16736 5316 16745
rect 2964 16668 3016 16720
rect 1584 16600 1636 16652
rect 2228 16532 2280 16584
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 2136 16464 2188 16516
rect 4436 16668 4488 16720
rect 5356 16711 5408 16720
rect 5356 16677 5365 16711
rect 5365 16677 5399 16711
rect 5399 16677 5408 16711
rect 5356 16668 5408 16677
rect 8024 16668 8076 16720
rect 3976 16643 4028 16652
rect 3976 16609 3985 16643
rect 3985 16609 4019 16643
rect 4019 16609 4028 16643
rect 3976 16600 4028 16609
rect 6276 16600 6328 16652
rect 6552 16600 6604 16652
rect 8116 16532 8168 16584
rect 3700 16464 3752 16516
rect 7564 16464 7616 16516
rect 2412 16396 2464 16448
rect 2504 16396 2556 16448
rect 7932 16396 7984 16448
rect 8576 16396 8628 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2964 16192 3016 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 8116 16192 8168 16244
rect 112 16056 164 16108
rect 3976 16124 4028 16176
rect 3516 16056 3568 16108
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 6000 16056 6052 16108
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8576 15988 8628 16040
rect 2136 15963 2188 15972
rect 2136 15929 2145 15963
rect 2145 15929 2179 15963
rect 2179 15929 2188 15963
rect 2136 15920 2188 15929
rect 2320 15920 2372 15972
rect 3516 15963 3568 15972
rect 3516 15929 3525 15963
rect 3525 15929 3559 15963
rect 3559 15929 3568 15963
rect 3516 15920 3568 15929
rect 4344 15963 4396 15972
rect 4344 15929 4353 15963
rect 4353 15929 4387 15963
rect 4387 15929 4396 15963
rect 5264 15963 5316 15972
rect 4344 15920 4396 15929
rect 5264 15929 5273 15963
rect 5273 15929 5307 15963
rect 5307 15929 5316 15963
rect 5264 15920 5316 15929
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 6828 15852 6880 15904
rect 7840 15920 7892 15972
rect 8024 15852 8076 15904
rect 8392 15852 8444 15904
rect 9312 15895 9364 15904
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2504 15648 2556 15700
rect 3700 15691 3752 15700
rect 3700 15657 3709 15691
rect 3709 15657 3743 15691
rect 3743 15657 3752 15691
rect 3700 15648 3752 15657
rect 5264 15648 5316 15700
rect 1676 15623 1728 15632
rect 1676 15589 1685 15623
rect 1685 15589 1719 15623
rect 1719 15589 1728 15623
rect 1676 15580 1728 15589
rect 3516 15580 3568 15632
rect 6644 15623 6696 15632
rect 6644 15589 6653 15623
rect 6653 15589 6687 15623
rect 6687 15589 6696 15623
rect 6644 15580 6696 15589
rect 8024 15623 8076 15632
rect 8024 15589 8033 15623
rect 8033 15589 8067 15623
rect 8067 15589 8076 15623
rect 8024 15580 8076 15589
rect 2412 15512 2464 15564
rect 5448 15555 5500 15564
rect 2780 15444 2832 15496
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 9312 15512 9364 15564
rect 6828 15487 6880 15496
rect 6828 15453 6837 15487
rect 6837 15453 6871 15487
rect 6871 15453 6880 15487
rect 6828 15444 6880 15453
rect 1860 15376 1912 15428
rect 2136 15419 2188 15428
rect 2136 15385 2145 15419
rect 2145 15385 2179 15419
rect 2179 15385 2188 15419
rect 2136 15376 2188 15385
rect 2688 15308 2740 15360
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 2780 15104 2832 15156
rect 2136 15036 2188 15088
rect 3792 15104 3844 15156
rect 5448 15104 5500 15156
rect 5172 15036 5224 15088
rect 6828 15036 6880 15088
rect 2320 14968 2372 15020
rect 2872 14968 2924 15020
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 6644 14968 6696 15020
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 2688 14832 2740 14884
rect 3700 14875 3752 14884
rect 3700 14841 3709 14875
rect 3709 14841 3743 14875
rect 3743 14841 3752 14875
rect 3700 14832 3752 14841
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 5264 14875 5316 14884
rect 3792 14832 3844 14841
rect 5264 14841 5273 14875
rect 5273 14841 5307 14875
rect 5307 14841 5316 14875
rect 5264 14832 5316 14841
rect 5356 14875 5408 14884
rect 5356 14841 5365 14875
rect 5365 14841 5399 14875
rect 5399 14841 5408 14875
rect 5356 14832 5408 14841
rect 8392 14764 8444 14816
rect 9864 14764 9916 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 4344 14560 4396 14612
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 5356 14603 5408 14612
rect 5356 14569 5365 14603
rect 5365 14569 5399 14603
rect 5399 14569 5408 14603
rect 5356 14560 5408 14569
rect 1768 14535 1820 14544
rect 1768 14501 1777 14535
rect 1777 14501 1811 14535
rect 1811 14501 1820 14535
rect 1768 14492 1820 14501
rect 2320 14535 2372 14544
rect 2320 14501 2329 14535
rect 2329 14501 2363 14535
rect 2363 14501 2372 14535
rect 2320 14492 2372 14501
rect 6460 14560 6512 14612
rect 7196 14603 7248 14612
rect 7196 14569 7205 14603
rect 7205 14569 7239 14603
rect 7239 14569 7248 14603
rect 7196 14560 7248 14569
rect 6276 14492 6328 14544
rect 2688 14424 2740 14476
rect 8392 14492 8444 14544
rect 9864 14492 9916 14544
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5264 14356 5316 14408
rect 5540 14356 5592 14408
rect 9680 14399 9732 14408
rect 2504 14220 2556 14272
rect 3700 14263 3752 14272
rect 3700 14229 3709 14263
rect 3709 14229 3743 14263
rect 3743 14229 3752 14263
rect 3700 14220 3752 14229
rect 3976 14220 4028 14272
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 8484 14220 8536 14272
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1768 14016 1820 14068
rect 6460 14016 6512 14068
rect 8392 14016 8444 14068
rect 9680 14016 9732 14068
rect 2320 13880 2372 13932
rect 9772 13948 9824 14000
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 2228 13787 2280 13796
rect 2228 13753 2237 13787
rect 2237 13753 2271 13787
rect 2271 13753 2280 13787
rect 2228 13744 2280 13753
rect 4344 13744 4396 13796
rect 6644 13812 6696 13864
rect 8392 13812 8444 13864
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 10876 13855 10928 13864
rect 2504 13676 2556 13728
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 6644 13719 6696 13728
rect 6644 13685 6653 13719
rect 6653 13685 6687 13719
rect 6687 13685 6696 13719
rect 6644 13676 6696 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 8576 13719 8628 13728
rect 8576 13685 8585 13719
rect 8585 13685 8619 13719
rect 8619 13685 8628 13719
rect 8576 13676 8628 13685
rect 9128 13744 9180 13796
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 10692 13744 10744 13796
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13472 1728 13524
rect 5540 13472 5592 13524
rect 9772 13472 9824 13524
rect 10876 13472 10928 13524
rect 3332 13404 3384 13456
rect 3792 13404 3844 13456
rect 5172 13404 5224 13456
rect 5816 13404 5868 13456
rect 6552 13404 6604 13456
rect 9312 13404 9364 13456
rect 10692 13447 10744 13456
rect 10692 13413 10701 13447
rect 10701 13413 10735 13447
rect 10735 13413 10744 13447
rect 10692 13404 10744 13413
rect 1584 13336 1636 13388
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 4252 13268 4304 13320
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 6000 13268 6052 13320
rect 6644 13268 6696 13320
rect 7656 13336 7708 13388
rect 9864 13336 9916 13388
rect 11888 13336 11940 13388
rect 2228 13200 2280 13252
rect 7932 13200 7984 13252
rect 9128 13200 9180 13252
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 9680 13200 9732 13252
rect 4068 13132 4120 13184
rect 6920 13132 6972 13184
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 9404 13175 9456 13184
rect 7012 13132 7064 13141
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 9588 13132 9640 13184
rect 10140 13132 10192 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 2412 12928 2464 12980
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 1492 12792 1544 12844
rect 2504 12792 2556 12844
rect 2596 12792 2648 12844
rect 4160 12724 4212 12776
rect 6000 12792 6052 12844
rect 5264 12724 5316 12776
rect 7656 12792 7708 12844
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 8392 12724 8444 12776
rect 9036 12792 9088 12844
rect 9312 12767 9364 12776
rect 2504 12699 2556 12708
rect 2504 12665 2513 12699
rect 2513 12665 2547 12699
rect 2547 12665 2556 12699
rect 2504 12656 2556 12665
rect 4252 12656 4304 12708
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 3792 12588 3844 12640
rect 6552 12588 6604 12640
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9496 12792 9548 12844
rect 9680 12724 9732 12776
rect 11060 12767 11112 12776
rect 8668 12656 8720 12708
rect 9772 12588 9824 12640
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 12900 12767 12952 12776
rect 10692 12656 10744 12708
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 11888 12699 11940 12708
rect 11888 12665 11897 12699
rect 11897 12665 11931 12699
rect 11931 12665 11940 12699
rect 11888 12656 11940 12665
rect 18604 12656 18656 12708
rect 11152 12588 11204 12640
rect 12716 12588 12768 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 1952 12384 2004 12393
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 6828 12384 6880 12436
rect 7104 12384 7156 12436
rect 11060 12427 11112 12436
rect 2780 12316 2832 12368
rect 4252 12359 4304 12368
rect 4252 12325 4261 12359
rect 4261 12325 4295 12359
rect 4295 12325 4304 12359
rect 4252 12316 4304 12325
rect 4804 12359 4856 12368
rect 4804 12325 4813 12359
rect 4813 12325 4847 12359
rect 4847 12325 4856 12359
rect 4804 12316 4856 12325
rect 6000 12316 6052 12368
rect 6920 12316 6972 12368
rect 9680 12316 9732 12368
rect 1584 12248 1636 12300
rect 6644 12291 6696 12300
rect 6644 12257 6653 12291
rect 6653 12257 6687 12291
rect 6687 12257 6696 12291
rect 6644 12248 6696 12257
rect 6736 12248 6788 12300
rect 8116 12248 8168 12300
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 11152 12384 11204 12436
rect 10508 12316 10560 12368
rect 11704 12291 11756 12300
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 2596 12180 2648 12232
rect 2872 12180 2924 12232
rect 1768 12112 1820 12164
rect 3792 12112 3844 12164
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 9864 12180 9916 12232
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 11796 12248 11848 12300
rect 13176 12248 13228 12300
rect 13820 12291 13872 12300
rect 13820 12257 13829 12291
rect 13829 12257 13863 12291
rect 13863 12257 13872 12291
rect 13820 12248 13872 12257
rect 12348 12180 12400 12232
rect 12992 12180 13044 12232
rect 13452 12180 13504 12232
rect 1860 12044 1912 12096
rect 4344 12044 4396 12096
rect 8024 12112 8076 12164
rect 9496 12112 9548 12164
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7840 12044 7892 12096
rect 10140 12044 10192 12096
rect 10876 12044 10928 12096
rect 13084 12044 13136 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 3240 11840 3292 11892
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 6736 11840 6788 11892
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 2780 11815 2832 11824
rect 2780 11781 2789 11815
rect 2789 11781 2823 11815
rect 2823 11781 2832 11815
rect 2780 11772 2832 11781
rect 1768 11747 1820 11756
rect 1768 11713 1777 11747
rect 1777 11713 1811 11747
rect 1811 11713 1820 11747
rect 1768 11704 1820 11713
rect 2504 11704 2556 11756
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 4896 11704 4948 11756
rect 5264 11704 5316 11756
rect 6644 11704 6696 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 13728 11840 13780 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 10048 11772 10100 11824
rect 12900 11772 12952 11824
rect 13176 11772 13228 11824
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 11980 11704 12032 11756
rect 12992 11704 13044 11756
rect 1952 11568 2004 11620
rect 3332 11611 3384 11620
rect 3332 11577 3341 11611
rect 3341 11577 3375 11611
rect 3375 11577 3384 11611
rect 3332 11568 3384 11577
rect 4896 11611 4948 11620
rect 3240 11500 3292 11552
rect 4896 11577 4905 11611
rect 4905 11577 4939 11611
rect 4939 11577 4948 11611
rect 4896 11568 4948 11577
rect 6000 11568 6052 11620
rect 4160 11500 4212 11552
rect 9128 11636 9180 11688
rect 9680 11636 9732 11688
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 9220 11568 9272 11620
rect 6552 11500 6604 11509
rect 8484 11500 8536 11552
rect 9036 11500 9088 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 11152 11636 11204 11688
rect 13084 11636 13136 11688
rect 13176 11636 13228 11688
rect 11244 11611 11296 11620
rect 11244 11577 11253 11611
rect 11253 11577 11287 11611
rect 11287 11577 11296 11611
rect 11244 11568 11296 11577
rect 13268 11568 13320 11620
rect 11060 11500 11112 11552
rect 11612 11500 11664 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 3608 11339 3660 11348
rect 3608 11305 3617 11339
rect 3617 11305 3651 11339
rect 3651 11305 3660 11339
rect 3608 11296 3660 11305
rect 2044 11271 2096 11280
rect 2044 11237 2053 11271
rect 2053 11237 2087 11271
rect 2087 11237 2096 11271
rect 2044 11228 2096 11237
rect 2780 11228 2832 11280
rect 4896 11296 4948 11348
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 6000 11296 6052 11348
rect 6736 11296 6788 11348
rect 8852 11296 8904 11348
rect 9680 11296 9732 11348
rect 11704 11296 11756 11348
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 6552 11228 6604 11280
rect 3240 11160 3292 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 13084 11228 13136 11280
rect 10784 11160 10836 11212
rect 11520 11203 11572 11212
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 8484 11024 8536 11076
rect 9588 11092 9640 11144
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 13636 11160 13688 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 15476 11160 15528 11212
rect 11428 11092 11480 11144
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 11888 11092 11940 11144
rect 9312 11024 9364 11076
rect 10876 11024 10928 11076
rect 1860 10956 1912 11008
rect 3332 10999 3384 11008
rect 3332 10965 3341 10999
rect 3341 10965 3375 10999
rect 3375 10965 3384 10999
rect 3332 10956 3384 10965
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 13544 11024 13596 11076
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1952 10752 2004 10804
rect 7656 10752 7708 10804
rect 11428 10752 11480 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 2228 10684 2280 10736
rect 6000 10684 6052 10736
rect 8576 10684 8628 10736
rect 10140 10684 10192 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 10784 10684 10836 10736
rect 10968 10684 11020 10736
rect 14096 10684 14148 10736
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 5816 10616 5868 10668
rect 7564 10616 7616 10668
rect 9404 10616 9456 10668
rect 3424 10548 3476 10600
rect 1308 10480 1360 10532
rect 1860 10480 1912 10532
rect 2228 10523 2280 10532
rect 2228 10489 2237 10523
rect 2237 10489 2271 10523
rect 2271 10489 2280 10523
rect 2228 10480 2280 10489
rect 2044 10412 2096 10464
rect 2412 10412 2464 10464
rect 3516 10412 3568 10464
rect 4528 10412 4580 10464
rect 5172 10480 5224 10532
rect 6552 10523 6604 10532
rect 6552 10489 6561 10523
rect 6561 10489 6595 10523
rect 6595 10489 6604 10523
rect 6552 10480 6604 10489
rect 6000 10412 6052 10464
rect 7380 10591 7432 10600
rect 6736 10480 6788 10532
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9496 10548 9548 10600
rect 13360 10548 13412 10600
rect 14556 10616 14608 10668
rect 15844 10548 15896 10600
rect 10692 10480 10744 10532
rect 11796 10480 11848 10532
rect 11980 10480 12032 10532
rect 7840 10412 7892 10464
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 11520 10412 11572 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 14740 10480 14792 10532
rect 15476 10480 15528 10532
rect 14464 10412 14516 10464
rect 15660 10412 15712 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1676 10140 1728 10192
rect 3516 10208 3568 10260
rect 3884 10208 3936 10260
rect 4804 10208 4856 10260
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 8392 10208 8444 10260
rect 9312 10208 9364 10260
rect 10692 10208 10744 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 8852 10140 8904 10192
rect 8944 10140 8996 10192
rect 13636 10208 13688 10260
rect 11520 10140 11572 10192
rect 5080 10072 5132 10124
rect 5264 10115 5316 10124
rect 5264 10081 5273 10115
rect 5273 10081 5307 10115
rect 5307 10081 5316 10115
rect 5264 10072 5316 10081
rect 5356 10072 5408 10124
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 7932 10072 7984 10124
rect 9404 10072 9456 10124
rect 9956 10072 10008 10124
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 12256 10072 12308 10124
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 13636 10072 13688 10124
rect 16488 10072 16540 10124
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7656 10004 7708 10056
rect 9036 10004 9088 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 15384 10004 15436 10056
rect 2320 9936 2372 9988
rect 5448 9936 5500 9988
rect 11888 9936 11940 9988
rect 4528 9868 4580 9920
rect 7840 9868 7892 9920
rect 8668 9868 8720 9920
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 11796 9868 11848 9920
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 16580 9868 16632 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 5264 9664 5316 9716
rect 7380 9664 7432 9716
rect 9496 9664 9548 9716
rect 11428 9664 11480 9716
rect 12164 9664 12216 9716
rect 13084 9664 13136 9716
rect 6828 9596 6880 9648
rect 7840 9596 7892 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 13636 9596 13688 9648
rect 2228 9528 2280 9580
rect 2596 9528 2648 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 9036 9528 9088 9580
rect 3424 9460 3476 9512
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 6000 9460 6052 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 12624 9528 12676 9580
rect 2136 9392 2188 9444
rect 2412 9392 2464 9444
rect 11612 9460 11664 9512
rect 12348 9460 12400 9512
rect 12532 9460 12584 9512
rect 15476 9503 15528 9512
rect 11152 9392 11204 9444
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 14004 9392 14056 9444
rect 15476 9469 15485 9503
rect 15485 9469 15519 9503
rect 15519 9469 15528 9503
rect 15476 9460 15528 9469
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 10140 9324 10192 9376
rect 12256 9324 12308 9376
rect 18236 9392 18288 9444
rect 16488 9324 16540 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 5356 9163 5408 9172
rect 5356 9129 5365 9163
rect 5365 9129 5399 9163
rect 5399 9129 5408 9163
rect 5356 9120 5408 9129
rect 7656 9120 7708 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 2504 9052 2556 9104
rect 4528 9052 4580 9104
rect 6276 9052 6328 9104
rect 9864 9052 9916 9104
rect 11336 9120 11388 9172
rect 12532 9120 12584 9172
rect 12808 9120 12860 9172
rect 13820 9120 13872 9172
rect 12900 9095 12952 9104
rect 12900 9061 12909 9095
rect 12909 9061 12943 9095
rect 12943 9061 12952 9095
rect 12900 9052 12952 9061
rect 12992 9052 13044 9104
rect 13912 9052 13964 9104
rect 15476 9095 15528 9104
rect 15476 9061 15485 9095
rect 15485 9061 15519 9095
rect 15519 9061 15528 9095
rect 15476 9052 15528 9061
rect 3884 8984 3936 9036
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 16948 8984 17000 9036
rect 18420 8984 18472 9036
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 5264 8916 5316 8968
rect 6552 8916 6604 8968
rect 12440 8916 12492 8968
rect 13636 8916 13688 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 17500 8916 17552 8968
rect 2964 8848 3016 8900
rect 4160 8848 4212 8900
rect 4896 8848 4948 8900
rect 5080 8848 5132 8900
rect 9128 8848 9180 8900
rect 11152 8891 11204 8900
rect 11152 8857 11161 8891
rect 11161 8857 11195 8891
rect 11195 8857 11204 8891
rect 11152 8848 11204 8857
rect 11796 8848 11848 8900
rect 13820 8848 13872 8900
rect 1952 8780 2004 8832
rect 2136 8823 2188 8832
rect 2136 8789 2145 8823
rect 2145 8789 2179 8823
rect 2179 8789 2188 8823
rect 2136 8780 2188 8789
rect 3148 8780 3200 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5172 8780 5224 8832
rect 12348 8780 12400 8832
rect 12532 8780 12584 8832
rect 14004 8823 14056 8832
rect 14004 8789 14013 8823
rect 14013 8789 14047 8823
rect 14047 8789 14056 8823
rect 14004 8780 14056 8789
rect 17132 8780 17184 8832
rect 18880 8780 18932 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2504 8576 2556 8628
rect 4988 8576 5040 8628
rect 6276 8619 6328 8628
rect 6276 8585 6285 8619
rect 6285 8585 6319 8619
rect 6319 8585 6328 8619
rect 6276 8576 6328 8585
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 2320 8551 2372 8560
rect 2320 8517 2329 8551
rect 2329 8517 2363 8551
rect 2363 8517 2372 8551
rect 2320 8508 2372 8517
rect 4896 8508 4948 8560
rect 5080 8440 5132 8492
rect 3148 8372 3200 8424
rect 8668 8576 8720 8628
rect 9404 8619 9456 8628
rect 9404 8585 9413 8619
rect 9413 8585 9447 8619
rect 9447 8585 9456 8619
rect 9404 8576 9456 8585
rect 9772 8576 9824 8628
rect 11152 8576 11204 8628
rect 12532 8576 12584 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 18420 8576 18472 8628
rect 7564 8508 7616 8560
rect 7840 8508 7892 8560
rect 8852 8508 8904 8560
rect 9956 8508 10008 8560
rect 12440 8508 12492 8560
rect 7472 8440 7524 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 9680 8440 9732 8492
rect 12992 8440 13044 8492
rect 13176 8440 13228 8492
rect 10048 8372 10100 8424
rect 11336 8415 11388 8424
rect 1768 8347 1820 8356
rect 1768 8313 1777 8347
rect 1777 8313 1811 8347
rect 1811 8313 1820 8347
rect 1768 8304 1820 8313
rect 1952 8304 2004 8356
rect 2596 8236 2648 8288
rect 5264 8347 5316 8356
rect 5264 8313 5273 8347
rect 5273 8313 5307 8347
rect 5307 8313 5316 8347
rect 5264 8304 5316 8313
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 6644 8304 6696 8356
rect 7932 8304 7984 8356
rect 8300 8347 8352 8356
rect 8300 8313 8309 8347
rect 8309 8313 8343 8347
rect 8343 8313 8352 8347
rect 8300 8304 8352 8313
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 14740 8440 14792 8492
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 16212 8372 16264 8424
rect 8852 8236 8904 8288
rect 11428 8236 11480 8288
rect 14280 8304 14332 8356
rect 15476 8304 15528 8356
rect 13176 8236 13228 8288
rect 14372 8236 14424 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4068 8032 4120 8084
rect 5356 8032 5408 8084
rect 8392 8032 8444 8084
rect 11520 8032 11572 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12900 8032 12952 8084
rect 13176 8032 13228 8084
rect 14188 8032 14240 8084
rect 14648 8032 14700 8084
rect 3148 8007 3200 8016
rect 3148 7973 3157 8007
rect 3157 7973 3191 8007
rect 3191 7973 3200 8007
rect 3148 7964 3200 7973
rect 4528 7964 4580 8016
rect 6184 7964 6236 8016
rect 9036 7964 9088 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2688 7939 2740 7948
rect 2688 7905 2697 7939
rect 2697 7905 2731 7939
rect 2731 7905 2740 7939
rect 2688 7896 2740 7905
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 4620 7939 4672 7948
rect 1768 7828 1820 7880
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 8944 7896 8996 7948
rect 9404 7896 9456 7948
rect 4712 7828 4764 7880
rect 2044 7692 2096 7744
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 6644 7803 6696 7812
rect 6644 7769 6653 7803
rect 6653 7769 6687 7803
rect 6687 7769 6696 7803
rect 6644 7760 6696 7769
rect 8116 7828 8168 7880
rect 9036 7828 9088 7880
rect 9772 7896 9824 7948
rect 11336 7964 11388 8016
rect 11428 8007 11480 8016
rect 11428 7973 11437 8007
rect 11437 7973 11471 8007
rect 11471 7973 11480 8007
rect 11428 7964 11480 7973
rect 12072 7964 12124 8016
rect 13360 7964 13412 8016
rect 13636 8007 13688 8016
rect 13636 7973 13645 8007
rect 13645 7973 13679 8007
rect 13679 7973 13688 8007
rect 13636 7964 13688 7973
rect 15384 8007 15436 8016
rect 15384 7973 15393 8007
rect 15393 7973 15427 8007
rect 15427 7973 15436 8007
rect 15384 7964 15436 7973
rect 15568 7964 15620 8016
rect 11152 7896 11204 7948
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 11888 7828 11940 7880
rect 11060 7760 11112 7812
rect 13268 7828 13320 7880
rect 17960 7939 18012 7948
rect 17960 7905 17969 7939
rect 17969 7905 18003 7939
rect 18003 7905 18012 7939
rect 17960 7896 18012 7905
rect 18696 7896 18748 7948
rect 23848 7896 23900 7948
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 7564 7735 7616 7744
rect 5540 7692 5592 7701
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 7932 7692 7984 7744
rect 8668 7692 8720 7744
rect 10232 7692 10284 7744
rect 11796 7692 11848 7744
rect 13728 7692 13780 7744
rect 16948 7692 17000 7744
rect 24216 7692 24268 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2964 7531 3016 7540
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 4712 7531 4764 7540
rect 2688 7463 2740 7472
rect 2688 7429 2697 7463
rect 2697 7429 2731 7463
rect 2731 7429 2740 7463
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 5448 7488 5500 7540
rect 7564 7488 7616 7540
rect 10784 7488 10836 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 11888 7488 11940 7540
rect 13360 7488 13412 7540
rect 15568 7488 15620 7540
rect 2688 7420 2740 7429
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 5172 7420 5224 7472
rect 5264 7420 5316 7472
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 5540 7352 5592 7404
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 10232 7463 10284 7472
rect 10232 7429 10241 7463
rect 10241 7429 10275 7463
rect 10275 7429 10284 7463
rect 10232 7420 10284 7429
rect 11244 7420 11296 7472
rect 4252 7284 4304 7336
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 8668 7284 8720 7336
rect 9772 7284 9824 7336
rect 5264 7259 5316 7268
rect 5264 7225 5273 7259
rect 5273 7225 5307 7259
rect 5307 7225 5316 7259
rect 5264 7216 5316 7225
rect 5448 7216 5500 7268
rect 6000 7148 6052 7200
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 6828 7148 6880 7200
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 7012 7216 7064 7225
rect 8300 7216 8352 7268
rect 13176 7352 13228 7404
rect 15384 7420 15436 7472
rect 10140 7284 10192 7336
rect 10692 7259 10744 7268
rect 10692 7225 10701 7259
rect 10701 7225 10735 7259
rect 10735 7225 10744 7259
rect 10692 7216 10744 7225
rect 11612 7216 11664 7268
rect 12532 7216 12584 7268
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9680 7148 9732 7200
rect 10048 7148 10100 7200
rect 12072 7148 12124 7200
rect 13176 7148 13228 7200
rect 14832 7284 14884 7336
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 16120 7259 16172 7268
rect 16120 7225 16129 7259
rect 16129 7225 16163 7259
rect 16163 7225 16172 7259
rect 16120 7216 16172 7225
rect 18052 7259 18104 7268
rect 18052 7225 18061 7259
rect 18061 7225 18095 7259
rect 18095 7225 18104 7259
rect 18052 7216 18104 7225
rect 14096 7148 14148 7200
rect 14832 7191 14884 7200
rect 14832 7157 14841 7191
rect 14841 7157 14875 7191
rect 14875 7157 14884 7191
rect 14832 7148 14884 7157
rect 15292 7148 15344 7200
rect 17132 7191 17184 7200
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 18236 7284 18288 7336
rect 17868 7148 17920 7157
rect 18696 7148 18748 7200
rect 19156 7148 19208 7200
rect 20904 7284 20956 7336
rect 21088 7191 21140 7200
rect 21088 7157 21097 7191
rect 21097 7157 21131 7191
rect 21131 7157 21140 7191
rect 21088 7148 21140 7157
rect 21640 7148 21692 7200
rect 22008 7148 22060 7200
rect 23848 7191 23900 7200
rect 23848 7157 23857 7191
rect 23857 7157 23891 7191
rect 23891 7157 23900 7191
rect 23848 7148 23900 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2044 6919 2096 6928
rect 2044 6885 2053 6919
rect 2053 6885 2087 6919
rect 2087 6885 2096 6919
rect 2044 6876 2096 6885
rect 5540 6944 5592 6996
rect 7012 6944 7064 6996
rect 8116 6944 8168 6996
rect 9220 6944 9272 6996
rect 9312 6944 9364 6996
rect 6184 6876 6236 6928
rect 7380 6876 7432 6928
rect 12716 6987 12768 6996
rect 11152 6876 11204 6928
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 13268 6944 13320 6996
rect 16212 6987 16264 6996
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 13452 6876 13504 6928
rect 3056 6808 3108 6860
rect 3792 6808 3844 6860
rect 7564 6808 7616 6860
rect 8668 6808 8720 6860
rect 9864 6808 9916 6860
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 4252 6740 4304 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 8576 6740 8628 6792
rect 10048 6783 10100 6792
rect 4620 6715 4672 6724
rect 4620 6681 4629 6715
rect 4629 6681 4663 6715
rect 4663 6681 4672 6715
rect 4620 6672 4672 6681
rect 8668 6672 8720 6724
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 13176 6808 13228 6860
rect 14280 6876 14332 6928
rect 18144 6876 18196 6928
rect 19064 6876 19116 6928
rect 16120 6808 16172 6860
rect 16764 6808 16816 6860
rect 20812 6851 20864 6860
rect 20812 6817 20821 6851
rect 20821 6817 20855 6851
rect 20855 6817 20864 6851
rect 20812 6808 20864 6817
rect 21824 6808 21876 6860
rect 24216 6808 24268 6860
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 11888 6740 11940 6792
rect 12256 6740 12308 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 16948 6740 17000 6792
rect 19340 6740 19392 6792
rect 23848 6740 23900 6792
rect 12348 6672 12400 6724
rect 1400 6604 1452 6656
rect 4436 6604 4488 6656
rect 4896 6647 4948 6656
rect 4896 6613 4905 6647
rect 4905 6613 4939 6647
rect 4939 6613 4948 6647
rect 4896 6604 4948 6613
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7932 6647 7984 6656
rect 7932 6613 7941 6647
rect 7941 6613 7975 6647
rect 7975 6613 7984 6647
rect 7932 6604 7984 6613
rect 8852 6604 8904 6656
rect 10140 6604 10192 6656
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 13176 6672 13228 6724
rect 17132 6672 17184 6724
rect 18788 6672 18840 6724
rect 24124 6672 24176 6724
rect 19156 6604 19208 6656
rect 19248 6604 19300 6656
rect 26792 6604 26844 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2872 6400 2924 6452
rect 3792 6400 3844 6452
rect 5540 6400 5592 6452
rect 7104 6400 7156 6452
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 7932 6400 7984 6452
rect 9496 6400 9548 6452
rect 10784 6400 10836 6452
rect 11336 6400 11388 6452
rect 13176 6400 13228 6452
rect 13268 6400 13320 6452
rect 14832 6400 14884 6452
rect 15292 6400 15344 6452
rect 16764 6443 16816 6452
rect 16764 6409 16773 6443
rect 16773 6409 16807 6443
rect 16807 6409 16816 6443
rect 16764 6400 16816 6409
rect 17960 6400 18012 6452
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19340 6400 19392 6452
rect 21824 6400 21876 6452
rect 24216 6400 24268 6452
rect 3056 6332 3108 6384
rect 9680 6332 9732 6384
rect 10140 6375 10192 6384
rect 10140 6341 10149 6375
rect 10149 6341 10183 6375
rect 10183 6341 10192 6375
rect 10140 6332 10192 6341
rect 2504 6264 2556 6316
rect 3240 6264 3292 6316
rect 4068 6264 4120 6316
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 8576 6196 8628 6248
rect 10048 6196 10100 6248
rect 3148 6060 3200 6112
rect 5448 6128 5500 6180
rect 9220 6128 9272 6180
rect 9864 6171 9916 6180
rect 9864 6137 9873 6171
rect 9873 6137 9907 6171
rect 9907 6137 9916 6171
rect 9864 6128 9916 6137
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 8116 6060 8168 6112
rect 9772 6060 9824 6112
rect 11980 6332 12032 6384
rect 14740 6332 14792 6384
rect 12716 6264 12768 6316
rect 12992 6264 13044 6316
rect 14372 6264 14424 6316
rect 15108 6264 15160 6316
rect 19248 6332 19300 6384
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 19432 6264 19484 6316
rect 14188 6196 14240 6248
rect 14832 6196 14884 6248
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 21548 6196 21600 6248
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 12624 6171 12676 6180
rect 12624 6137 12633 6171
rect 12633 6137 12667 6171
rect 12667 6137 12676 6171
rect 12624 6128 12676 6137
rect 13176 6171 13228 6180
rect 13176 6137 13185 6171
rect 13185 6137 13219 6171
rect 13219 6137 13228 6171
rect 13176 6128 13228 6137
rect 11428 6060 11480 6112
rect 11888 6060 11940 6112
rect 14648 6128 14700 6180
rect 15476 6128 15528 6180
rect 15936 6171 15988 6180
rect 15936 6137 15945 6171
rect 15945 6137 15979 6171
rect 15979 6137 15988 6171
rect 18144 6171 18196 6180
rect 15936 6128 15988 6137
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 16856 6060 16908 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17960 6060 18012 6112
rect 18972 6128 19024 6180
rect 21456 6128 21508 6180
rect 20444 6060 20496 6112
rect 20812 6060 20864 6112
rect 21088 6060 21140 6112
rect 23940 6060 23992 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 2780 5856 2832 5908
rect 1676 5831 1728 5840
rect 1676 5797 1685 5831
rect 1685 5797 1719 5831
rect 1719 5797 1728 5831
rect 1676 5788 1728 5797
rect 2044 5788 2096 5840
rect 4436 5856 4488 5908
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 6644 5856 6696 5908
rect 8668 5856 8720 5908
rect 11428 5856 11480 5908
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 15108 5899 15160 5908
rect 15108 5865 15117 5899
rect 15117 5865 15151 5899
rect 15151 5865 15160 5899
rect 15108 5856 15160 5865
rect 16212 5856 16264 5908
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 18144 5899 18196 5908
rect 3240 5831 3292 5840
rect 3240 5797 3249 5831
rect 3249 5797 3283 5831
rect 3283 5797 3292 5831
rect 3240 5788 3292 5797
rect 4160 5763 4212 5772
rect 4160 5729 4178 5763
rect 4178 5729 4212 5763
rect 4160 5720 4212 5729
rect 4712 5720 4764 5772
rect 5356 5763 5408 5772
rect 5356 5729 5365 5763
rect 5365 5729 5399 5763
rect 5399 5729 5408 5763
rect 5356 5720 5408 5729
rect 6000 5788 6052 5840
rect 9036 5788 9088 5840
rect 9220 5788 9272 5840
rect 11244 5831 11296 5840
rect 11244 5797 11253 5831
rect 11253 5797 11287 5831
rect 11287 5797 11296 5831
rect 11244 5788 11296 5797
rect 11980 5788 12032 5840
rect 13176 5788 13228 5840
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 19984 5856 20036 5908
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 11704 5720 11756 5772
rect 12532 5720 12584 5772
rect 13360 5720 13412 5772
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 15292 5763 15344 5772
rect 2964 5652 3016 5704
rect 6828 5652 6880 5704
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 13452 5652 13504 5704
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 16488 5695 16540 5704
rect 1860 5584 1912 5636
rect 12624 5584 12676 5636
rect 14004 5584 14056 5636
rect 5264 5559 5316 5568
rect 5264 5525 5273 5559
rect 5273 5525 5307 5559
rect 5307 5525 5316 5559
rect 5264 5516 5316 5525
rect 8852 5516 8904 5568
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10140 5516 10192 5525
rect 13544 5516 13596 5568
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 17868 5788 17920 5840
rect 19064 5788 19116 5840
rect 19524 5788 19576 5840
rect 19156 5720 19208 5772
rect 20904 5720 20956 5772
rect 20996 5763 21048 5772
rect 20996 5729 21005 5763
rect 21005 5729 21039 5763
rect 21039 5729 21048 5763
rect 22468 5763 22520 5772
rect 20996 5720 21048 5729
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 23296 5720 23348 5772
rect 18420 5652 18472 5704
rect 18512 5584 18564 5636
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 16304 5516 16356 5568
rect 23388 5516 23440 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 5540 5312 5592 5364
rect 7472 5312 7524 5364
rect 9772 5312 9824 5364
rect 10048 5312 10100 5364
rect 15476 5312 15528 5364
rect 18052 5312 18104 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 664 5244 716 5296
rect 4160 5244 4212 5296
rect 1860 5176 1912 5228
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2044 5040 2096 5092
rect 3148 5108 3200 5160
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 4620 5108 4672 5160
rect 7196 5244 7248 5296
rect 11336 5287 11388 5296
rect 11336 5253 11345 5287
rect 11345 5253 11379 5287
rect 11379 5253 11388 5287
rect 11336 5244 11388 5253
rect 13636 5287 13688 5296
rect 13636 5253 13645 5287
rect 13645 5253 13679 5287
rect 13679 5253 13688 5287
rect 13636 5244 13688 5253
rect 13912 5244 13964 5296
rect 15200 5244 15252 5296
rect 5264 5108 5316 5160
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 8116 5108 8168 5160
rect 2688 5083 2740 5092
rect 2688 5049 2697 5083
rect 2697 5049 2731 5083
rect 2731 5049 2740 5083
rect 2688 5040 2740 5049
rect 4896 5040 4948 5092
rect 8300 5083 8352 5092
rect 8300 5049 8309 5083
rect 8309 5049 8343 5083
rect 8343 5049 8352 5083
rect 10140 5108 10192 5160
rect 12164 5176 12216 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 15384 5176 15436 5228
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16396 5244 16448 5296
rect 20996 5312 21048 5364
rect 25596 5244 25648 5296
rect 17684 5176 17736 5228
rect 18420 5176 18472 5228
rect 19156 5176 19208 5228
rect 19340 5176 19392 5228
rect 10692 5108 10744 5160
rect 14096 5108 14148 5160
rect 9496 5083 9548 5092
rect 8300 5040 8352 5049
rect 9496 5049 9505 5083
rect 9505 5049 9539 5083
rect 9539 5049 9548 5083
rect 9496 5040 9548 5049
rect 12164 5040 12216 5092
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 17776 5108 17828 5160
rect 12624 5040 12676 5049
rect 1860 4972 1912 5024
rect 3332 4972 3384 5024
rect 5264 5015 5316 5024
rect 5264 4981 5273 5015
rect 5273 4981 5307 5015
rect 5307 4981 5316 5015
rect 5264 4972 5316 4981
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 11980 4972 12032 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 16212 5040 16264 5092
rect 15752 4972 15804 5024
rect 16120 4972 16172 5024
rect 16856 4972 16908 5024
rect 17592 4972 17644 5024
rect 18052 4972 18104 5024
rect 18328 4972 18380 5024
rect 19248 4972 19300 5024
rect 20720 5108 20772 5160
rect 23940 5151 23992 5160
rect 23940 5117 23949 5151
rect 23949 5117 23983 5151
rect 23983 5117 23992 5151
rect 23940 5108 23992 5117
rect 22192 5040 22244 5092
rect 23296 5040 23348 5092
rect 20536 4972 20588 5024
rect 22468 5015 22520 5024
rect 22468 4981 22477 5015
rect 22477 4981 22511 5015
rect 22511 4981 22520 5015
rect 22468 4972 22520 4981
rect 23480 4972 23532 5024
rect 25412 4972 25464 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 3884 4768 3936 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 6000 4768 6052 4820
rect 7932 4768 7984 4820
rect 8852 4768 8904 4820
rect 9220 4768 9272 4820
rect 10692 4811 10744 4820
rect 2136 4743 2188 4752
rect 2136 4709 2145 4743
rect 2145 4709 2179 4743
rect 2179 4709 2188 4743
rect 2136 4700 2188 4709
rect 4528 4700 4580 4752
rect 6184 4700 6236 4752
rect 10140 4700 10192 4752
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 11704 4768 11756 4820
rect 12440 4768 12492 4820
rect 11888 4700 11940 4752
rect 12624 4700 12676 4752
rect 12900 4700 12952 4752
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 3792 4632 3844 4684
rect 5264 4632 5316 4684
rect 6644 4632 6696 4684
rect 7104 4632 7156 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 13452 4700 13504 4752
rect 14832 4700 14884 4752
rect 15936 4700 15988 4752
rect 16120 4700 16172 4752
rect 16488 4743 16540 4752
rect 16488 4709 16497 4743
rect 16497 4709 16531 4743
rect 16531 4709 16540 4743
rect 16488 4700 16540 4709
rect 18420 4700 18472 4752
rect 18512 4743 18564 4752
rect 18512 4709 18521 4743
rect 18521 4709 18555 4743
rect 18555 4709 18564 4743
rect 18512 4700 18564 4709
rect 23296 4700 23348 4752
rect 14004 4632 14056 4684
rect 14740 4632 14792 4684
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 16396 4632 16448 4684
rect 17040 4632 17092 4684
rect 19064 4675 19116 4684
rect 8668 4564 8720 4616
rect 9956 4564 10008 4616
rect 11336 4564 11388 4616
rect 14096 4564 14148 4616
rect 14188 4564 14240 4616
rect 19064 4641 19073 4675
rect 19073 4641 19107 4675
rect 19107 4641 19116 4675
rect 19064 4632 19116 4641
rect 20812 4632 20864 4684
rect 22008 4632 22060 4684
rect 22560 4675 22612 4684
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 23020 4632 23072 4684
rect 25504 4632 25556 4684
rect 18696 4564 18748 4616
rect 20260 4564 20312 4616
rect 21732 4564 21784 4616
rect 13452 4496 13504 4548
rect 14556 4496 14608 4548
rect 19248 4496 19300 4548
rect 24952 4496 25004 4548
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 4252 4428 4304 4480
rect 7196 4428 7248 4480
rect 11428 4428 11480 4480
rect 15384 4428 15436 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 24676 4428 24728 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1676 4224 1728 4276
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 8300 4224 8352 4276
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 9588 4224 9640 4276
rect 6920 4088 6972 4140
rect 10692 4156 10744 4208
rect 17316 4224 17368 4276
rect 2044 4063 2096 4072
rect 2044 4029 2053 4063
rect 2053 4029 2087 4063
rect 2087 4029 2096 4063
rect 2044 4020 2096 4029
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 9128 4063 9180 4072
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 7656 3952 7708 4004
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 14096 4156 14148 4208
rect 17592 4156 17644 4208
rect 17960 4156 18012 4208
rect 18604 4224 18656 4276
rect 19984 4224 20036 4276
rect 22560 4267 22612 4276
rect 22560 4233 22569 4267
rect 22569 4233 22603 4267
rect 22603 4233 22612 4267
rect 22560 4224 22612 4233
rect 24124 4224 24176 4276
rect 25504 4267 25556 4276
rect 25504 4233 25513 4267
rect 25513 4233 25547 4267
rect 25547 4233 25556 4267
rect 25504 4224 25556 4233
rect 21088 4156 21140 4208
rect 11060 4088 11112 4140
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 12440 4088 12492 4097
rect 14372 4088 14424 4140
rect 18696 4088 18748 4140
rect 23572 4088 23624 4140
rect 3424 3884 3476 3936
rect 4528 3927 4580 3936
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 6184 3927 6236 3936
rect 4528 3884 4580 3893
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9772 3952 9824 4004
rect 12164 4020 12216 4072
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 18144 4020 18196 4072
rect 24124 4063 24176 4072
rect 11888 3995 11940 4004
rect 10048 3927 10100 3936
rect 9036 3884 9088 3893
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10140 3884 10192 3936
rect 11888 3961 11897 3995
rect 11897 3961 11931 3995
rect 11931 3961 11940 3995
rect 11888 3952 11940 3961
rect 11980 3952 12032 4004
rect 14188 3952 14240 4004
rect 15936 3952 15988 4004
rect 17960 3952 18012 4004
rect 18512 3952 18564 4004
rect 21364 3995 21416 4004
rect 21364 3961 21373 3995
rect 21373 3961 21407 3995
rect 21407 3961 21416 3995
rect 21364 3952 21416 3961
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 14464 3927 14516 3936
rect 14464 3893 14473 3927
rect 14473 3893 14507 3927
rect 14507 3893 14516 3927
rect 14464 3884 14516 3893
rect 16948 3884 17000 3936
rect 17040 3927 17092 3936
rect 17040 3893 17049 3927
rect 17049 3893 17083 3927
rect 17083 3893 17092 3927
rect 17408 3927 17460 3936
rect 17040 3884 17092 3893
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 18880 3884 18932 3936
rect 19432 3884 19484 3936
rect 20628 3884 20680 3936
rect 20812 3927 20864 3936
rect 20812 3893 20821 3927
rect 20821 3893 20855 3927
rect 20855 3893 20864 3927
rect 20812 3884 20864 3893
rect 21088 3884 21140 3936
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 23020 3952 23072 4004
rect 21548 3884 21600 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1860 3680 1912 3732
rect 2044 3680 2096 3732
rect 2780 3680 2832 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 5632 3680 5684 3732
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 3424 3612 3476 3664
rect 1676 3544 1728 3596
rect 3516 3476 3568 3528
rect 3056 3451 3108 3460
rect 3056 3417 3065 3451
rect 3065 3417 3099 3451
rect 3099 3417 3108 3451
rect 3884 3612 3936 3664
rect 4252 3655 4304 3664
rect 4252 3621 4261 3655
rect 4261 3621 4295 3655
rect 4295 3621 4304 3655
rect 4804 3655 4856 3664
rect 4252 3612 4304 3621
rect 4804 3621 4813 3655
rect 4813 3621 4847 3655
rect 4847 3621 4856 3655
rect 4804 3612 4856 3621
rect 6184 3612 6236 3664
rect 8024 3612 8076 3664
rect 9036 3612 9088 3664
rect 12348 3680 12400 3732
rect 14280 3723 14332 3732
rect 10048 3612 10100 3664
rect 11244 3612 11296 3664
rect 11612 3612 11664 3664
rect 13176 3655 13228 3664
rect 13176 3621 13185 3655
rect 13185 3621 13219 3655
rect 13219 3621 13228 3655
rect 13176 3612 13228 3621
rect 13360 3612 13412 3664
rect 13820 3612 13872 3664
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 14740 3680 14792 3732
rect 17408 3680 17460 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 19156 3680 19208 3732
rect 15292 3612 15344 3664
rect 16212 3612 16264 3664
rect 17224 3655 17276 3664
rect 17224 3621 17233 3655
rect 17233 3621 17267 3655
rect 17267 3621 17276 3655
rect 17224 3612 17276 3621
rect 18972 3655 19024 3664
rect 18972 3621 18981 3655
rect 18981 3621 19015 3655
rect 19015 3621 19024 3655
rect 18972 3612 19024 3621
rect 19248 3612 19300 3664
rect 20812 3544 20864 3596
rect 22284 3544 22336 3596
rect 24216 3587 24268 3596
rect 24216 3553 24225 3587
rect 24225 3553 24259 3587
rect 24259 3553 24268 3587
rect 24216 3544 24268 3553
rect 5908 3476 5960 3528
rect 6276 3476 6328 3528
rect 7932 3476 7984 3528
rect 11888 3476 11940 3528
rect 12992 3476 13044 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 16396 3476 16448 3528
rect 16488 3476 16540 3528
rect 17132 3519 17184 3528
rect 17132 3485 17141 3519
rect 17141 3485 17175 3519
rect 17175 3485 17184 3519
rect 17132 3476 17184 3485
rect 3056 3408 3108 3417
rect 6920 3408 6972 3460
rect 9680 3408 9732 3460
rect 9956 3408 10008 3460
rect 14832 3408 14884 3460
rect 17040 3408 17092 3460
rect 7012 3340 7064 3392
rect 8576 3340 8628 3392
rect 9404 3340 9456 3392
rect 10876 3340 10928 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13452 3340 13504 3392
rect 17776 3476 17828 3528
rect 18880 3519 18932 3528
rect 18880 3485 18889 3519
rect 18889 3485 18923 3519
rect 18923 3485 18932 3519
rect 18880 3476 18932 3485
rect 19156 3519 19208 3528
rect 19156 3485 19165 3519
rect 19165 3485 19199 3519
rect 19199 3485 19208 3519
rect 19156 3476 19208 3485
rect 20536 3476 20588 3528
rect 20904 3519 20956 3528
rect 20904 3485 20913 3519
rect 20913 3485 20947 3519
rect 20947 3485 20956 3519
rect 20904 3476 20956 3485
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 17960 3408 18012 3460
rect 20076 3408 20128 3460
rect 18420 3340 18472 3392
rect 19800 3383 19852 3392
rect 19800 3349 19809 3383
rect 19809 3349 19843 3383
rect 19843 3349 19852 3383
rect 19800 3340 19852 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1584 3136 1636 3188
rect 3700 3136 3752 3188
rect 3056 3111 3108 3120
rect 3056 3077 3065 3111
rect 3065 3077 3099 3111
rect 3099 3077 3108 3111
rect 3056 3068 3108 3077
rect 3424 3068 3476 3120
rect 2228 3000 2280 3052
rect 8484 3136 8536 3188
rect 9496 3179 9548 3188
rect 9496 3145 9505 3179
rect 9505 3145 9539 3179
rect 9539 3145 9548 3179
rect 9496 3136 9548 3145
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14188 3136 14240 3145
rect 14464 3136 14516 3188
rect 6184 3000 6236 3052
rect 8024 3068 8076 3120
rect 8576 3068 8628 3120
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 9404 3000 9456 3052
rect 9588 3068 9640 3120
rect 12808 3068 12860 3120
rect 11244 3043 11296 3052
rect 11244 3009 11253 3043
rect 11253 3009 11287 3043
rect 11287 3009 11296 3043
rect 11244 3000 11296 3009
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 17040 3136 17092 3188
rect 19248 3179 19300 3188
rect 19248 3145 19257 3179
rect 19257 3145 19291 3179
rect 19291 3145 19300 3179
rect 19248 3136 19300 3145
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 24768 3136 24820 3188
rect 17224 3111 17276 3120
rect 17224 3077 17233 3111
rect 17233 3077 17267 3111
rect 17267 3077 17276 3111
rect 17224 3068 17276 3077
rect 18696 3068 18748 3120
rect 18788 3068 18840 3120
rect 16396 3000 16448 3052
rect 17408 3000 17460 3052
rect 19156 3000 19208 3052
rect 19248 3000 19300 3052
rect 22192 3000 22244 3052
rect 1676 2864 1728 2916
rect 2504 2864 2556 2916
rect 3148 2796 3200 2848
rect 3608 2796 3660 2848
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 4804 2796 4856 2848
rect 9772 2932 9824 2984
rect 7012 2907 7064 2916
rect 7012 2873 7021 2907
rect 7021 2873 7055 2907
rect 7055 2873 7064 2907
rect 7012 2864 7064 2873
rect 7104 2864 7156 2916
rect 7656 2796 7708 2848
rect 8576 2907 8628 2916
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 10140 2864 10192 2916
rect 12808 2907 12860 2916
rect 12808 2873 12817 2907
rect 12817 2873 12851 2907
rect 12851 2873 12860 2907
rect 12808 2864 12860 2873
rect 12900 2907 12952 2916
rect 12900 2873 12909 2907
rect 12909 2873 12943 2907
rect 12943 2873 12952 2907
rect 16028 2932 16080 2984
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 23388 2975 23440 2984
rect 12900 2864 12952 2873
rect 14188 2864 14240 2916
rect 16304 2907 16356 2916
rect 16304 2873 16313 2907
rect 16313 2873 16347 2907
rect 16347 2873 16356 2907
rect 16304 2864 16356 2873
rect 8760 2796 8812 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 18604 2864 18656 2916
rect 19340 2864 19392 2916
rect 21364 2907 21416 2916
rect 21364 2873 21373 2907
rect 21373 2873 21407 2907
rect 21407 2873 21416 2907
rect 21364 2864 21416 2873
rect 21180 2839 21232 2848
rect 21180 2805 21189 2839
rect 21189 2805 21223 2839
rect 21223 2805 21232 2839
rect 23388 2941 23397 2975
rect 23397 2941 23431 2975
rect 23431 2941 23440 2975
rect 23388 2932 23440 2941
rect 24860 2975 24912 2984
rect 24860 2941 24878 2975
rect 24878 2941 24912 2975
rect 24860 2932 24912 2941
rect 22284 2864 22336 2916
rect 23848 2839 23900 2848
rect 21180 2796 21232 2805
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1308 2592 1360 2644
rect 3976 2592 4028 2644
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 8300 2592 8352 2644
rect 8760 2592 8812 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 11888 2592 11940 2644
rect 13176 2592 13228 2644
rect 15292 2635 15344 2644
rect 15292 2601 15301 2635
rect 15301 2601 15335 2635
rect 15335 2601 15344 2635
rect 15292 2592 15344 2601
rect 17132 2592 17184 2644
rect 18880 2592 18932 2644
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 4712 2524 4764 2576
rect 5448 2567 5500 2576
rect 5448 2533 5457 2567
rect 5457 2533 5491 2567
rect 5491 2533 5500 2567
rect 5448 2524 5500 2533
rect 6736 2567 6788 2576
rect 6736 2533 6745 2567
rect 6745 2533 6779 2567
rect 6779 2533 6788 2567
rect 6736 2524 6788 2533
rect 7196 2524 7248 2576
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 10876 2524 10928 2576
rect 16488 2524 16540 2576
rect 18144 2524 18196 2576
rect 18512 2567 18564 2576
rect 1860 2456 1912 2508
rect 3884 2499 3936 2508
rect 3884 2465 3893 2499
rect 3893 2465 3927 2499
rect 3927 2465 3936 2499
rect 3884 2456 3936 2465
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 8944 2499 8996 2508
rect 8944 2465 8953 2499
rect 8953 2465 8987 2499
rect 8987 2465 8996 2499
rect 8944 2456 8996 2465
rect 15568 2499 15620 2508
rect 15568 2465 15577 2499
rect 15577 2465 15611 2499
rect 15611 2465 15620 2499
rect 15568 2456 15620 2465
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 5540 2320 5592 2372
rect 1860 2295 1912 2304
rect 1860 2261 1869 2295
rect 1869 2261 1903 2295
rect 1903 2261 1912 2295
rect 1860 2252 1912 2261
rect 7104 2388 7156 2440
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 9588 2388 9640 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 12992 2431 13044 2440
rect 11152 2320 11204 2372
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 16948 2388 17000 2440
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 18696 2524 18748 2576
rect 19248 2456 19300 2508
rect 19432 2456 19484 2508
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 21640 2456 21692 2508
rect 23940 2456 23992 2508
rect 24676 2456 24728 2508
rect 16028 2320 16080 2372
rect 20812 2320 20864 2372
rect 22652 2320 22704 2372
rect 8852 2252 8904 2304
rect 12808 2252 12860 2304
rect 16396 2252 16448 2304
rect 18420 2252 18472 2304
rect 22008 2252 22060 2304
rect 24676 2252 24728 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 3424 2048 3476 2100
rect 6644 2048 6696 2100
rect 12716 2048 12768 2100
rect 18420 2048 18472 2100
rect 4620 1980 4672 2032
rect 8944 1980 8996 2032
rect 14004 1980 14056 2032
rect 16856 1980 16908 2032
rect 14740 1912 14792 1964
rect 21732 1912 21784 1964
rect 14004 144 14056 196
rect 6736 76 6788 128
rect 9956 76 10008 128
rect 18236 76 18288 128
rect 9128 8 9180 60
rect 10968 8 11020 60
<< metal2 >>
rect 1122 26888 1178 26897
rect 1122 26823 1178 26832
rect 110 24304 166 24313
rect 110 24239 166 24248
rect 18 19136 74 19145
rect 18 19071 74 19080
rect 32 18698 60 19071
rect 124 18970 152 24239
rect 1136 23866 1164 26823
rect 1582 25800 1638 25809
rect 1582 25735 1638 25744
rect 1596 24410 1624 25735
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 2686 24848 2742 24857
rect 2686 24783 2742 24792
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1492 24268 1544 24274
rect 1492 24210 1544 24216
rect 1124 23860 1176 23866
rect 1124 23802 1176 23808
rect 1504 23730 1532 24210
rect 2700 23866 2728 24783
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1412 22982 1440 23598
rect 1400 22976 1452 22982
rect 1400 22918 1452 22924
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1490 21720 1546 21729
rect 1596 21690 1624 22607
rect 1490 21655 1546 21664
rect 1584 21684 1636 21690
rect 1504 21146 1532 21655
rect 1584 21626 1636 21632
rect 1492 21140 1544 21146
rect 1492 21082 1544 21088
rect 1582 20632 1638 20641
rect 1582 20567 1638 20576
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 112 18964 164 18970
rect 112 18906 164 18912
rect 1412 18834 1440 20198
rect 1596 20058 1624 20567
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1582 19680 1638 19689
rect 1582 19615 1638 19624
rect 1596 19514 1624 19615
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 20 18692 72 18698
rect 20 18634 72 18640
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1582 17504 1638 17513
rect 1582 17439 1638 17448
rect 1596 16658 1624 17439
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16250 1624 16594
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 112 16108 164 16114
rect 112 16050 164 16056
rect 124 16017 152 16050
rect 110 16008 166 16017
rect 110 15943 166 15952
rect 1688 15638 1716 18022
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1688 15162 1716 15574
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1780 14550 1808 17478
rect 1872 15434 1900 20198
rect 1964 17338 1992 22918
rect 2044 21344 2096 21350
rect 2044 21286 2096 21292
rect 2056 21146 2084 21286
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 2228 21004 2280 21010
rect 2228 20946 2280 20952
rect 2596 21004 2648 21010
rect 2596 20946 2648 20952
rect 2240 20602 2268 20946
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2240 20058 2268 20538
rect 2608 20262 2636 20946
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2332 19514 2360 19858
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18970 2084 19110
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2148 18816 2176 19246
rect 2056 18788 2176 18816
rect 2504 18828 2556 18834
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1676 14408 1728 14414
rect 1582 14376 1638 14385
rect 1676 14350 1728 14356
rect 1582 14311 1638 14320
rect 1596 13394 1624 14311
rect 1688 13530 1716 14350
rect 1780 14074 1808 14486
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 12986 1624 13330
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 18 12200 74 12209
rect 18 12135 74 12144
rect 32 6633 60 12135
rect 1308 10532 1360 10538
rect 1308 10474 1360 10480
rect 18 6624 74 6633
rect 18 6559 74 6568
rect 664 5296 716 5302
rect 664 5238 716 5244
rect 110 2544 166 2553
rect 166 2502 244 2530
rect 110 2479 166 2488
rect 216 785 244 2502
rect 202 776 258 785
rect 202 711 258 720
rect 386 82 442 480
rect 676 82 704 5238
rect 1320 2650 1348 10474
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 6662 1440 7890
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 1308 2644 1360 2650
rect 1308 2586 1360 2592
rect 386 54 704 82
rect 1122 82 1178 480
rect 1412 82 1440 6598
rect 1504 4154 1532 12786
rect 1964 12442 1992 16934
rect 2056 13814 2084 18788
rect 2504 18770 2556 18776
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 16590 2268 17682
rect 2516 17542 2544 18770
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2148 15978 2176 16458
rect 2136 15972 2188 15978
rect 2136 15914 2188 15920
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15094 2176 15370
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2056 13786 2176 13814
rect 2240 13802 2268 16526
rect 2332 15978 2360 16730
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2516 16454 2544 16526
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2424 15570 2452 16390
rect 2516 15706 2544 16390
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14550 2360 14962
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2332 13938 2360 14486
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1582 12336 1638 12345
rect 1582 12271 1584 12280
rect 1636 12271 1638 12280
rect 1584 12242 1636 12248
rect 1596 11354 1624 12242
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1780 11762 1808 12106
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1872 11132 1900 12038
rect 1964 11626 1992 12378
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 1952 11144 2004 11150
rect 1872 11104 1952 11132
rect 1952 11086 2004 11092
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1872 10538 1900 10950
rect 1964 10810 1992 11086
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 2056 10470 2084 11222
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1676 10192 1728 10198
rect 1596 10152 1676 10180
rect 1596 9382 1624 10152
rect 1676 10134 1728 10140
rect 2148 9568 2176 13786
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 13258 2268 13738
rect 2516 13734 2544 14214
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2424 12986 2452 13262
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2424 12696 2452 12922
rect 2516 12850 2544 13670
rect 2608 12850 2636 20198
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3344 19514 3372 19858
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3344 19242 3372 19450
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 3436 18426 3464 23666
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2700 15366 2728 18022
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16794 2912 16934
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2976 16726 3004 18090
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2976 16250 3004 16662
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 14890 2728 15302
rect 2792 15162 2820 15438
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2884 15026 2912 15302
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2700 14482 2728 14826
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2504 12708 2556 12714
rect 2424 12668 2504 12696
rect 2504 12650 2556 12656
rect 2608 12238 2636 12786
rect 2792 12374 2820 13330
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2516 11762 2544 12174
rect 2792 11830 2820 12310
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2780 11280 2832 11286
rect 2780 11222 2832 11228
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2240 10538 2268 10678
rect 2792 10674 2820 11222
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2320 9988 2372 9994
rect 2320 9930 2372 9936
rect 2228 9580 2280 9586
rect 2148 9540 2228 9568
rect 2228 9522 2280 9528
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 7410 1624 9318
rect 2148 8838 2176 9386
rect 2332 9110 2360 9930
rect 2424 9450 2452 10406
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 1964 8362 1992 8774
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1780 7886 1808 8298
rect 1964 8090 1992 8298
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1964 7342 1992 8026
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 2056 6934 2084 7686
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2056 5846 2084 6870
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 1688 4826 1716 5782
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5234 1900 5578
rect 2056 5234 2084 5782
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 4282 1716 4762
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1504 4126 1624 4154
rect 1596 3194 1624 4126
rect 1872 3738 1900 4966
rect 2056 4826 2084 5034
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2056 4078 2084 4762
rect 2148 4758 2176 8774
rect 2332 8566 2360 9046
rect 2516 8634 2544 9046
rect 2608 8974 2636 9522
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2516 8276 2544 8570
rect 2596 8288 2648 8294
rect 2516 8248 2596 8276
rect 2596 8230 2648 8236
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5914 2544 6258
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2226 4992 2282 5001
rect 2226 4927 2282 4936
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2056 3738 2084 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1688 2922 1716 3538
rect 2240 3058 2268 4927
rect 2608 4672 2636 8230
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2700 7478 2728 7890
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2884 6458 2912 12174
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2976 7954 3004 8842
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2976 7546 3004 7890
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 3068 6866 3096 18022
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 3252 11898 3280 17206
rect 3344 13462 3372 18158
rect 3528 17882 3556 19110
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3988 18086 4016 18770
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17066 3464 17614
rect 3528 17202 3556 17818
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3516 16108 3568 16114
rect 3620 16096 3648 17138
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3712 16114 3740 16458
rect 3568 16068 3648 16096
rect 3700 16108 3752 16114
rect 3516 16050 3568 16056
rect 3700 16050 3752 16056
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3528 15638 3556 15914
rect 3712 15706 3740 16050
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3804 14890 3832 15098
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3712 14278 3740 14826
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12209 3464 12582
rect 3422 12200 3478 12209
rect 3422 12135 3478 12144
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3252 11558 3280 11834
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11218 3280 11494
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3344 11014 3372 11562
rect 3620 11354 3648 11698
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3422 11248 3478 11257
rect 3422 11183 3478 11192
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8430 3188 8774
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 8022 3188 8366
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3068 6390 3096 6802
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2780 5908 2832 5914
rect 2832 5868 3004 5896
rect 2780 5850 2832 5856
rect 2976 5710 3004 5868
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3160 5166 3188 6054
rect 3252 5846 3280 6258
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2700 5001 2728 5034
rect 3344 5030 3372 10950
rect 3436 10606 3464 11183
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10266 3556 10406
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3436 9382 3464 9454
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 7206 3464 9318
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 5166 3464 7142
rect 3514 5264 3570 5273
rect 3514 5199 3570 5208
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3332 5024 3384 5030
rect 2686 4992 2742 5001
rect 3332 4966 3384 4972
rect 2686 4927 2742 4936
rect 2780 4684 2832 4690
rect 2608 4644 2780 4672
rect 2780 4626 2832 4632
rect 2792 3738 2820 4626
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3436 3670 3464 3878
rect 3528 3738 3556 5199
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 3126 3096 3402
rect 3436 3126 3464 3606
rect 3528 3534 3556 3674
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3712 3194 3740 14214
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3804 12986 3832 13398
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12170 3832 12582
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3790 10296 3846 10305
rect 3896 10266 3924 17478
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3988 16182 4016 16594
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4356 15026 4384 15914
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3790 10231 3846 10240
rect 3884 10260 3936 10266
rect 3804 6866 3832 10231
rect 3884 10202 3936 10208
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3896 9042 3924 9318
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3896 8090 3924 8978
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3896 4826 3924 5102
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 3738 3832 4626
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3896 3670 3924 4422
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1872 2310 1900 2450
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1122 54 1440 82
rect 1872 82 1900 2246
rect 1950 82 2006 480
rect 1872 54 2006 82
rect 2516 82 2544 2858
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2608 1057 2636 2518
rect 2594 1048 2650 1057
rect 2594 983 2650 992
rect 2778 82 2834 480
rect 2516 54 2834 82
rect 3160 82 3188 2790
rect 3436 2106 3464 3062
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3514 2544 3570 2553
rect 3514 2479 3570 2488
rect 3528 2446 3556 2479
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3620 513 3648 2790
rect 3882 2680 3938 2689
rect 3988 2650 4016 14214
rect 4080 13190 4108 14350
rect 4356 13802 4384 14554
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4172 12782 4200 13359
rect 4448 13326 4476 16662
rect 4252 13320 4304 13326
rect 4436 13320 4488 13326
rect 4304 13280 4384 13308
rect 4252 13262 4304 13268
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12374 4292 12650
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4172 11558 4200 12174
rect 4264 11898 4292 12310
rect 4356 12102 4384 13280
rect 4436 13262 4488 13268
rect 4816 12374 4844 19178
rect 4908 17882 4936 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5000 16998 5028 17682
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 14618 5028 16934
rect 5184 15094 5212 17614
rect 5276 17202 5304 18022
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5552 17270 5580 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 16794 5304 17138
rect 6012 17066 6040 18158
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 6000 17060 6052 17066
rect 6000 17002 6052 17008
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5368 16726 5396 17002
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16114 6040 17002
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5276 15706 5304 15914
rect 6288 15910 6316 16594
rect 6564 16561 6592 16594
rect 6550 16552 6606 16561
rect 7576 16522 7604 17070
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 6550 16487 6606 16496
rect 7564 16516 7616 16522
rect 6564 16250 6592 16487
rect 7564 16458 7616 16464
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 7576 16114 7604 16458
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7840 15972 7892 15978
rect 7944 15960 7972 16390
rect 7892 15932 7972 15960
rect 7840 15914 7892 15920
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15162 5488 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5276 14414 5304 14826
rect 5368 14618 5396 14826
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 6288 14550 6316 15846
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6656 15026 6684 15574
rect 6840 15502 6868 15846
rect 7944 15570 7972 15932
rect 8036 15910 8064 16662
rect 8128 16590 8156 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 16250 8156 16526
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8588 16046 8616 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8036 15638 8064 15846
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6840 15094 6868 15438
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7208 14618 7236 14894
rect 8404 14822 8432 15846
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13734 5580 14350
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6472 14074 6500 14554
rect 8404 14550 8432 14758
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8404 14074 8432 14486
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5184 13462 5212 13670
rect 5552 13530 5580 13670
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5828 13462 5856 13670
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5816 13456 5868 13462
rect 6472 13444 6500 14010
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 6656 13734 6684 13806
rect 8404 13734 8432 13806
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 6552 13456 6604 13462
rect 6472 13416 6552 13444
rect 5816 13398 5868 13404
rect 6552 13398 6604 13404
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12850 6040 13262
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5276 12442 5304 12718
rect 6564 12646 6592 13398
rect 6656 13326 6684 13670
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4816 11744 4844 12310
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 4896 11756 4948 11762
rect 4816 11716 4896 11744
rect 4896 11698 4948 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4908 11354 4936 11562
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4540 9926 4568 10406
rect 4816 10266 4844 11086
rect 5184 10538 5212 11290
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 5276 10130 5304 11698
rect 6012 11626 6040 12310
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6012 11354 6040 11562
rect 6564 11558 6592 12582
rect 6656 12306 6684 13262
rect 6932 13190 6960 13670
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12782 7052 13126
rect 7668 12850 7696 13330
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7944 12986 7972 13194
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6656 11762 6684 12242
rect 6748 11898 6776 12242
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6564 11286 6592 11494
rect 6748 11354 6776 11834
rect 6840 11762 6868 12378
rect 6920 12368 6972 12374
rect 7024 12356 7052 12718
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6972 12328 7052 12356
rect 6920 12310 6972 12316
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6642 11248 6698 11257
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5828 10130 5856 10610
rect 6012 10470 6040 10678
rect 6564 10538 6592 11222
rect 6642 11183 6698 11192
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 8906 4200 9454
rect 4540 9110 4568 9862
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4540 8294 4568 9046
rect 5092 8906 5120 10066
rect 5276 9722 5304 10066
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5368 9178 5396 10066
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4908 8566 4936 8842
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5000 8634 5028 8774
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5092 8498 5120 8842
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4080 6322 4108 8026
rect 4540 8022 4568 8230
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4264 6798 4292 7278
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4632 6730 4660 7890
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4724 7546 4752 7822
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4724 7449 4752 7482
rect 5184 7478 5212 8774
rect 5276 8362 5304 8910
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 7478 5304 8298
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5172 7472 5224 7478
rect 4710 7440 4766 7449
rect 5172 7414 5224 7420
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 4710 7375 4766 7384
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4448 5914 4476 6598
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5302 4200 5714
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4632 5166 4660 6666
rect 4724 5778 4752 7375
rect 5264 7268 5316 7274
rect 5368 7256 5396 8026
rect 5460 7546 5488 9930
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9518 6040 10406
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6288 8634 6316 9046
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8634 6592 8910
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8362 6684 11183
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6748 10266 6776 10474
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9654 6868 9998
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5460 7274 5488 7482
rect 5552 7410 5580 7686
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5316 7228 5396 7256
rect 5448 7268 5500 7274
rect 5264 7210 5316 7216
rect 5448 7210 5500 7216
rect 6196 7206 6224 7958
rect 6656 7818 6684 8298
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 7024 7274 7052 7890
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6254 4936 6598
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4802 5808 4858 5817
rect 4712 5772 4764 5778
rect 4802 5743 4858 5752
rect 4712 5714 4764 5720
rect 4620 5160 4672 5166
rect 4816 5137 4844 5743
rect 4620 5102 4672 5108
rect 4802 5128 4858 5137
rect 4908 5098 4936 6190
rect 5460 6186 5488 6734
rect 5552 6458 5580 6938
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5914 5488 6122
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 6012 5846 6040 7142
rect 6196 6934 6224 7142
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6196 6118 6224 6870
rect 6840 6662 6868 7142
rect 7024 7002 7052 7210
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6361 6868 6598
rect 7116 6458 7144 12378
rect 7668 12102 7696 12786
rect 8404 12782 8432 13670
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8024 12164 8076 12170
rect 8024 12106 8076 12112
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7668 10810 7696 12038
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 9722 7420 10542
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7576 9586 7604 10610
rect 7852 10470 7880 12038
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 8498 7512 9454
rect 7668 9178 7696 9998
rect 7852 9926 7880 10406
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9654 7880 9862
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7852 8566 7880 9590
rect 7944 9178 7972 10066
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7576 7750 7604 8502
rect 7944 8362 7972 9114
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7576 7546 7604 7686
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7392 6458 7420 6870
rect 7576 6866 7604 7482
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7944 6662 7972 7686
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5276 5166 5304 5510
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 4802 5063 4858 5072
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 3670 4292 4422
rect 4540 3942 4568 4694
rect 5276 4690 5304 4966
rect 5368 4826 5396 5714
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4802 4176 4858 4185
rect 5552 4154 5580 5306
rect 6012 4826 6040 5782
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6196 4758 6224 6054
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5552 4126 5672 4154
rect 4802 4111 4858 4120
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4816 3670 4844 4111
rect 5644 4078 5672 4126
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 3738 5672 4014
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 4252 3664 4304 3670
rect 4804 3664 4856 3670
rect 4252 3606 4304 3612
rect 4724 3624 4804 3652
rect 4264 2689 4292 3606
rect 4250 2680 4306 2689
rect 3882 2615 3938 2624
rect 3976 2644 4028 2650
rect 3896 2514 3924 2615
rect 4250 2615 4306 2624
rect 3976 2586 4028 2592
rect 4724 2582 4752 3624
rect 4804 3606 4856 3612
rect 5920 3534 5948 3946
rect 6196 3942 6224 4694
rect 6656 4690 6684 5850
rect 6840 5710 6868 6054
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 7208 5302 7236 5714
rect 7484 5370 7512 5714
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6656 4282 6684 4626
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6932 4146 6960 4966
rect 7116 4690 7144 5102
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3670 6224 3878
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6090 3224 6146 3233
rect 6090 3159 6146 3168
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 3606 504 3662 513
rect 3514 82 3570 480
rect 3606 439 3662 448
rect 3160 54 3570 82
rect 386 0 442 54
rect 1122 0 1178 54
rect 1950 0 2006 54
rect 2778 0 2834 54
rect 3514 0 3570 54
rect 4342 82 4398 480
rect 4632 82 4660 1974
rect 4342 54 4660 82
rect 4816 82 4844 2790
rect 5368 649 5396 2858
rect 6104 2689 6132 3159
rect 6196 3058 6224 3606
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6090 2680 6146 2689
rect 6288 2650 6316 3470
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6932 3058 6960 3402
rect 7012 3392 7064 3398
rect 7208 3369 7236 4422
rect 7746 4312 7802 4321
rect 7746 4247 7802 4256
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7668 3738 7696 3946
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7012 3334 7064 3340
rect 7194 3360 7250 3369
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7024 2922 7052 3334
rect 7194 3295 7250 3304
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 6734 2680 6790 2689
rect 6090 2615 6146 2624
rect 6276 2644 6328 2650
rect 6734 2615 6790 2624
rect 6276 2586 6328 2592
rect 6748 2582 6776 2615
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 5460 1057 5488 2518
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 5446 1048 5502 1057
rect 5446 983 5502 992
rect 5354 640 5410 649
rect 5354 575 5410 584
rect 5170 82 5226 480
rect 4816 54 5226 82
rect 5552 82 5580 2314
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6656 1057 6684 2042
rect 7024 1737 7052 2858
rect 7116 2446 7144 2858
rect 7208 2689 7236 3295
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7194 2680 7250 2689
rect 7194 2615 7250 2624
rect 7208 2582 7236 2615
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7668 2446 7696 2790
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7010 1728 7066 1737
rect 7010 1663 7066 1672
rect 6642 1048 6698 1057
rect 6642 983 6698 992
rect 5906 82 5962 480
rect 5552 54 5962 82
rect 4342 0 4398 54
rect 5170 0 5226 54
rect 5906 0 5962 54
rect 6734 128 6790 480
rect 6734 76 6736 128
rect 6788 76 6790 128
rect 6734 0 6790 76
rect 7562 82 7618 480
rect 7760 82 7788 4247
rect 7944 3534 7972 4762
rect 8036 4154 8064 12106
rect 8128 11898 8156 12242
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8496 11558 8524 14214
rect 8588 13734 8616 15982
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15570 9352 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8680 12714 8708 14894
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 14550 9904 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13870 9076 14214
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9048 12850 9076 13806
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13258 9168 13738
rect 9692 13546 9720 14010
rect 9876 14006 9904 14486
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9508 13518 9720 13546
rect 9784 13530 9812 13942
rect 10888 13870 10916 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 9772 13524 9824 13530
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 9140 11694 9168 13194
rect 9324 12782 9352 13398
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8404 10606 8432 11086
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8496 10470 8524 11018
rect 8588 10742 8616 11154
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8864 10606 8892 11290
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8404 9518 8432 10202
rect 8864 10198 8892 10542
rect 8852 10192 8904 10198
rect 8758 10160 8814 10169
rect 8852 10134 8904 10140
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8758 10095 8814 10104
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 9654 8708 9862
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8680 9042 8708 9590
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8680 8634 8708 8978
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8390 8528 8446 8537
rect 8390 8463 8446 8472
rect 8668 8492 8720 8498
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7002 8156 7822
rect 8312 7274 8340 8298
rect 8404 8090 8432 8463
rect 8668 8434 8720 8440
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8680 7857 8708 8434
rect 8666 7848 8722 7857
rect 8588 7806 8666 7834
rect 8390 7712 8446 7721
rect 8390 7647 8446 7656
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5166 8156 6054
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8312 4690 8340 5034
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4282 8340 4626
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8036 4126 8340 4154
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 2650 7972 3470
rect 8036 3126 8064 3606
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8312 2650 8340 4126
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7562 54 7788 82
rect 8298 82 8354 480
rect 8404 82 8432 7647
rect 8588 6798 8616 7806
rect 8666 7783 8722 7792
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7478 8708 7686
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6866 8708 7278
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 6254 8616 6734
rect 8680 6730 8708 6802
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8680 5914 8708 6258
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 3194 8524 5646
rect 8772 5001 8800 10095
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8864 8294 8892 8502
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 6662 8892 8230
rect 8956 7954 8984 10134
rect 9048 10062 9076 11494
rect 9140 11014 9168 11630
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9586 9076 9998
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 8022 9076 9522
rect 9140 8906 9168 10950
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 9048 7886 9076 7958
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 5574 8892 6598
rect 9048 5846 9076 7142
rect 9232 7002 9260 11562
rect 9324 11082 9352 12718
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9416 10674 9444 13126
rect 9508 12850 9536 13518
rect 9772 13466 9824 13472
rect 10704 13462 10732 13738
rect 10888 13530 10916 13806
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9680 13252 9732 13258
rect 9732 13212 9812 13240
rect 9680 13194 9732 13200
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9496 12164 9548 12170
rect 9600 12152 9628 13126
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12374 9720 12718
rect 9784 12646 9812 13212
rect 9876 12986 9904 13330
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9864 12980 9916 12986
rect 9916 12940 9996 12968
rect 9864 12922 9916 12928
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9548 12124 9628 12152
rect 9496 12106 9548 12112
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10606 9536 12106
rect 9692 11694 9720 12310
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9692 11354 9720 11630
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9324 7002 9352 10202
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 8634 9444 10066
rect 9508 9926 9536 10542
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9722 9536 9862
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9416 7954 9444 8570
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9232 6186 9260 6938
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9232 5846 9260 6122
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8758 4992 8814 5001
rect 8758 4927 8814 4936
rect 8864 4826 8892 5510
rect 9232 4826 9260 5782
rect 9508 5778 9536 6394
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8680 4282 8708 4558
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 3670 9076 3878
rect 9140 3738 9168 4014
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8588 3126 8616 3334
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8588 2922 8616 3062
rect 9416 3058 9444 3334
rect 9508 3194 9536 5034
rect 9600 4729 9628 11086
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9042 9720 9998
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8498 9720 8978
rect 9784 8634 9812 12582
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 9110 9904 12174
rect 9968 10130 9996 12940
rect 10152 12102 10180 13126
rect 10704 12714 10732 13398
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 11072 12442 11100 12718
rect 11900 12714 11928 13330
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12442 11192 12582
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10060 11558 10088 11766
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9784 7954 9812 8570
rect 9956 8560 10008 8566
rect 10060 8548 10088 11494
rect 10152 11336 10180 12038
rect 10520 11694 10548 12310
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11762 10916 12038
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10508 11688 10560 11694
rect 11152 11688 11204 11694
rect 10560 11648 10824 11676
rect 10508 11630 10560 11636
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10152 11308 10272 11336
rect 10244 10742 10272 11308
rect 10796 11218 10824 11648
rect 11152 11630 11204 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10784 10736 10836 10742
rect 10784 10678 10836 10684
rect 10152 10130 10180 10678
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 10474
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 9382 10180 10066
rect 10796 9926 10824 10678
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10008 8520 10088 8548
rect 9956 8502 10008 8508
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9784 7342 9812 7890
rect 10060 7449 10088 8366
rect 10046 7440 10102 7449
rect 10046 7375 10102 7384
rect 10152 7342 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7478 10272 7686
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 9772 7336 9824 7342
rect 10140 7336 10192 7342
rect 9824 7296 9904 7324
rect 9772 7278 9824 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6390 9720 7142
rect 9876 6866 9904 7296
rect 10140 7278 10192 7284
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9876 6186 9904 6802
rect 10060 6798 10088 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6254 10088 6734
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10152 6390 10180 6598
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5370 9812 6054
rect 10060 5710 10088 6190
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 5370 10088 5646
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10152 5166 10180 5510
rect 10704 5166 10732 7210
rect 10796 6662 10824 7482
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6458 10824 6598
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4826 10732 5102
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10140 4752 10192 4758
rect 9586 4720 9642 4729
rect 10140 4694 10192 4700
rect 9586 4655 9642 4664
rect 9600 4282 9628 4655
rect 9956 4616 10008 4622
rect 9678 4584 9734 4593
rect 9956 4558 10008 4564
rect 9678 4519 9734 4528
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9692 3466 9720 4519
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9784 3194 9812 3946
rect 9968 3466 9996 4558
rect 10152 3942 10180 4694
rect 10704 4214 10732 4762
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10060 3670 10088 3878
rect 10048 3664 10100 3670
rect 10152 3641 10180 3878
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10048 3606 10100 3612
rect 10138 3632 10194 3641
rect 10138 3567 10194 3576
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 10888 3398 10916 11018
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8588 2417 8616 2858
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2650 8800 2790
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8574 2408 8630 2417
rect 8574 2343 8630 2352
rect 8850 2408 8906 2417
rect 8850 2343 8906 2352
rect 8864 2310 8892 2343
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8956 2038 8984 2450
rect 9600 2446 9628 3062
rect 9784 2990 9812 3130
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9588 2440 9640 2446
rect 9968 2417 9996 2518
rect 10152 2446 10180 2858
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10888 2582 10916 2790
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10140 2440 10192 2446
rect 9588 2382 9640 2388
rect 9954 2408 10010 2417
rect 10140 2382 10192 2388
rect 9954 2343 10010 2352
rect 8944 2032 8996 2038
rect 8944 1974 8996 1980
rect 8298 54 8432 82
rect 9126 60 9182 480
rect 7562 0 7618 54
rect 8298 0 8354 54
rect 9126 8 9128 60
rect 9180 8 9182 60
rect 9126 0 9182 8
rect 9954 128 10010 480
rect 9954 76 9956 128
rect 10008 76 10010 128
rect 9954 0 10010 76
rect 10690 96 10746 480
rect 10980 66 11008 10678
rect 11072 7818 11100 11494
rect 11164 10266 11192 11630
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11164 9450 11192 10202
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 8906 11192 9386
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 7954 11192 8570
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 7546 11100 7754
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11256 7478 11284 11562
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11440 10810 11468 11086
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10470 11560 11154
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10198 11560 10406
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11440 9722 11468 10066
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 8430 11376 9114
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11348 8022 11376 8366
rect 11440 8294 11468 8978
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 8022 11468 8230
rect 11532 8090 11560 10134
rect 11624 9518 11652 11494
rect 11716 11354 11744 12242
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11716 11257 11744 11290
rect 11702 11248 11758 11257
rect 11702 11183 11758 11192
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11624 7954 11652 9454
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11624 7274 11652 7890
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11164 4154 11192 6870
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11256 5846 11284 6802
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11520 6656 11572 6662
rect 11440 6616 11520 6644
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11348 5302 11376 6394
rect 11440 6118 11468 6616
rect 11520 6598 11572 6604
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5914 11468 6054
rect 11624 5914 11652 6734
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11072 4146 11192 4154
rect 11060 4140 11192 4146
rect 11112 4126 11192 4140
rect 11060 4082 11112 4088
rect 11150 4040 11206 4049
rect 11150 3975 11206 3984
rect 11164 2650 11192 3975
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11256 3058 11284 3606
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 2961 11284 2994
rect 11242 2952 11298 2961
rect 11242 2887 11298 2896
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11164 2378 11192 2586
rect 11348 2553 11376 4558
rect 11440 4486 11468 5850
rect 11716 5778 11744 11086
rect 11808 10538 11836 12242
rect 12268 12209 12296 13262
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12348 12232 12400 12238
rect 12254 12200 12310 12209
rect 12348 12174 12400 12180
rect 12254 12135 12310 12144
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11900 9994 11928 11086
rect 11992 10538 12020 11698
rect 12360 11354 12388 12174
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11808 8906 11836 9862
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 4826 11744 5714
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11624 2854 11652 3606
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11334 2544 11390 2553
rect 11334 2479 11390 2488
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11624 921 11652 2790
rect 11610 912 11666 921
rect 11610 847 11666 856
rect 11518 82 11574 480
rect 11808 82 11836 7686
rect 11900 7546 11928 7822
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11900 6798 11928 7482
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11992 6390 12020 9998
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 12084 7206 12112 7958
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 4758 11928 6054
rect 12084 5953 12112 7142
rect 12070 5944 12126 5953
rect 12070 5879 12126 5888
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5030 12020 5782
rect 12176 5234 12204 9658
rect 12268 9382 12296 10066
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9518 12572 9862
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 6798 12296 9318
rect 12360 8838 12388 9454
rect 12544 9178 12572 9454
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 7313 12388 8774
rect 12452 8566 12480 8910
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8634 12572 8774
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12452 8090 12480 8502
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12346 7304 12402 7313
rect 12346 7239 12402 7248
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12268 5137 12296 6734
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12254 5128 12310 5137
rect 12164 5092 12216 5098
rect 12254 5063 12310 5072
rect 12164 5034 12216 5040
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11992 4010 12020 4966
rect 12176 4078 12204 5034
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 11900 3913 11928 3946
rect 11886 3904 11942 3913
rect 11886 3839 11942 3848
rect 12360 3738 12388 6666
rect 12544 6066 12572 7210
rect 12636 6186 12664 9522
rect 12728 7002 12756 12582
rect 12912 12345 12940 12718
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 12898 12336 12954 12345
rect 12898 12271 12954 12280
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 11824 12952 11830
rect 12820 11784 12900 11812
rect 12820 9178 12848 11784
rect 12900 11766 12952 11772
rect 13004 11762 13032 12174
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12820 7970 12848 9114
rect 12912 9110 12940 10406
rect 13004 9110 13032 11698
rect 13096 11694 13124 12038
rect 13188 11830 13216 12242
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11286 13124 11494
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13096 9722 13124 10066
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9568 13216 11630
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13096 9540 13216 9568
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12912 8090 12940 9046
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12820 7942 12940 7970
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12728 6322 12756 6938
rect 12806 6760 12862 6769
rect 12806 6695 12862 6704
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12544 6038 12756 6066
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12544 5234 12572 5714
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12636 5098 12664 5578
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12452 4146 12480 4762
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 2854 11928 3470
rect 12636 3398 12664 4694
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11900 2650 11928 2790
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12636 1329 12664 3334
rect 12728 2106 12756 6038
rect 12820 3126 12848 6695
rect 12912 4758 12940 7942
rect 13004 6322 13032 8434
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 12912 2922 12940 3334
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12820 2310 12848 2858
rect 13004 2689 13032 3470
rect 12990 2680 13046 2689
rect 12990 2615 13046 2624
rect 13004 2446 13032 2615
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12820 1601 12848 2246
rect 12806 1592 12862 1601
rect 12806 1527 12862 1536
rect 12622 1320 12678 1329
rect 12622 1255 12678 1264
rect 13096 626 13124 9540
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8498 13216 9386
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 8090 13216 8230
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13188 7410 13216 8026
rect 13280 7886 13308 11562
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 8634 13400 10542
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13372 8022 13400 8570
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13188 7206 13216 7346
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6866 13216 7142
rect 13280 7002 13308 7822
rect 13372 7546 13400 7958
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13464 7018 13492 12174
rect 13832 11898 13860 12242
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13556 10169 13584 11018
rect 13648 10810 13676 11154
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13648 10266 13676 10746
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13542 10160 13598 10169
rect 13542 10095 13598 10104
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13372 6990 13492 7018
rect 13176 6860 13228 6866
rect 13228 6820 13308 6848
rect 13176 6802 13228 6808
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13188 6458 13216 6666
rect 13280 6458 13308 6820
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13188 5846 13216 6122
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 13188 5234 13216 5782
rect 13372 5778 13400 6990
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13464 5914 13492 6870
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13464 5710 13492 5850
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13464 4758 13492 5646
rect 13556 5574 13584 9998
rect 13648 9654 13676 10066
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8022 13676 8910
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13740 7750 13768 11834
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 14108 10742 14136 11154
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13832 8906 13860 9114
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13924 7857 13952 9046
rect 14016 8838 14044 9386
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 13910 7848 13966 7857
rect 13910 7783 13966 7792
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13634 7304 13690 7313
rect 13634 7239 13690 7248
rect 13648 5778 13676 7239
rect 13726 7168 13782 7177
rect 13726 7103 13782 7112
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13648 5302 13676 5714
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13174 4448 13230 4457
rect 13174 4383 13230 4392
rect 13188 3670 13216 4383
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3670 13400 3878
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13188 2650 13216 3606
rect 13464 3534 13492 4490
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3058 13492 3334
rect 13634 3088 13690 3097
rect 13452 3052 13504 3058
rect 13740 3074 13768 7103
rect 13924 5302 13952 7783
rect 14016 5642 14044 8774
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14200 8090 14228 8366
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 14108 5166 14136 7142
rect 14292 6934 14320 8298
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 14280 6928 14332 6934
rect 14200 6876 14280 6882
rect 14200 6870 14332 6876
rect 14200 6854 14320 6870
rect 14200 6254 14228 6854
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4729 14228 4966
rect 14186 4720 14242 4729
rect 14004 4684 14056 4690
rect 14186 4655 14242 4664
rect 14004 4626 14056 4632
rect 14016 3942 14044 4626
rect 14200 4622 14228 4655
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14108 4214 14136 4558
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13690 3046 13768 3074
rect 13634 3023 13690 3032
rect 13452 2994 13504 3000
rect 13832 2854 13860 3606
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13832 2553 13860 2790
rect 13818 2544 13874 2553
rect 13818 2479 13874 2488
rect 14016 2038 14044 3878
rect 14200 3194 14228 3946
rect 14292 3738 14320 6734
rect 14384 6322 14412 8230
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14384 4146 14412 5646
rect 14476 4593 14504 10406
rect 14568 7721 14596 10610
rect 15488 10538 15516 11154
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 14752 8809 14780 10474
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14738 8664 14794 8673
rect 14956 8656 15252 8676
rect 14738 8599 14794 8608
rect 14752 8498 14780 8599
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14554 7712 14610 7721
rect 14554 7647 14610 7656
rect 14660 6186 14688 8026
rect 15396 8022 15424 9998
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15488 9110 15516 9454
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15488 8634 15516 9046
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7478 15424 7958
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 14832 7336 14884 7342
rect 14830 7304 14832 7313
rect 14884 7304 14886 7313
rect 14830 7239 14886 7248
rect 14844 7206 14872 7239
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14844 6458 14872 7142
rect 15304 6798 15332 7142
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6458 15332 6734
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14752 4690 14780 6326
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 4758 14872 6190
rect 15120 5914 15148 6258
rect 15488 6186 15516 8298
rect 15580 8022 15608 9386
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15580 7546 15608 7958
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15200 5296 15252 5302
rect 15304 5284 15332 5714
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5370 15516 5510
rect 15672 5409 15700 10406
rect 15658 5400 15714 5409
rect 15476 5364 15528 5370
rect 15658 5335 15714 5344
rect 15476 5306 15528 5312
rect 15252 5256 15332 5284
rect 15566 5264 15622 5273
rect 15200 5238 15252 5244
rect 15384 5228 15436 5234
rect 15566 5199 15622 5208
rect 15384 5170 15436 5176
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14462 4584 14518 4593
rect 14462 4519 14518 4528
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14200 2922 14228 3130
rect 14292 3058 14320 3674
rect 14476 3194 14504 3878
rect 14568 3369 14596 4490
rect 14752 3738 14780 4626
rect 15396 4486 15424 5170
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15292 3664 15344 3670
rect 15396 3641 15424 4422
rect 15292 3606 15344 3612
rect 15382 3632 15438 3641
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14738 2272 14794 2281
rect 14738 2207 14794 2216
rect 14004 2032 14056 2038
rect 13818 2000 13874 2009
rect 14004 1974 14056 1980
rect 14752 1970 14780 2207
rect 13818 1935 13874 1944
rect 14740 1964 14792 1970
rect 13096 598 13216 626
rect 10690 0 10746 40
rect 10968 60 11020 66
rect 10968 2 11020 8
rect 11518 54 11836 82
rect 12346 82 12402 480
rect 12530 368 12586 377
rect 12530 303 12586 312
rect 12544 82 12572 303
rect 12346 54 12572 82
rect 13082 82 13138 480
rect 13188 82 13216 598
rect 13082 54 13216 82
rect 13832 82 13860 1935
rect 14740 1906 14792 1912
rect 13910 82 13966 480
rect 14004 196 14056 202
rect 14004 138 14056 144
rect 14016 105 14044 138
rect 13832 54 13966 82
rect 11518 0 11574 54
rect 12346 0 12402 54
rect 13082 0 13138 54
rect 13910 0 13966 54
rect 14002 96 14058 105
rect 14002 31 14058 40
rect 14738 82 14794 480
rect 14844 82 14872 3402
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15304 2650 15332 3606
rect 15382 3567 15438 3576
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15580 2514 15608 5199
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14738 54 14872 82
rect 15566 82 15622 480
rect 15764 82 15792 4966
rect 15856 4593 15884 10542
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9382 16528 10066
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 18418 9888 18474 9897
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 9081 16528 9318
rect 16486 9072 16542 9081
rect 16486 9007 16542 9016
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 7886 16068 8910
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16040 6905 16068 7822
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16026 6896 16082 6905
rect 16132 6866 16160 7210
rect 16224 7002 16252 8366
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16026 6831 16082 6840
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5234 15976 6122
rect 16224 5914 16252 6938
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16224 5098 16252 5850
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4758 16160 4966
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 15842 4584 15898 4593
rect 15842 4519 15898 4528
rect 15948 4010 15976 4694
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16040 2378 16068 2926
rect 16132 2825 16160 3839
rect 16224 3670 16252 4626
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16316 2922 16344 5510
rect 16396 5296 16448 5302
rect 16396 5238 16448 5244
rect 16408 4690 16436 5238
rect 16500 4758 16528 5646
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16592 4154 16620 9862
rect 18418 9823 18474 9832
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16960 8634 16988 8978
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17144 8537 17172 8774
rect 17130 8528 17186 8537
rect 17130 8463 17186 8472
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7342 16988 7686
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16776 6458 16804 6802
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16960 6322 16988 6734
rect 17144 6730 17172 7142
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17420 6118 17448 6938
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16868 5030 16896 5850
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16500 4126 16620 4154
rect 16500 3534 16528 4126
rect 17052 3942 17080 4626
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17328 4282 17356 4422
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17512 4185 17540 8910
rect 18248 8634 18276 9386
rect 18432 9042 18460 9823
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18432 8634 18460 8978
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 5846 17908 7142
rect 17972 7002 18000 7890
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17972 6458 18000 6938
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 6118 18000 6394
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 18064 5370 18092 7210
rect 18156 6934 18184 7822
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5914 18184 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4214 17632 4966
rect 17592 4208 17644 4214
rect 17498 4176 17554 4185
rect 17592 4150 17644 4156
rect 17498 4111 17554 4120
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 16396 3528 16448 3534
rect 16394 3496 16396 3505
rect 16488 3528 16540 3534
rect 16448 3496 16450 3505
rect 16488 3470 16540 3476
rect 16394 3431 16450 3440
rect 16408 3058 16436 3431
rect 16486 3360 16542 3369
rect 16486 3295 16542 3304
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16118 2816 16174 2825
rect 16118 2751 16174 2760
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 15566 54 15792 82
rect 16132 82 16160 2751
rect 16500 2582 16528 3295
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16960 2446 16988 3878
rect 17052 3466 17080 3878
rect 17420 3738 17448 3878
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 3194 17080 3402
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17144 2650 17172 3470
rect 17236 3126 17264 3606
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17420 3058 17448 3674
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17406 2680 17462 2689
rect 17132 2644 17184 2650
rect 17406 2615 17462 2624
rect 17132 2586 17184 2592
rect 17420 2514 17448 2615
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 1193 16436 2246
rect 16856 2032 16908 2038
rect 16856 1974 16908 1980
rect 16394 1184 16450 1193
rect 16394 1119 16450 1128
rect 16302 82 16358 480
rect 16132 54 16358 82
rect 16868 82 16896 1974
rect 17130 82 17186 480
rect 16868 54 17186 82
rect 17696 82 17724 5170
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 3534 17816 5102
rect 18064 5030 18092 5306
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17972 4010 18000 4150
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17972 3466 18000 3946
rect 18064 3738 18092 4014
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 18156 2582 18184 4014
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 17958 82 18014 480
rect 18248 134 18276 7278
rect 18420 5704 18472 5710
rect 18616 5692 18644 12650
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7206 18736 7890
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 5817 18736 7142
rect 18788 6724 18840 6730
rect 18788 6666 18840 6672
rect 18800 6322 18828 6666
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18616 5664 18828 5692
rect 18420 5646 18472 5652
rect 18432 5234 18460 5646
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18340 649 18368 4966
rect 18432 4758 18460 5170
rect 18524 4758 18552 5578
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18512 4752 18564 4758
rect 18512 4694 18564 4700
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 2446 18460 3334
rect 18524 2582 18552 3946
rect 18616 2922 18644 4218
rect 18708 4146 18736 4558
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18800 3126 18828 5664
rect 18892 3942 18920 8774
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 21822 7984 21878 7993
rect 21822 7919 21878 7928
rect 23848 7948 23900 7954
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19430 7168 19486 7177
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19076 6458 19104 6870
rect 19168 6662 19196 7142
rect 19430 7103 19486 7112
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19260 6390 19288 6598
rect 19352 6458 19380 6734
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19444 6322 19472 7103
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18984 3670 19012 6122
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5914 20024 6190
rect 20824 6118 20852 6802
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19614 5808 19670 5817
rect 19076 5370 19104 5782
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19168 5234 19196 5714
rect 19536 5273 19564 5782
rect 19614 5743 19670 5752
rect 19522 5264 19578 5273
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19340 5228 19392 5234
rect 19522 5199 19578 5208
rect 19340 5170 19392 5176
rect 19062 5128 19118 5137
rect 19062 5063 19118 5072
rect 19076 4690 19104 5063
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 19076 4154 19104 4626
rect 19260 4554 19288 4966
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19352 4162 19380 5170
rect 19628 5148 19656 5743
rect 19076 4126 19196 4154
rect 19168 3738 19196 4126
rect 19306 4134 19380 4162
rect 19536 5120 19656 5148
rect 19306 4026 19334 4134
rect 19260 3998 19334 4026
rect 19260 3777 19288 3998
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19246 3768 19302 3777
rect 19156 3732 19208 3738
rect 19246 3703 19302 3712
rect 19156 3674 19208 3680
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 19248 3664 19300 3670
rect 19248 3606 19300 3612
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18708 2582 18736 3062
rect 18892 2650 18920 3470
rect 19168 3058 19196 3470
rect 19260 3194 19288 3606
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 19260 2689 19288 2994
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 19352 2825 19380 2858
rect 19338 2816 19394 2825
rect 19338 2751 19394 2760
rect 19246 2680 19302 2689
rect 18880 2644 18932 2650
rect 19246 2615 19302 2624
rect 18880 2586 18932 2592
rect 18512 2576 18564 2582
rect 18512 2518 18564 2524
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 19260 2514 19288 2615
rect 19444 2514 19472 3878
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18432 2310 18460 2382
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18420 2100 18472 2106
rect 18420 2042 18472 2048
rect 18326 640 18382 649
rect 18326 575 18382 584
rect 17696 54 18014 82
rect 18236 128 18288 134
rect 18236 70 18288 76
rect 18432 82 18460 2042
rect 19536 626 19564 5120
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4282 20024 5850
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 2990 19840 3334
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19536 598 19656 626
rect 18694 82 18750 480
rect 18432 54 18750 82
rect 14738 0 14794 54
rect 15566 0 15622 54
rect 16302 0 16358 54
rect 17130 0 17186 54
rect 17958 0 18014 54
rect 18694 0 18750 54
rect 19522 82 19578 480
rect 19628 82 19656 598
rect 19522 54 19656 82
rect 20088 82 20116 3402
rect 20272 921 20300 4558
rect 20456 3777 20484 6054
rect 20916 5778 20944 7278
rect 21088 7200 21140 7206
rect 21640 7200 21692 7206
rect 21088 7142 21140 7148
rect 21546 7168 21602 7177
rect 21100 6769 21128 7142
rect 21640 7142 21692 7148
rect 21546 7103 21602 7112
rect 21086 6760 21142 6769
rect 21086 6695 21142 6704
rect 21560 6254 21588 7103
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21008 5370 21036 5714
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20442 3768 20498 3777
rect 20442 3703 20498 3712
rect 20548 3534 20576 4966
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20640 3369 20668 3878
rect 20626 3360 20682 3369
rect 20626 3295 20682 3304
rect 20732 2961 20760 5102
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 3942 20852 4626
rect 21100 4214 21128 6054
rect 21088 4208 21140 4214
rect 21088 4150 21140 4156
rect 21468 4049 21496 6122
rect 21454 4040 21510 4049
rect 21364 4004 21416 4010
rect 21454 3975 21510 3984
rect 21364 3946 21416 3952
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20824 3194 20852 3538
rect 20904 3528 20956 3534
rect 20904 3470 20956 3476
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20824 3097 20852 3130
rect 20810 3088 20866 3097
rect 20810 3023 20866 3032
rect 20718 2952 20774 2961
rect 20718 2887 20774 2896
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 20258 912 20314 921
rect 20258 847 20314 856
rect 20350 82 20406 480
rect 20088 54 20406 82
rect 20824 82 20852 2314
rect 20916 1737 20944 3470
rect 21100 1873 21128 3878
rect 21376 3233 21404 3946
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21362 3224 21418 3233
rect 21362 3159 21418 3168
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21086 1864 21142 1873
rect 21086 1799 21142 1808
rect 20902 1728 20958 1737
rect 20902 1663 20958 1672
rect 21192 1057 21220 2790
rect 21178 1048 21234 1057
rect 21178 983 21234 992
rect 21376 513 21404 2858
rect 21560 1601 21588 3878
rect 21652 2514 21680 7142
rect 21836 6866 21864 7919
rect 23848 7890 23900 7896
rect 23860 7206 23888 7890
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 21836 6458 21864 6802
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 22020 4690 22048 7142
rect 23860 6905 23888 7142
rect 23846 6896 23902 6905
rect 24228 6866 24256 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23846 6831 23902 6840
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 21744 1970 21772 4558
rect 22204 3058 22232 5034
rect 22480 5030 22508 5714
rect 23308 5098 23336 5714
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23296 5092 23348 5098
rect 23296 5034 23348 5040
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 23020 4684 23072 4690
rect 23020 4626 23072 4632
rect 22572 4282 22600 4626
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 23032 4010 23060 4626
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22296 2922 22324 3538
rect 22468 3528 22520 3534
rect 23032 3505 23060 3946
rect 22468 3470 22520 3476
rect 23018 3496 23074 3505
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22296 2825 22324 2858
rect 22282 2816 22338 2825
rect 22282 2751 22338 2760
rect 22480 2417 22508 3470
rect 23018 3431 23074 3440
rect 22466 2408 22522 2417
rect 22466 2343 22522 2352
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 21732 1964 21784 1970
rect 21732 1906 21784 1912
rect 21546 1592 21602 1601
rect 21546 1527 21602 1536
rect 21362 504 21418 513
rect 21086 82 21142 480
rect 21362 439 21418 448
rect 20824 54 21142 82
rect 19522 0 19578 54
rect 20350 0 20406 54
rect 21086 0 21142 54
rect 21914 82 21970 480
rect 22020 82 22048 2246
rect 21914 54 22048 82
rect 22664 82 22692 2314
rect 23308 785 23336 4694
rect 23400 2990 23428 5510
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 3641 23520 4966
rect 23860 4154 23888 6734
rect 24124 6724 24176 6730
rect 24124 6666 24176 6672
rect 24136 6254 24164 6666
rect 24228 6458 24256 6802
rect 26792 6656 26844 6662
rect 26792 6598 26844 6604
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23952 5166 23980 6054
rect 24766 5808 24822 5817
rect 24766 5743 24822 5752
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 24676 4480 24728 4486
rect 24122 4448 24178 4457
rect 24676 4422 24728 4428
rect 24122 4383 24178 4392
rect 24136 4282 24164 4383
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 23572 4140 23624 4146
rect 23860 4126 23980 4154
rect 23572 4082 23624 4088
rect 23478 3632 23534 3641
rect 23478 3567 23534 3576
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23294 776 23350 785
rect 23294 711 23350 720
rect 22742 82 22798 480
rect 22664 54 22798 82
rect 21914 0 21970 54
rect 22742 0 22798 54
rect 23478 82 23534 480
rect 23584 241 23612 4082
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23570 232 23626 241
rect 23570 167 23626 176
rect 23860 82 23888 2790
rect 23952 2514 23980 4126
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24044 1329 24072 3470
rect 24136 2009 24164 4014
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 3194 24256 3538
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24228 2553 24256 3130
rect 24214 2544 24270 2553
rect 24688 2514 24716 4422
rect 24780 3194 24808 5743
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24214 2479 24270 2488
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24122 2000 24178 2009
rect 24122 1935 24178 1944
rect 24030 1320 24086 1329
rect 24030 1255 24086 1264
rect 23478 54 23888 82
rect 24306 82 24362 480
rect 24688 82 24716 2246
rect 24872 105 24900 2926
rect 24306 54 24716 82
rect 24858 96 24914 105
rect 23478 0 23534 54
rect 24306 0 24362 54
rect 24964 82 24992 4490
rect 25134 82 25190 480
rect 25424 377 25452 4966
rect 25504 4684 25556 4690
rect 25504 4626 25556 4632
rect 25516 4282 25544 4626
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 25410 368 25466 377
rect 25410 303 25466 312
rect 24964 54 25190 82
rect 25608 82 25636 5238
rect 25870 82 25926 480
rect 25608 54 25926 82
rect 24858 31 24914 40
rect 25134 0 25190 54
rect 25870 0 25926 54
rect 26698 82 26754 480
rect 26804 82 26832 6598
rect 27342 1184 27398 1193
rect 27342 1119 27398 1128
rect 26698 54 26832 82
rect 27356 82 27384 1119
rect 27526 82 27582 480
rect 27356 54 27582 82
rect 26698 0 26754 54
rect 27526 0 27582 54
<< via2 >>
rect 1122 26832 1178 26888
rect 110 24248 166 24304
rect 18 19080 74 19136
rect 1582 25744 1638 25800
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 2686 24792 2742 24848
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 1582 22616 1638 22672
rect 1490 21664 1546 21720
rect 1582 20576 1638 20632
rect 1582 19624 1638 19680
rect 1582 17448 1638 17504
rect 110 15952 166 16008
rect 1582 14320 1638 14376
rect 18 12144 74 12200
rect 18 6568 74 6624
rect 110 2488 166 2544
rect 202 720 258 776
rect 1582 12300 1638 12336
rect 1582 12280 1584 12300
rect 1584 12280 1636 12300
rect 1636 12280 1638 12300
rect 2226 4936 2282 4992
rect 3422 12144 3478 12200
rect 3422 11192 3478 11248
rect 3514 5208 3570 5264
rect 2686 4936 2742 4992
rect 3790 10240 3846 10296
rect 2594 992 2650 1048
rect 3514 2488 3570 2544
rect 3882 2624 3938 2680
rect 4158 13368 4214 13424
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6550 16496 6606 16552
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6642 11192 6698 11248
rect 4710 7384 4766 7440
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4802 5752 4858 5808
rect 4802 5072 4858 5128
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6826 6296 6882 6352
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4802 4120 4858 4176
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4250 2624 4306 2680
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6090 3168 6146 3224
rect 3606 448 3662 504
rect 6090 2624 6146 2680
rect 7746 4256 7802 4312
rect 7194 3304 7250 3360
rect 6734 2624 6790 2680
rect 5446 992 5502 1048
rect 5354 584 5410 640
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7194 2624 7250 2680
rect 7010 1672 7066 1728
rect 6642 992 6698 1048
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 8758 10104 8814 10160
rect 8390 8472 8446 8528
rect 8390 7656 8446 7712
rect 8666 7792 8722 7848
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 8758 4936 8814 4992
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10046 7384 10102 7440
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9586 4664 9642 4720
rect 9678 4528 9734 4584
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3576 10194 3632
rect 8574 2352 8630 2408
rect 8850 2352 8906 2408
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9954 2352 10010 2408
rect 10690 40 10746 96
rect 11702 11192 11758 11248
rect 11150 3984 11206 4040
rect 11242 2896 11298 2952
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 12254 12144 12310 12200
rect 11334 2488 11390 2544
rect 11610 856 11666 912
rect 12070 5888 12126 5944
rect 12346 7248 12402 7304
rect 12254 5072 12310 5128
rect 11886 3848 11942 3904
rect 12898 12280 12954 12336
rect 12806 6704 12862 6760
rect 12990 2624 13046 2680
rect 12806 1536 12862 1592
rect 12622 1264 12678 1320
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 13542 10104 13598 10160
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 13910 7792 13966 7848
rect 13634 7248 13690 7304
rect 13726 7112 13782 7168
rect 13174 4392 13230 4448
rect 13634 3032 13690 3088
rect 14186 4664 14242 4720
rect 13818 2488 13874 2544
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14738 8744 14794 8800
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14738 8608 14794 8664
rect 14554 7656 14610 7712
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14830 7284 14832 7304
rect 14832 7284 14884 7304
rect 14884 7284 14886 7304
rect 14830 7248 14886 7284
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15658 5344 15714 5400
rect 15566 5208 15622 5264
rect 14462 4528 14518 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14554 3304 14610 3360
rect 14738 2216 14794 2272
rect 13818 1944 13874 2000
rect 12530 312 12586 368
rect 14002 40 14058 96
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15382 3576 15438 3632
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16486 9016 16542 9072
rect 16026 6840 16082 6896
rect 15842 4528 15898 4584
rect 16118 3848 16174 3904
rect 18418 9832 18474 9888
rect 17130 8472 17186 8528
rect 17498 4120 17554 4176
rect 16394 3476 16396 3496
rect 16396 3476 16448 3496
rect 16448 3476 16450 3496
rect 16394 3440 16450 3476
rect 16486 3304 16542 3360
rect 16118 2760 16174 2816
rect 17406 2624 17462 2680
rect 16394 1128 16450 1184
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 18694 5752 18750 5808
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 21822 7928 21878 7984
rect 19430 7112 19486 7168
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19614 5752 19670 5808
rect 19522 5208 19578 5264
rect 19062 5072 19118 5128
rect 19246 3712 19302 3768
rect 19338 2760 19394 2816
rect 19246 2624 19302 2680
rect 18326 584 18382 640
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 21546 7112 21602 7168
rect 21086 6704 21142 6760
rect 20442 3712 20498 3768
rect 20626 3304 20682 3360
rect 21454 3984 21510 4040
rect 20810 3032 20866 3088
rect 20718 2896 20774 2952
rect 20258 856 20314 912
rect 21362 3168 21418 3224
rect 21086 1808 21142 1864
rect 20902 1672 20958 1728
rect 21178 992 21234 1048
rect 23846 6840 23902 6896
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 22282 2760 22338 2816
rect 23018 3440 23074 3496
rect 22466 2352 22522 2408
rect 21546 1536 21602 1592
rect 21362 448 21418 504
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24766 5752 24822 5808
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24122 4392 24178 4448
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23478 3576 23534 3632
rect 23294 720 23350 776
rect 23570 176 23626 232
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24214 2488 24270 2544
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24122 1944 24178 2000
rect 24030 1264 24086 1320
rect 24858 40 24914 96
rect 25410 312 25466 368
rect 27342 1128 27398 1184
<< metal3 >>
rect 0 27344 480 27464
rect 62 26890 122 27344
rect 1117 26890 1183 26893
rect 62 26888 1183 26890
rect 62 26832 1122 26888
rect 1178 26832 1183 26888
rect 62 26830 1183 26832
rect 1117 26827 1183 26830
rect 0 26256 480 26376
rect 62 25802 122 26256
rect 1577 25802 1643 25805
rect 62 25800 1643 25802
rect 62 25744 1582 25800
rect 1638 25744 1643 25800
rect 62 25742 1643 25744
rect 1577 25739 1643 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25304 480 25424
rect 62 24850 122 25304
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 2681 24850 2747 24853
rect 62 24848 2747 24850
rect 62 24792 2686 24848
rect 2742 24792 2747 24848
rect 62 24790 2747 24792
rect 2681 24787 2747 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24304 480 24336
rect 0 24248 110 24304
rect 166 24248 480 24304
rect 0 24216 480 24248
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 62 22674 122 23128
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1577 22674 1643 22677
rect 62 22672 1643 22674
rect 62 22616 1582 22672
rect 1638 22616 1643 22672
rect 62 22614 1643 22616
rect 1577 22611 1643 22614
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1485 21722 1551 21725
rect 62 21720 1551 21722
rect 62 21664 1490 21720
rect 1546 21664 1551 21720
rect 62 21662 1551 21664
rect 1485 21659 1551 21662
rect 10277 21248 10597 21249
rect 0 21088 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 62 20634 122 21088
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1577 20634 1643 20637
rect 62 20632 1643 20634
rect 62 20576 1582 20632
rect 1638 20576 1643 20632
rect 62 20574 1643 20576
rect 1577 20571 1643 20574
rect 10277 20160 10597 20161
rect 0 20000 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 62 19682 122 20000
rect 1577 19682 1643 19685
rect 62 19680 1643 19682
rect 62 19624 1582 19680
rect 1638 19624 1643 19680
rect 62 19622 1643 19624
rect 1577 19619 1643 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19136 480 19168
rect 0 19080 18 19136
rect 74 19080 480 19136
rect 0 19048 480 19080
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 17960 480 18080
rect 10277 17984 10597 17985
rect 62 17506 122 17960
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 1577 17506 1643 17509
rect 62 17504 1643 17506
rect 62 17448 1582 17504
rect 1638 17448 1643 17504
rect 62 17446 1643 17448
rect 1577 17443 1643 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17008 480 17128
rect 62 16554 122 17008
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 6545 16554 6611 16557
rect 62 16552 6611 16554
rect 62 16496 6550 16552
rect 6606 16496 6611 16552
rect 62 16494 6611 16496
rect 6545 16491 6611 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16008 480 16040
rect 0 15952 110 16008
rect 166 15952 480 16008
rect 0 15920 480 15952
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 62 14378 122 14832
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14378 1643 14381
rect 62 14376 1643 14378
rect 62 14320 1582 14376
rect 1638 14320 1643 14376
rect 62 14318 1643 14320
rect 1577 14315 1643 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13880 480 14000
rect 62 13426 122 13880
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4153 13426 4219 13429
rect 62 13424 4219 13426
rect 62 13368 4158 13424
rect 4214 13368 4219 13424
rect 62 13366 4219 13368
rect 4153 13363 4219 13366
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12792 480 12912
rect 62 12338 122 12792
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 1577 12338 1643 12341
rect 12893 12338 12959 12341
rect 62 12336 1643 12338
rect 62 12280 1582 12336
rect 1638 12280 1643 12336
rect 62 12278 1643 12280
rect 1577 12275 1643 12278
rect 1718 12336 12959 12338
rect 1718 12280 12898 12336
rect 12954 12280 12959 12336
rect 1718 12278 12959 12280
rect 13 12202 79 12205
rect 1718 12202 1778 12278
rect 12893 12275 12959 12278
rect 13 12200 1778 12202
rect 13 12144 18 12200
rect 74 12144 1778 12200
rect 13 12142 1778 12144
rect 3417 12202 3483 12205
rect 12249 12202 12315 12205
rect 3417 12200 12315 12202
rect 3417 12144 3422 12200
rect 3478 12144 12254 12200
rect 12310 12144 12315 12200
rect 3417 12142 12315 12144
rect 13 12139 79 12142
rect 3417 12139 3483 12142
rect 12249 12139 12315 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11704 480 11824
rect 62 11250 122 11704
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3417 11250 3483 11253
rect 62 11248 3483 11250
rect 62 11192 3422 11248
rect 3478 11192 3483 11248
rect 62 11190 3483 11192
rect 3417 11187 3483 11190
rect 6637 11250 6703 11253
rect 11697 11250 11763 11253
rect 6637 11248 11763 11250
rect 6637 11192 6642 11248
rect 6698 11192 11702 11248
rect 11758 11192 11763 11248
rect 6637 11190 11763 11192
rect 6637 11187 6703 11190
rect 11697 11187 11763 11190
rect 5610 10912 5930 10913
rect 0 10752 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 62 10298 122 10752
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 3785 10298 3851 10301
rect 62 10296 3851 10298
rect 62 10240 3790 10296
rect 3846 10240 3851 10296
rect 62 10238 3851 10240
rect 3785 10235 3851 10238
rect 8753 10162 8819 10165
rect 13537 10162 13603 10165
rect 8753 10160 13603 10162
rect 8753 10104 8758 10160
rect 8814 10104 13542 10160
rect 13598 10104 13603 10160
rect 8753 10102 13603 10104
rect 8753 10099 8819 10102
rect 13537 10099 13603 10102
rect 238 9964 244 10028
rect 308 10026 314 10028
rect 308 9966 6194 10026
rect 308 9964 314 9966
rect 6134 9890 6194 9966
rect 9622 9890 9628 9892
rect 6134 9830 9628 9890
rect 9622 9828 9628 9830
rect 9692 9828 9698 9892
rect 18270 9828 18276 9892
rect 18340 9890 18346 9892
rect 18413 9890 18479 9893
rect 18340 9888 18479 9890
rect 18340 9832 18418 9888
rect 18474 9832 18479 9888
rect 18340 9830 18479 9832
rect 18340 9828 18346 9830
rect 18413 9827 18479 9830
rect 5610 9824 5930 9825
rect 0 9664 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 62 9630 168 9664
rect 108 9484 168 9630
rect 54 9420 60 9484
rect 124 9422 168 9484
rect 124 9420 130 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12382 9012 12388 9076
rect 12452 9074 12458 9076
rect 16481 9074 16547 9077
rect 12452 9072 16547 9074
rect 12452 9016 16486 9072
rect 16542 9016 16547 9072
rect 12452 9014 16547 9016
rect 12452 9012 12458 9014
rect 16481 9011 16547 9014
rect 0 8712 480 8832
rect 12014 8740 12020 8804
rect 12084 8802 12090 8804
rect 14733 8802 14799 8805
rect 12084 8800 14799 8802
rect 12084 8744 14738 8800
rect 14794 8744 14799 8800
rect 12084 8742 14799 8744
rect 12084 8740 12090 8742
rect 14733 8739 14799 8742
rect 5610 8736 5930 8737
rect 62 8530 122 8712
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 14733 8666 14799 8669
rect 8204 8664 14799 8666
rect 8204 8608 14738 8664
rect 14794 8608 14799 8664
rect 8204 8606 14799 8608
rect 8204 8530 8264 8606
rect 14733 8603 14799 8606
rect 62 8470 8264 8530
rect 8385 8530 8451 8533
rect 8518 8530 8524 8532
rect 8385 8528 8524 8530
rect 8385 8472 8390 8528
rect 8446 8472 8524 8528
rect 8385 8470 8524 8472
rect 8385 8467 8451 8470
rect 8518 8468 8524 8470
rect 8588 8468 8594 8532
rect 15878 8468 15884 8532
rect 15948 8530 15954 8532
rect 17125 8530 17191 8533
rect 15948 8528 17191 8530
rect 15948 8472 17130 8528
rect 17186 8472 17191 8528
rect 15948 8470 17191 8472
rect 15948 8468 15954 8470
rect 17125 8467 17191 8470
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 62 8062 4170 8122
rect 62 7744 122 8062
rect 4110 7986 4170 8062
rect 21817 7986 21883 7989
rect 4110 7984 21883 7986
rect 4110 7928 21822 7984
rect 21878 7928 21883 7984
rect 4110 7926 21883 7928
rect 21817 7923 21883 7926
rect 8661 7850 8727 7853
rect 13905 7850 13971 7853
rect 8661 7848 13971 7850
rect 8661 7792 8666 7848
rect 8722 7792 13910 7848
rect 13966 7792 13971 7848
rect 8661 7790 13971 7792
rect 8661 7787 8727 7790
rect 13905 7787 13971 7790
rect 0 7624 480 7744
rect 8385 7714 8451 7717
rect 14549 7714 14615 7717
rect 8385 7712 14615 7714
rect 8385 7656 8390 7712
rect 8446 7656 14554 7712
rect 14610 7656 14615 7712
rect 8385 7654 14615 7656
rect 8385 7651 8451 7654
rect 14549 7651 14615 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 4705 7442 4771 7445
rect 10041 7442 10107 7445
rect 4705 7440 10107 7442
rect 4705 7384 4710 7440
rect 4766 7384 10046 7440
rect 10102 7384 10107 7440
rect 4705 7382 10107 7384
rect 4705 7379 4771 7382
rect 10041 7379 10107 7382
rect 12341 7306 12407 7309
rect 13629 7306 13695 7309
rect 14825 7306 14891 7309
rect 12341 7304 14891 7306
rect 12341 7248 12346 7304
rect 12402 7248 13634 7304
rect 13690 7248 14830 7304
rect 14886 7248 14891 7304
rect 12341 7246 14891 7248
rect 12341 7243 12407 7246
rect 13629 7243 13695 7246
rect 14825 7243 14891 7246
rect 13721 7170 13787 7173
rect 19425 7170 19491 7173
rect 13721 7168 19491 7170
rect 13721 7112 13726 7168
rect 13782 7112 19430 7168
rect 19486 7112 19491 7168
rect 13721 7110 19491 7112
rect 13721 7107 13787 7110
rect 19425 7107 19491 7110
rect 21398 7108 21404 7172
rect 21468 7170 21474 7172
rect 21541 7170 21607 7173
rect 21468 7168 21607 7170
rect 21468 7112 21546 7168
rect 21602 7112 21607 7168
rect 21468 7110 21607 7112
rect 21468 7108 21474 7110
rect 21541 7107 21607 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 16021 6898 16087 6901
rect 23841 6898 23907 6901
rect 16021 6896 23907 6898
rect 16021 6840 16026 6896
rect 16082 6840 23846 6896
rect 23902 6840 23907 6896
rect 16021 6838 23907 6840
rect 16021 6835 16087 6838
rect 23841 6835 23907 6838
rect 12801 6762 12867 6765
rect 21081 6762 21147 6765
rect 12801 6760 21147 6762
rect 12801 6704 12806 6760
rect 12862 6704 21086 6760
rect 21142 6704 21147 6760
rect 12801 6702 21147 6704
rect 12801 6699 12867 6702
rect 21081 6699 21147 6702
rect 0 6624 480 6656
rect 0 6568 18 6624
rect 74 6568 480 6624
rect 0 6536 480 6568
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 6821 6354 6887 6357
rect 7046 6354 7052 6356
rect 6821 6352 7052 6354
rect 6821 6296 6826 6352
rect 6882 6296 7052 6352
rect 6821 6294 7052 6296
rect 6821 6291 6887 6294
rect 7046 6292 7052 6294
rect 7116 6292 7122 6356
rect 9622 6082 9628 6084
rect 62 6022 9628 6082
rect 62 5704 122 6022
rect 9622 6020 9628 6022
rect 9692 6020 9698 6084
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 12065 5946 12131 5949
rect 12065 5944 19074 5946
rect 12065 5888 12070 5944
rect 12126 5888 19074 5944
rect 12065 5886 19074 5888
rect 12065 5883 12131 5886
rect 4797 5810 4863 5813
rect 18689 5810 18755 5813
rect 4797 5808 18755 5810
rect 4797 5752 4802 5808
rect 4858 5752 18694 5808
rect 18750 5752 18755 5808
rect 4797 5750 18755 5752
rect 19014 5810 19074 5886
rect 19609 5810 19675 5813
rect 19014 5808 19675 5810
rect 19014 5752 19614 5808
rect 19670 5752 19675 5808
rect 19014 5750 19675 5752
rect 4797 5747 4863 5750
rect 18689 5747 18755 5750
rect 19609 5747 19675 5750
rect 23422 5748 23428 5812
rect 23492 5810 23498 5812
rect 24761 5810 24827 5813
rect 23492 5808 24827 5810
rect 23492 5752 24766 5808
rect 24822 5752 24827 5808
rect 23492 5750 24827 5752
rect 23492 5748 23498 5750
rect 24761 5747 24827 5750
rect 0 5584 480 5704
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 15653 5402 15719 5405
rect 15334 5400 15719 5402
rect 15334 5344 15658 5400
rect 15714 5344 15719 5400
rect 15334 5342 15719 5344
rect 3509 5266 3575 5269
rect 15334 5266 15394 5342
rect 15653 5339 15719 5342
rect 3509 5264 15394 5266
rect 3509 5208 3514 5264
rect 3570 5208 15394 5264
rect 3509 5206 15394 5208
rect 15561 5266 15627 5269
rect 19517 5266 19583 5269
rect 15561 5264 19583 5266
rect 15561 5208 15566 5264
rect 15622 5208 19522 5264
rect 19578 5208 19583 5264
rect 15561 5206 19583 5208
rect 3509 5203 3575 5206
rect 15561 5203 15627 5206
rect 19517 5203 19583 5206
rect 4797 5130 4863 5133
rect 62 5128 4863 5130
rect 62 5072 4802 5128
rect 4858 5072 4863 5128
rect 62 5070 4863 5072
rect 62 4616 122 5070
rect 4797 5067 4863 5070
rect 12249 5130 12315 5133
rect 19057 5130 19123 5133
rect 12249 5128 19123 5130
rect 12249 5072 12254 5128
rect 12310 5072 19062 5128
rect 19118 5072 19123 5128
rect 12249 5070 19123 5072
rect 12249 5067 12315 5070
rect 19057 5067 19123 5070
rect 2221 4994 2287 4997
rect 2681 4994 2747 4997
rect 8753 4994 8819 4997
rect 2221 4992 8819 4994
rect 2221 4936 2226 4992
rect 2282 4936 2686 4992
rect 2742 4936 8758 4992
rect 8814 4936 8819 4992
rect 2221 4934 8819 4936
rect 2221 4931 2287 4934
rect 2681 4931 2747 4934
rect 8753 4931 8819 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 9581 4722 9647 4725
rect 14181 4722 14247 4725
rect 9581 4720 14247 4722
rect 9581 4664 9586 4720
rect 9642 4664 14186 4720
rect 14242 4664 14247 4720
rect 9581 4662 14247 4664
rect 9581 4659 9647 4662
rect 14181 4659 14247 4662
rect 0 4496 480 4616
rect 9673 4586 9739 4589
rect 14457 4586 14523 4589
rect 15837 4586 15903 4589
rect 9673 4584 14523 4586
rect 9673 4528 9678 4584
rect 9734 4528 14462 4584
rect 14518 4528 14523 4584
rect 9673 4526 14523 4528
rect 9673 4523 9739 4526
rect 14457 4523 14523 4526
rect 14782 4584 15903 4586
rect 14782 4528 15842 4584
rect 15898 4528 15903 4584
rect 14782 4526 15903 4528
rect 13169 4450 13235 4453
rect 13486 4450 13492 4452
rect 13169 4448 13492 4450
rect 13169 4392 13174 4448
rect 13230 4392 13492 4448
rect 13169 4390 13492 4392
rect 13169 4387 13235 4390
rect 13486 4388 13492 4390
rect 13556 4388 13562 4452
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 7741 4314 7807 4317
rect 14782 4314 14842 4526
rect 15837 4523 15903 4526
rect 23422 4388 23428 4452
rect 23492 4450 23498 4452
rect 24117 4450 24183 4453
rect 23492 4448 24183 4450
rect 23492 4392 24122 4448
rect 24178 4392 24183 4448
rect 23492 4390 24183 4392
rect 23492 4388 23498 4390
rect 24117 4387 24183 4390
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 7741 4312 14842 4314
rect 7741 4256 7746 4312
rect 7802 4256 14842 4312
rect 7741 4254 14842 4256
rect 7741 4251 7807 4254
rect 4797 4178 4863 4181
rect 17493 4178 17559 4181
rect 4797 4176 17559 4178
rect 4797 4120 4802 4176
rect 4858 4120 17498 4176
rect 17554 4120 17559 4176
rect 4797 4118 17559 4120
rect 4797 4115 4863 4118
rect 17493 4115 17559 4118
rect 11145 4042 11211 4045
rect 21449 4042 21515 4045
rect 11145 4040 21515 4042
rect 11145 3984 11150 4040
rect 11206 3984 21454 4040
rect 21510 3984 21515 4040
rect 11145 3982 21515 3984
rect 11145 3979 11211 3982
rect 21449 3979 21515 3982
rect 11881 3906 11947 3909
rect 16113 3906 16179 3909
rect 11881 3904 16179 3906
rect 11881 3848 11886 3904
rect 11942 3848 16118 3904
rect 16174 3848 16179 3904
rect 11881 3846 16179 3848
rect 11881 3843 11947 3846
rect 16113 3843 16179 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 19241 3770 19307 3773
rect 13770 3768 19307 3770
rect 13770 3712 19246 3768
rect 19302 3712 19307 3768
rect 13770 3710 19307 3712
rect 10133 3634 10199 3637
rect 13770 3634 13830 3710
rect 19241 3707 19307 3710
rect 20110 3708 20116 3772
rect 20180 3770 20186 3772
rect 20437 3770 20503 3773
rect 20180 3768 20503 3770
rect 20180 3712 20442 3768
rect 20498 3712 20503 3768
rect 20180 3710 20503 3712
rect 20180 3708 20186 3710
rect 20437 3707 20503 3710
rect 10133 3632 13830 3634
rect 10133 3576 10138 3632
rect 10194 3576 13830 3632
rect 10133 3574 13830 3576
rect 15377 3634 15443 3637
rect 23473 3634 23539 3637
rect 15377 3632 23539 3634
rect 15377 3576 15382 3632
rect 15438 3576 23478 3632
rect 23534 3576 23539 3632
rect 15377 3574 23539 3576
rect 10133 3571 10199 3574
rect 15377 3571 15443 3574
rect 23473 3571 23539 3574
rect 0 3408 480 3528
rect 16389 3498 16455 3501
rect 23013 3498 23079 3501
rect 16389 3496 23079 3498
rect 16389 3440 16394 3496
rect 16450 3440 23018 3496
rect 23074 3440 23079 3496
rect 16389 3438 23079 3440
rect 16389 3435 16455 3438
rect 23013 3435 23079 3438
rect 62 3090 122 3408
rect 7189 3362 7255 3365
rect 14549 3362 14615 3365
rect 7189 3360 14615 3362
rect 7189 3304 7194 3360
rect 7250 3304 14554 3360
rect 14610 3304 14615 3360
rect 7189 3302 14615 3304
rect 7189 3299 7255 3302
rect 14549 3299 14615 3302
rect 16481 3362 16547 3365
rect 20621 3362 20687 3365
rect 16481 3360 20687 3362
rect 16481 3304 16486 3360
rect 16542 3304 20626 3360
rect 20682 3304 20687 3360
rect 16481 3302 20687 3304
rect 16481 3299 16547 3302
rect 20621 3299 20687 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 6085 3226 6151 3229
rect 6085 3224 13830 3226
rect 6085 3168 6090 3224
rect 6146 3168 13830 3224
rect 6085 3166 13830 3168
rect 6085 3163 6151 3166
rect 13629 3090 13695 3093
rect 62 3088 13695 3090
rect 62 3032 13634 3088
rect 13690 3032 13695 3088
rect 62 3030 13695 3032
rect 13770 3090 13830 3166
rect 15878 3164 15884 3228
rect 15948 3226 15954 3228
rect 21357 3226 21423 3229
rect 15948 3224 21423 3226
rect 15948 3168 21362 3224
rect 21418 3168 21423 3224
rect 15948 3166 21423 3168
rect 15948 3164 15954 3166
rect 21357 3163 21423 3166
rect 20805 3090 20871 3093
rect 13770 3088 20871 3090
rect 13770 3032 20810 3088
rect 20866 3032 20871 3088
rect 13770 3030 20871 3032
rect 13629 3027 13695 3030
rect 20805 3027 20871 3030
rect 11237 2954 11303 2957
rect 20713 2954 20779 2957
rect 11237 2952 20779 2954
rect 11237 2896 11242 2952
rect 11298 2896 20718 2952
rect 20774 2896 20779 2952
rect 11237 2894 20779 2896
rect 11237 2891 11303 2894
rect 20713 2891 20779 2894
rect 16113 2818 16179 2821
rect 19333 2818 19399 2821
rect 16113 2816 19399 2818
rect 16113 2760 16118 2816
rect 16174 2760 19338 2816
rect 19394 2760 19399 2816
rect 16113 2758 19399 2760
rect 16113 2755 16179 2758
rect 19333 2755 19399 2758
rect 22134 2756 22140 2820
rect 22204 2818 22210 2820
rect 22277 2818 22343 2821
rect 22204 2816 22343 2818
rect 22204 2760 22282 2816
rect 22338 2760 22343 2816
rect 22204 2758 22343 2760
rect 22204 2756 22210 2758
rect 22277 2755 22343 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3877 2682 3943 2685
rect 4245 2682 4311 2685
rect 6085 2682 6151 2685
rect 3877 2680 6151 2682
rect 3877 2624 3882 2680
rect 3938 2624 4250 2680
rect 4306 2624 6090 2680
rect 6146 2624 6151 2680
rect 3877 2622 6151 2624
rect 3877 2619 3943 2622
rect 4245 2619 4311 2622
rect 6085 2619 6151 2622
rect 6729 2682 6795 2685
rect 7189 2682 7255 2685
rect 6729 2680 7255 2682
rect 6729 2624 6734 2680
rect 6790 2624 7194 2680
rect 7250 2624 7255 2680
rect 6729 2622 7255 2624
rect 6729 2619 6795 2622
rect 7189 2619 7255 2622
rect 12985 2682 13051 2685
rect 16430 2682 16436 2684
rect 12985 2680 16436 2682
rect 12985 2624 12990 2680
rect 13046 2624 16436 2680
rect 12985 2622 16436 2624
rect 12985 2619 13051 2622
rect 16430 2620 16436 2622
rect 16500 2620 16506 2684
rect 17401 2682 17467 2685
rect 19241 2682 19307 2685
rect 17401 2680 19307 2682
rect 17401 2624 17406 2680
rect 17462 2624 19246 2680
rect 19302 2624 19307 2680
rect 17401 2622 19307 2624
rect 17401 2619 17467 2622
rect 19241 2619 19307 2622
rect 0 2544 480 2576
rect 0 2488 110 2544
rect 166 2488 480 2544
rect 0 2456 480 2488
rect 3509 2546 3575 2549
rect 11329 2546 11395 2549
rect 3509 2544 11395 2546
rect 3509 2488 3514 2544
rect 3570 2488 11334 2544
rect 11390 2488 11395 2544
rect 3509 2486 11395 2488
rect 3509 2483 3575 2486
rect 11329 2483 11395 2486
rect 13813 2546 13879 2549
rect 24209 2546 24275 2549
rect 13813 2544 24275 2546
rect 13813 2488 13818 2544
rect 13874 2488 24214 2544
rect 24270 2488 24275 2544
rect 13813 2486 24275 2488
rect 13813 2483 13879 2486
rect 24209 2483 24275 2486
rect 8569 2410 8635 2413
rect 8702 2410 8708 2412
rect 8569 2408 8708 2410
rect 8569 2352 8574 2408
rect 8630 2352 8708 2408
rect 8569 2350 8708 2352
rect 8569 2347 8635 2350
rect 8702 2348 8708 2350
rect 8772 2348 8778 2412
rect 8845 2410 8911 2413
rect 9949 2410 10015 2413
rect 22461 2410 22527 2413
rect 8845 2408 9690 2410
rect 8845 2352 8850 2408
rect 8906 2352 9690 2408
rect 8845 2350 9690 2352
rect 8845 2347 8911 2350
rect 9630 2274 9690 2350
rect 9949 2408 22527 2410
rect 9949 2352 9954 2408
rect 10010 2352 22466 2408
rect 22522 2352 22527 2408
rect 9949 2350 22527 2352
rect 9949 2347 10015 2350
rect 22461 2347 22527 2350
rect 14733 2274 14799 2277
rect 9630 2272 14799 2274
rect 9630 2216 14738 2272
rect 14794 2216 14799 2272
rect 9630 2214 14799 2216
rect 14733 2211 14799 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 13813 2002 13879 2005
rect 24117 2002 24183 2005
rect 13813 2000 24183 2002
rect 13813 1944 13818 2000
rect 13874 1944 24122 2000
rect 24178 1944 24183 2000
rect 13813 1942 24183 1944
rect 13813 1939 13879 1942
rect 24117 1939 24183 1942
rect 21081 1866 21147 1869
rect 13770 1864 21147 1866
rect 13770 1808 21086 1864
rect 21142 1808 21147 1864
rect 13770 1806 21147 1808
rect 54 1668 60 1732
rect 124 1730 130 1732
rect 7005 1730 7071 1733
rect 13770 1730 13830 1806
rect 21081 1803 21147 1806
rect 124 1670 674 1730
rect 124 1668 130 1670
rect 614 1594 674 1670
rect 7005 1728 13830 1730
rect 7005 1672 7010 1728
rect 7066 1672 13830 1728
rect 7005 1670 13830 1672
rect 7005 1667 7071 1670
rect 17534 1668 17540 1732
rect 17604 1730 17610 1732
rect 20897 1730 20963 1733
rect 17604 1728 20963 1730
rect 17604 1672 20902 1728
rect 20958 1672 20963 1728
rect 17604 1670 20963 1672
rect 17604 1668 17610 1670
rect 20897 1667 20963 1670
rect 12014 1594 12020 1596
rect 614 1534 12020 1594
rect 12014 1532 12020 1534
rect 12084 1532 12090 1596
rect 12801 1594 12867 1597
rect 21541 1594 21607 1597
rect 12801 1592 21607 1594
rect 12801 1536 12806 1592
rect 12862 1536 21546 1592
rect 21602 1536 21607 1592
rect 12801 1534 21607 1536
rect 12801 1531 12867 1534
rect 21541 1531 21607 1534
rect 0 1460 480 1488
rect 0 1396 60 1460
rect 124 1396 480 1460
rect 0 1368 480 1396
rect 12382 1322 12388 1324
rect 9630 1262 12388 1322
rect 9630 1186 9690 1262
rect 12382 1260 12388 1262
rect 12452 1260 12458 1324
rect 12617 1322 12683 1325
rect 24025 1322 24091 1325
rect 12617 1320 24091 1322
rect 12617 1264 12622 1320
rect 12678 1264 24030 1320
rect 24086 1264 24091 1320
rect 12617 1262 24091 1264
rect 12617 1259 12683 1262
rect 24025 1259 24091 1262
rect 62 1126 9690 1186
rect 16389 1186 16455 1189
rect 27337 1186 27403 1189
rect 16389 1184 27403 1186
rect 16389 1128 16394 1184
rect 16450 1128 27342 1184
rect 27398 1128 27403 1184
rect 16389 1126 27403 1128
rect 62 536 122 1126
rect 16389 1123 16455 1126
rect 27337 1123 27403 1126
rect 2589 1050 2655 1053
rect 4102 1050 4108 1052
rect 2589 1048 4108 1050
rect 2589 992 2594 1048
rect 2650 992 4108 1048
rect 2589 990 4108 992
rect 2589 987 2655 990
rect 4102 988 4108 990
rect 4172 988 4178 1052
rect 5441 1050 5507 1053
rect 5574 1050 5580 1052
rect 5441 1048 5580 1050
rect 5441 992 5446 1048
rect 5502 992 5580 1048
rect 5441 990 5580 992
rect 5441 987 5507 990
rect 5574 988 5580 990
rect 5644 988 5650 1052
rect 6637 1050 6703 1053
rect 21173 1050 21239 1053
rect 6637 1048 21239 1050
rect 6637 992 6642 1048
rect 6698 992 21178 1048
rect 21234 992 21239 1048
rect 6637 990 21239 992
rect 6637 987 6703 990
rect 21173 987 21239 990
rect 11605 914 11671 917
rect 20253 914 20319 917
rect 11605 912 20319 914
rect 11605 856 11610 912
rect 11666 856 20258 912
rect 20314 856 20319 912
rect 11605 854 20319 856
rect 11605 851 11671 854
rect 20253 851 20319 854
rect 197 778 263 781
rect 23289 778 23355 781
rect 197 776 23355 778
rect 197 720 202 776
rect 258 720 23294 776
rect 23350 720 23355 776
rect 197 718 23355 720
rect 197 715 263 718
rect 23289 715 23355 718
rect 5349 642 5415 645
rect 18321 642 18387 645
rect 5349 640 18387 642
rect 5349 584 5354 640
rect 5410 584 18326 640
rect 18382 584 18387 640
rect 5349 582 18387 584
rect 5349 579 5415 582
rect 18321 579 18387 582
rect 0 416 480 536
rect 3601 506 3667 509
rect 21357 506 21423 509
rect 3601 504 21423 506
rect 3601 448 3606 504
rect 3662 448 21362 504
rect 21418 448 21423 504
rect 3601 446 21423 448
rect 3601 443 3667 446
rect 21357 443 21423 446
rect 12525 370 12591 373
rect 25405 370 25471 373
rect 12525 368 25471 370
rect 12525 312 12530 368
rect 12586 312 25410 368
rect 25466 312 25471 368
rect 12525 310 25471 312
rect 12525 307 12591 310
rect 25405 307 25471 310
rect 23565 234 23631 237
rect 13770 232 23631 234
rect 13770 176 23570 232
rect 23626 176 23631 232
rect 13770 174 23631 176
rect 10685 98 10751 101
rect 13770 98 13830 174
rect 23565 171 23631 174
rect 10685 96 13830 98
rect 10685 40 10690 96
rect 10746 40 13830 96
rect 10685 38 13830 40
rect 13997 98 14063 101
rect 24853 98 24919 101
rect 13997 96 24919 98
rect 13997 40 14002 96
rect 14058 40 24858 96
rect 24914 40 24919 96
rect 13997 38 24919 40
rect 10685 35 10751 38
rect 13997 35 14063 38
rect 24853 35 24919 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 244 9964 308 10028
rect 9628 9828 9692 9892
rect 18276 9828 18340 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 60 9420 124 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 12388 9012 12452 9076
rect 12020 8740 12084 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 8524 8468 8588 8532
rect 15884 8468 15948 8532
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 21404 7108 21468 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 7052 6292 7116 6356
rect 9628 6020 9692 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 23428 5748 23492 5812
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 13492 4388 13556 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 23428 4388 23492 4452
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 20116 3708 20180 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 15884 3164 15948 3228
rect 22140 2756 22204 2820
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 16436 2620 16500 2684
rect 8708 2348 8772 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 60 1668 124 1732
rect 17540 1668 17604 1732
rect 12020 1532 12084 1596
rect 60 1396 124 1460
rect 12388 1260 12452 1324
rect 4108 988 4172 1052
rect 5580 988 5644 1052
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 243 10028 309 10029
rect 243 9964 244 10028
rect 308 9964 309 10028
rect 243 9963 309 9964
rect 246 9690 306 9963
rect 62 9630 306 9690
rect 5610 9824 5931 10848
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 62 9485 122 9630
rect 59 9484 125 9485
rect 59 9420 60 9484
rect 124 9420 125 9484
rect 59 9419 125 9420
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 10277 8192 10597 9216
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 12387 9076 12453 9077
rect 12387 9012 12388 9076
rect 12452 9012 12453 9076
rect 12387 9011 12453 9012
rect 12019 8804 12085 8805
rect 12019 8740 12020 8804
rect 12084 8740 12085 8804
rect 12019 8739 12085 8740
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 7051 6356 7117 6357
rect 7051 6292 7052 6356
rect 7116 6292 7117 6356
rect 7051 6291 7117 6292
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 7054 5218 7114 6291
rect 9630 6085 9690 7022
rect 9627 6084 9693 6085
rect 9627 6020 9628 6084
rect 9692 6020 9693 6084
rect 9627 6019 9693 6020
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2128 10597 2688
rect 59 1732 125 1733
rect 59 1668 60 1732
rect 124 1668 125 1732
rect 59 1667 125 1668
rect 62 1461 122 1667
rect 12022 1597 12082 8739
rect 12019 1596 12085 1597
rect 59 1460 125 1461
rect 59 1396 60 1460
rect 124 1396 125 1460
rect 59 1395 125 1396
rect 4110 1053 4170 1582
rect 12019 1532 12020 1596
rect 12084 1532 12085 1596
rect 12019 1531 12085 1532
rect 12390 1325 12450 9011
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 15883 3228 15949 3229
rect 15883 3164 15884 3228
rect 15948 3164 15949 3228
rect 15883 3163 15949 3164
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 12387 1324 12453 1325
rect 12387 1260 12388 1324
rect 12452 1260 12453 1324
rect 12387 1259 12453 1260
rect 15886 1138 15946 3163
rect 16438 2685 16498 3622
rect 19610 2752 19930 3776
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 22139 2820 22205 2821
rect 22139 2756 22140 2820
rect 22204 2756 22205 2820
rect 22139 2755 22205 2756
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 16435 2684 16501 2685
rect 16435 2620 16436 2684
rect 16500 2620 16501 2684
rect 16435 2619 16501 2620
rect 19610 2128 19930 2688
rect 22142 2498 22202 2755
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 4107 1052 4173 1053
rect 4107 988 4108 1052
rect 4172 988 4173 1052
rect 4107 987 4173 988
<< via4 >>
rect 9542 9892 9778 9978
rect 9542 9828 9628 9892
rect 9628 9828 9692 9892
rect 9692 9828 9778 9892
rect 9542 9742 9778 9828
rect 8438 8532 8674 8618
rect 8438 8468 8524 8532
rect 8524 8468 8588 8532
rect 8588 8468 8674 8532
rect 8438 8382 8674 8468
rect 9542 7022 9778 7258
rect 6966 4982 7202 5218
rect 8622 2412 8858 2498
rect 8622 2348 8708 2412
rect 8708 2348 8772 2412
rect 8772 2348 8858 2412
rect 8622 2262 8858 2348
rect 4022 1582 4258 1818
rect 18190 9892 18426 9978
rect 18190 9828 18276 9892
rect 18276 9828 18340 9892
rect 18340 9828 18426 9892
rect 18190 9742 18426 9828
rect 15798 8532 16034 8618
rect 15798 8468 15884 8532
rect 15884 8468 15948 8532
rect 15948 8468 16034 8532
rect 15798 8382 16034 8468
rect 13406 4452 13642 4538
rect 13406 4388 13492 4452
rect 13492 4388 13556 4452
rect 13556 4388 13642 4452
rect 13406 4302 13642 4388
rect 21318 7172 21554 7258
rect 21318 7108 21404 7172
rect 21404 7108 21468 7172
rect 21468 7108 21554 7172
rect 21318 7022 21554 7108
rect 23342 5812 23578 5898
rect 23342 5748 23428 5812
rect 23428 5748 23492 5812
rect 23492 5748 23578 5812
rect 23342 5662 23578 5748
rect 16350 3622 16586 3858
rect 23342 4452 23578 4538
rect 23342 4388 23428 4452
rect 23428 4388 23492 4452
rect 23492 4388 23578 4452
rect 23342 4302 23578 4388
rect 20030 3772 20266 3858
rect 20030 3708 20116 3772
rect 20116 3708 20180 3772
rect 20180 3708 20266 3772
rect 20030 3622 20266 3708
rect 22054 2262 22290 2498
rect 17454 1732 17690 1818
rect 17454 1668 17540 1732
rect 17540 1668 17604 1732
rect 17604 1668 17690 1732
rect 17454 1582 17690 1668
rect 5494 1052 5730 1138
rect 5494 988 5580 1052
rect 5580 988 5644 1052
rect 5644 988 5730 1052
rect 5494 902 5730 988
rect 15798 902 16034 1138
<< metal5 >>
rect 9500 9978 18468 10020
rect 9500 9742 9542 9978
rect 9778 9742 18190 9978
rect 18426 9742 18468 9978
rect 9500 9700 18468 9742
rect 8396 8618 16076 8660
rect 8396 8382 8438 8618
rect 8674 8382 15798 8618
rect 16034 8382 16076 8618
rect 8396 8340 16076 8382
rect 9500 7258 21596 7300
rect 9500 7022 9542 7258
rect 9778 7022 21318 7258
rect 21554 7022 21596 7258
rect 9500 6980 21596 7022
rect 13640 5898 23620 5940
rect 13640 5662 23342 5898
rect 23578 5662 23620 5898
rect 13640 5620 23620 5662
rect 13640 5260 13960 5620
rect 6924 5218 13960 5260
rect 6924 4982 6966 5218
rect 7202 4982 13960 5218
rect 6924 4940 13960 4982
rect 18378 4940 20124 5260
rect 18378 4580 18698 4940
rect 13364 4538 18698 4580
rect 13364 4302 13406 4538
rect 13642 4302 18698 4538
rect 13364 4260 18698 4302
rect 19804 4580 20124 4940
rect 19804 4538 23620 4580
rect 19804 4302 23342 4538
rect 23578 4302 23620 4538
rect 19068 3900 19480 4300
rect 19804 4260 23620 4302
rect 16308 3858 20308 3900
rect 16308 3622 16350 3858
rect 16586 3622 20030 3858
rect 20266 3622 20308 3858
rect 16308 3580 20308 3622
rect 8580 2498 22332 2540
rect 8580 2262 8622 2498
rect 8858 2262 22054 2498
rect 22290 2262 22332 2498
rect 8580 2220 22332 2262
rect 3980 1818 17732 1860
rect 3980 1582 4022 1818
rect 4258 1582 17454 1818
rect 17690 1582 17732 1818
rect 3980 1540 17732 1582
rect 5452 1138 16076 1180
rect 5452 902 5494 1138
rect 5730 902 15798 1138
rect 16034 902 16076 1138
rect 5452 860 16076 902
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _214_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_154
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_156 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _235_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_161
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_172
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_199
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_195
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_212
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_216
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _189_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_227 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_234
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_253
timestamp 1586364061
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_257
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_265
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_264 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_110
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_139
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 1472 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_13
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _112_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_79
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_83
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_243
timestamp 1586364061
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_248
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_252
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_267
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 2116 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_20
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_24
timestamp 1586364061
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_43
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_52
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_1  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_169
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_224
timestamp 1586364061
transform 1 0 21712 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_237
timestamp 1586364061
transform 1 0 22908 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_8  FILLER_4_248
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_22
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 130 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_175 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 774 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_256
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_267
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_13
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_18
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_14
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_24
timestamp 1586364061
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_28
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_37
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_39
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_35
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_43
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 866 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_73
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 314 592
use scs8hd_or4_4  _104_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_157
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_161
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 406 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_210
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_214
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_235
timestamp 1586364061
transform 1 0 22724 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_246
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_248
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_258
timestamp 1586364061
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_270
timestamp 1586364061
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_35
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_63
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_67
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_71
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_188
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_218
timestamp 1586364061
transform 1 0 21160 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_229
timestamp 1586364061
transform 1 0 22172 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_14
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_18
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_249
timestamp 1586364061
transform 1 0 24012 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_209
timestamp 1586364061
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_87
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_202
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_8
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_21
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_25
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_43
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_47
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_115
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_135
timestamp 1586364061
transform 1 0 13524 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_196
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_200
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_14
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 590 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_71
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_115
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_decap_6  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_23
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 406 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_17
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_25
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_29
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_6  FILLER_16_51
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_77
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_99
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_116
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_157
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_181
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_193
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_nor3_4  _168_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_115
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_178
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_76
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_130
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_12
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_26
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_41
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 8464 0 1 12512
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_113
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_124
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_154
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_178
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_14
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_26
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_120
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_13
timestamp 1586364061
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_17
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_25
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_53
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_36
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_94
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 590 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_66
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 130 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_70
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_70
timestamp 1586364061
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_87
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_117
timestamp 1586364061
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_25
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_52
timestamp 1586364061
transform 1 0 5888 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_63
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_75
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_16
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_38
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 130 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_42
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_47
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_59
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_71
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_29
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_41
timestamp 1586364061
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_14
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_42
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_54
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_19
timestamp 1586364061
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 15566 0 15622 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 16302 0 16358 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 17130 0 17186 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 17958 0 18014 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 18694 0 18750 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 19522 0 19578 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 13910 0 13966 480 6 bottom_left_grid_pin_13_
port 6 nsew default input
rlabel metal2 s 11518 0 11574 480 6 bottom_right_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 12346 0 12402 480 6 bottom_right_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 13082 0 13138 480 6 bottom_right_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 7562 0 7618 480 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 8298 0 8354 480 6 bottom_right_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 9126 0 9182 480 6 bottom_right_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 9954 0 10010 480 6 bottom_right_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 10690 0 10746 480 6 bottom_right_grid_pin_9_
port 14 nsew default input
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal2 s 386 0 442 480 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 1122 0 1178 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal2 s 2778 0 2834 480 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 5170 0 5226 480 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 25134 0 25190 480 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 25870 0 25926 480 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 26698 0 26754 480 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 data_in
port 51 nsew default input
rlabel metal2 s 14738 0 14794 480 6 enable
port 52 nsew default input
rlabel metal3 s 0 17960 480 18080 6 left_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal3 s 0 14832 480 14952 6 left_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 0 15920 480 16040 6 left_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 0 17008 480 17128 6 left_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 0 9664 480 9784 6 left_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 0 10752 480 10872 6 left_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 11704 480 11824 6 left_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 0 12792 480 12912 6 left_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 0 13880 480 14000 6 left_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
