VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__1_
  CLASS BLOCK ;
  FOREIGN sb_0__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.070 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.560 0.000 108.840 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.240 0.000 112.520 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.380 0.000 116.660 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.060 0.000 120.340 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.200 0.000 124.480 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.880 0.000 128.160 2.400 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.020 0.000 132.300 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.320 0.000 19.600 2.400 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.000 0.000 23.280 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.140 0.000 27.420 2.400 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.000 0.000 0.280 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.680 0.000 3.960 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.360 0.000 7.640 2.400 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.500 0.000 11.780 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.180 0.000 15.460 2.400 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.740 0.000 101.020 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 15.680 138.070 16.280 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 22.480 138.070 23.080 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 29.280 138.070 29.880 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 36.080 138.070 36.680 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 42.200 138.070 42.800 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 49.000 138.070 49.600 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 55.800 138.070 56.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 62.600 138.070 63.200 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 69.400 138.070 70.000 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 75.520 138.070 76.120 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 82.320 138.070 82.920 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 89.120 138.070 89.720 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 95.920 138.070 96.520 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 102.720 138.070 103.320 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 108.840 138.070 109.440 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 115.640 138.070 116.240 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 122.440 138.070 123.040 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.670 129.240 138.070 129.840 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.820 0.000 31.100 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.960 0.000 35.240 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.640 0.000 38.920 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.320 0.000 42.600 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.460 0.000 46.740 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.140 0.000 50.420 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.280 0.000 54.560 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.960 0.000 58.240 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.100 0.000 62.380 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.780 0.000 66.060 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.920 0.000 70.200 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.600 0.000 73.880 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.280 0.000 77.560 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.420 0.000 81.700 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.100 0.000 85.380 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.240 0.000 89.520 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.920 0.000 93.200 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.060 0.000 97.340 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.240 137.600 43.520 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.760 137.600 49.040 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.820 137.600 54.100 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.340 137.600 59.620 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.860 137.600 65.140 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.380 137.600 70.660 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.440 137.600 75.720 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.960 137.600 81.240 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.480 137.600 86.760 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.540 137.600 91.820 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.060 137.600 97.340 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.580 137.600 102.860 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.640 137.600 107.920 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.160 137.600 113.440 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.680 137.600 118.960 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.740 137.600 124.020 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.260 137.600 129.540 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.780 137.600 135.060 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.700 0.000 135.980 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.880 0.000 105.160 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 136.040 138.070 136.640 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 8.880 138.070 9.480 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.140 137.600 27.420 140.000 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.660 137.600 32.940 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.720 137.600 38.000 140.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.460 137.600 0.740 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.520 137.600 5.800 140.000 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.040 137.600 11.320 140.000 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.560 137.600 16.840 140.000 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.620 137.600 21.900 140.000 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.670 2.760 138.070 3.360 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 26.125 10.640 27.725 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 49.455 10.640 51.055 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 3.590 10.795 132.390 127.925 ;
      LAYER met1 ;
        RECT 0.440 0.040 136.000 137.660 ;
      LAYER met2 ;
        RECT 1.020 137.320 5.240 137.770 ;
        RECT 6.080 137.320 10.760 137.770 ;
        RECT 11.600 137.320 16.280 137.770 ;
        RECT 17.120 137.320 21.340 137.770 ;
        RECT 22.180 137.320 26.860 137.770 ;
        RECT 27.700 137.320 32.380 137.770 ;
        RECT 33.220 137.320 37.440 137.770 ;
        RECT 38.280 137.320 42.960 137.770 ;
        RECT 43.800 137.320 48.480 137.770 ;
        RECT 49.320 137.320 53.540 137.770 ;
        RECT 54.380 137.320 59.060 137.770 ;
        RECT 59.900 137.320 64.580 137.770 ;
        RECT 65.420 137.320 70.100 137.770 ;
        RECT 70.940 137.320 75.160 137.770 ;
        RECT 76.000 137.320 80.680 137.770 ;
        RECT 81.520 137.320 86.200 137.770 ;
        RECT 87.040 137.320 91.260 137.770 ;
        RECT 92.100 137.320 96.780 137.770 ;
        RECT 97.620 137.320 102.300 137.770 ;
        RECT 103.140 137.320 107.360 137.770 ;
        RECT 108.200 137.320 112.880 137.770 ;
        RECT 113.720 137.320 118.400 137.770 ;
        RECT 119.240 137.320 123.460 137.770 ;
        RECT 124.300 137.320 128.980 137.770 ;
        RECT 129.820 137.320 134.500 137.770 ;
        RECT 135.340 137.320 136.440 137.770 ;
        RECT 0.280 2.680 136.440 137.320 ;
        RECT 0.560 0.010 3.400 2.680 ;
        RECT 4.240 0.010 7.080 2.680 ;
        RECT 7.920 0.010 11.220 2.680 ;
        RECT 12.060 0.010 14.900 2.680 ;
        RECT 15.740 0.010 19.040 2.680 ;
        RECT 19.880 0.010 22.720 2.680 ;
        RECT 23.560 0.010 26.860 2.680 ;
        RECT 27.700 0.010 30.540 2.680 ;
        RECT 31.380 0.010 34.680 2.680 ;
        RECT 35.520 0.010 38.360 2.680 ;
        RECT 39.200 0.010 42.040 2.680 ;
        RECT 42.880 0.010 46.180 2.680 ;
        RECT 47.020 0.010 49.860 2.680 ;
        RECT 50.700 0.010 54.000 2.680 ;
        RECT 54.840 0.010 57.680 2.680 ;
        RECT 58.520 0.010 61.820 2.680 ;
        RECT 62.660 0.010 65.500 2.680 ;
        RECT 66.340 0.010 69.640 2.680 ;
        RECT 70.480 0.010 73.320 2.680 ;
        RECT 74.160 0.010 77.000 2.680 ;
        RECT 77.840 0.010 81.140 2.680 ;
        RECT 81.980 0.010 84.820 2.680 ;
        RECT 85.660 0.010 88.960 2.680 ;
        RECT 89.800 0.010 92.640 2.680 ;
        RECT 93.480 0.010 96.780 2.680 ;
        RECT 97.620 0.010 100.460 2.680 ;
        RECT 101.300 0.010 104.600 2.680 ;
        RECT 105.440 0.010 108.280 2.680 ;
        RECT 109.120 0.010 111.960 2.680 ;
        RECT 112.800 0.010 116.100 2.680 ;
        RECT 116.940 0.010 119.780 2.680 ;
        RECT 120.620 0.010 123.920 2.680 ;
        RECT 124.760 0.010 127.600 2.680 ;
        RECT 128.440 0.010 131.740 2.680 ;
        RECT 132.580 0.010 135.420 2.680 ;
        RECT 136.260 0.010 136.440 2.680 ;
      LAYER met3 ;
        RECT 10.095 135.640 135.270 136.040 ;
        RECT 10.095 130.240 136.720 135.640 ;
        RECT 10.095 128.840 135.270 130.240 ;
        RECT 10.095 123.440 136.720 128.840 ;
        RECT 10.095 122.040 135.270 123.440 ;
        RECT 10.095 116.640 136.720 122.040 ;
        RECT 10.095 115.240 135.270 116.640 ;
        RECT 10.095 109.840 136.720 115.240 ;
        RECT 10.095 108.440 135.270 109.840 ;
        RECT 10.095 103.720 136.720 108.440 ;
        RECT 10.095 102.320 135.270 103.720 ;
        RECT 10.095 96.920 136.720 102.320 ;
        RECT 10.095 95.520 135.270 96.920 ;
        RECT 10.095 90.120 136.720 95.520 ;
        RECT 10.095 88.720 135.270 90.120 ;
        RECT 10.095 83.320 136.720 88.720 ;
        RECT 10.095 81.920 135.270 83.320 ;
        RECT 10.095 76.520 136.720 81.920 ;
        RECT 10.095 75.120 135.270 76.520 ;
        RECT 10.095 70.400 136.720 75.120 ;
        RECT 10.095 69.000 135.270 70.400 ;
        RECT 10.095 63.600 136.720 69.000 ;
        RECT 10.095 62.200 135.270 63.600 ;
        RECT 10.095 56.800 136.720 62.200 ;
        RECT 10.095 55.400 135.270 56.800 ;
        RECT 10.095 50.000 136.720 55.400 ;
        RECT 10.095 48.600 135.270 50.000 ;
        RECT 10.095 43.200 136.720 48.600 ;
        RECT 10.095 41.800 135.270 43.200 ;
        RECT 10.095 37.080 136.720 41.800 ;
        RECT 10.095 35.680 135.270 37.080 ;
        RECT 10.095 30.280 136.720 35.680 ;
        RECT 10.095 28.880 135.270 30.280 ;
        RECT 10.095 23.480 136.720 28.880 ;
        RECT 10.095 22.080 135.270 23.480 ;
        RECT 10.095 16.680 136.720 22.080 ;
        RECT 10.095 15.280 135.270 16.680 ;
        RECT 10.095 9.880 136.720 15.280 ;
        RECT 10.095 8.480 135.270 9.880 ;
        RECT 10.095 3.760 136.720 8.480 ;
        RECT 10.095 2.895 135.270 3.760 ;
      LAYER met4 ;
        RECT 21.860 10.640 25.725 128.080 ;
        RECT 28.125 10.640 49.055 128.080 ;
        RECT 51.455 10.640 136.695 128.080 ;
      LAYER met5 ;
        RECT 21.650 11.100 85.810 33.100 ;
  END
END sb_0__1_
END LIBRARY

