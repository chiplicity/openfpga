magic
tech sky130A
magscale 1 2
timestamp 1605114789
<< locali >>
rect 38905 236879 38939 236981
rect 31947 236777 32005 236811
rect 26485 236607 26519 236777
rect 48473 236539 48507 236981
rect 96865 236811 96899 236913
rect 70587 236709 70645 236743
rect 77545 236675 77579 236777
rect 89965 236675 89999 236777
rect 80247 236641 80305 236675
rect 106433 236675 106467 236913
rect 48565 236471 48599 236573
rect 58133 236471 58167 236641
rect 123177 151539 123211 151913
rect 59421 134539 59455 144025
rect 59329 115159 59363 132941
rect 90609 37843 90643 44541
rect 137989 40563 138023 40665
rect 90701 22407 90735 28085
rect 74785 18055 74819 18361
rect 76073 18259 76107 18429
rect 106525 18327 106559 18429
rect 87205 17987 87239 18089
rect 96773 17987 96807 18293
rect 109745 18191 109779 18429
rect 145165 18259 145199 18361
rect 128547 18225 128605 18259
rect 116185 18055 116219 18157
rect 125753 18055 125787 18225
<< viali >>
rect 38905 236981 38939 237015
rect 38905 236845 38939 236879
rect 48473 236981 48507 237015
rect 26485 236777 26519 236811
rect 31913 236777 31947 236811
rect 32005 236777 32039 236811
rect 26485 236573 26519 236607
rect 96865 236913 96899 236947
rect 77545 236777 77579 236811
rect 70553 236709 70587 236743
rect 70645 236709 70679 236743
rect 89965 236777 89999 236811
rect 96865 236777 96899 236811
rect 106433 236913 106467 236947
rect 58133 236641 58167 236675
rect 77545 236641 77579 236675
rect 80213 236641 80247 236675
rect 80305 236641 80339 236675
rect 89965 236641 89999 236675
rect 106433 236641 106467 236675
rect 48473 236505 48507 236539
rect 48565 236573 48599 236607
rect 48565 236437 48599 236471
rect 58133 236437 58167 236471
rect 123177 151913 123211 151947
rect 123177 151505 123211 151539
rect 59421 144025 59455 144059
rect 59421 134505 59455 134539
rect 59329 132941 59363 132975
rect 59329 115125 59363 115159
rect 90609 44541 90643 44575
rect 137989 40665 138023 40699
rect 137989 40529 138023 40563
rect 90609 37809 90643 37843
rect 90701 28085 90735 28119
rect 90701 22373 90735 22407
rect 76073 18429 76107 18463
rect 74785 18361 74819 18395
rect 106525 18429 106559 18463
rect 76073 18225 76107 18259
rect 96773 18293 96807 18327
rect 106525 18293 106559 18327
rect 109745 18429 109779 18463
rect 74785 18021 74819 18055
rect 87205 18089 87239 18123
rect 87205 17953 87239 17987
rect 145165 18361 145199 18395
rect 125753 18225 125787 18259
rect 128513 18225 128547 18259
rect 128605 18225 128639 18259
rect 145165 18225 145199 18259
rect 109745 18157 109779 18191
rect 116185 18157 116219 18191
rect 116185 18021 116219 18055
rect 125753 18021 125787 18055
rect 96773 17953 96807 17987
<< metal1 >>
rect 99610 244248 99616 244300
rect 99668 244288 99674 244300
rect 99794 244288 99800 244300
rect 99668 244260 99800 244288
rect 99668 244248 99674 244260
rect 99794 244248 99800 244260
rect 99852 244248 99858 244300
rect 89858 241324 89864 241376
rect 89916 241364 89922 241376
rect 171830 241364 171836 241376
rect 89916 241336 171836 241364
rect 89916 241324 89922 241336
rect 171830 241324 171836 241336
rect 171888 241324 171894 241376
rect 174038 241324 174044 241376
rect 174096 241364 174102 241376
rect 207802 241364 207808 241376
rect 174096 241336 207808 241364
rect 174096 241324 174102 241336
rect 207802 241324 207808 241336
rect 207860 241324 207866 241376
rect 27850 241120 27856 241172
rect 27908 241160 27914 241172
rect 29138 241160 29144 241172
rect 27908 241132 29144 241160
rect 27908 241120 27914 241132
rect 29138 241120 29144 241132
rect 29196 241120 29202 241172
rect 135858 240712 135864 240764
rect 135916 240752 135922 240764
rect 136778 240752 136784 240764
rect 135916 240724 136784 240752
rect 135916 240712 135922 240724
rect 136778 240712 136784 240724
rect 136836 240712 136842 240764
rect 38893 237015 38951 237021
rect 38893 236981 38905 237015
rect 38939 237012 38951 237015
rect 48461 237015 48519 237021
rect 48461 237012 48473 237015
rect 38939 236984 48473 237012
rect 38939 236981 38951 236984
rect 38893 236975 38951 236981
rect 48461 236981 48473 236984
rect 48507 236981 48519 237015
rect 48461 236975 48519 236981
rect 96853 236947 96911 236953
rect 96853 236913 96865 236947
rect 96899 236944 96911 236947
rect 106421 236947 106479 236953
rect 106421 236944 106433 236947
rect 96899 236916 106433 236944
rect 96899 236913 96911 236916
rect 96853 236907 96911 236913
rect 106421 236913 106433 236916
rect 106467 236913 106479 236947
rect 106421 236907 106479 236913
rect 38893 236879 38951 236885
rect 38893 236876 38905 236879
rect 32192 236848 38905 236876
rect 26473 236811 26531 236817
rect 26473 236777 26485 236811
rect 26519 236808 26531 236811
rect 31901 236811 31959 236817
rect 31901 236808 31913 236811
rect 26519 236780 31913 236808
rect 26519 236777 26531 236780
rect 26473 236771 26531 236777
rect 31901 236777 31913 236780
rect 31947 236777 31959 236811
rect 31901 236771 31959 236777
rect 31993 236811 32051 236817
rect 31993 236777 32005 236811
rect 32039 236808 32051 236811
rect 32192 236808 32220 236848
rect 38893 236845 38905 236848
rect 38939 236845 38951 236879
rect 38893 236839 38951 236845
rect 77533 236811 77591 236817
rect 77533 236808 77545 236811
rect 32039 236780 32220 236808
rect 72672 236780 77545 236808
rect 32039 236777 32051 236780
rect 31993 236771 32051 236777
rect 62534 236740 62540 236752
rect 60896 236712 62540 236740
rect 12762 236632 12768 236684
rect 12820 236672 12826 236684
rect 30426 236672 30432 236684
rect 12820 236644 30432 236672
rect 12820 236632 12826 236644
rect 30426 236632 30432 236644
rect 30484 236632 30490 236684
rect 58121 236675 58179 236681
rect 58121 236641 58133 236675
rect 58167 236672 58179 236675
rect 60896 236672 60924 236712
rect 62534 236700 62540 236712
rect 62592 236740 62598 236752
rect 70541 236743 70599 236749
rect 70541 236740 70553 236743
rect 62592 236712 70553 236740
rect 62592 236700 62598 236712
rect 70541 236709 70553 236712
rect 70587 236709 70599 236743
rect 70541 236703 70599 236709
rect 70633 236743 70691 236749
rect 70633 236709 70645 236743
rect 70679 236740 70691 236743
rect 72672 236740 72700 236780
rect 77533 236777 77545 236780
rect 77579 236777 77591 236811
rect 77533 236771 77591 236777
rect 89953 236811 90011 236817
rect 89953 236777 89965 236811
rect 89999 236808 90011 236811
rect 96853 236811 96911 236817
rect 96853 236808 96865 236811
rect 89999 236780 96865 236808
rect 89999 236777 90011 236780
rect 89953 236771 90011 236777
rect 96853 236777 96865 236780
rect 96899 236777 96911 236811
rect 96853 236771 96911 236777
rect 70679 236712 72700 236740
rect 70679 236709 70691 236712
rect 70633 236703 70691 236709
rect 58167 236644 60924 236672
rect 77533 236675 77591 236681
rect 58167 236641 58179 236644
rect 58121 236635 58179 236641
rect 77533 236641 77545 236675
rect 77579 236672 77591 236675
rect 80201 236675 80259 236681
rect 80201 236672 80213 236675
rect 77579 236644 80213 236672
rect 77579 236641 77591 236644
rect 77533 236635 77591 236641
rect 80201 236641 80213 236644
rect 80247 236641 80259 236675
rect 80201 236635 80259 236641
rect 80293 236675 80351 236681
rect 80293 236641 80305 236675
rect 80339 236672 80351 236675
rect 89953 236675 90011 236681
rect 89953 236672 89965 236675
rect 80339 236644 89965 236672
rect 80339 236641 80351 236644
rect 80293 236635 80351 236641
rect 89953 236641 89965 236644
rect 89999 236641 90011 236675
rect 89953 236635 90011 236641
rect 106421 236675 106479 236681
rect 106421 236641 106433 236675
rect 106467 236672 106479 236675
rect 107430 236672 107436 236684
rect 106467 236644 107436 236672
rect 106467 236641 106479 236644
rect 106421 236635 106479 236641
rect 107430 236632 107436 236644
rect 107488 236672 107494 236684
rect 146530 236672 146536 236684
rect 107488 236644 146536 236672
rect 107488 236632 107494 236644
rect 146530 236632 146536 236644
rect 146588 236632 146594 236684
rect 23434 236564 23440 236616
rect 23492 236604 23498 236616
rect 26473 236607 26531 236613
rect 26473 236604 26485 236607
rect 23492 236576 26485 236604
rect 23492 236564 23498 236576
rect 26473 236573 26485 236576
rect 26519 236573 26531 236607
rect 48553 236607 48611 236613
rect 48553 236604 48565 236607
rect 26473 236567 26531 236573
rect 48476 236576 48565 236604
rect 48476 236545 48504 236576
rect 48553 236573 48565 236576
rect 48599 236573 48611 236607
rect 48553 236567 48611 236573
rect 72838 236564 72844 236616
rect 72896 236604 72902 236616
rect 121414 236604 121420 236616
rect 72896 236576 121420 236604
rect 72896 236564 72902 236576
rect 121414 236564 121420 236576
rect 121472 236564 121478 236616
rect 208906 236564 208912 236616
rect 208964 236604 208970 236616
rect 218290 236604 218296 236616
rect 208964 236576 218296 236604
rect 208964 236564 208970 236576
rect 218290 236564 218296 236576
rect 218348 236564 218354 236616
rect 48461 236539 48519 236545
rect 48461 236505 48473 236539
rect 48507 236505 48519 236539
rect 48461 236499 48519 236505
rect 48553 236471 48611 236477
rect 48553 236437 48565 236471
rect 48599 236468 48611 236471
rect 58121 236471 58179 236477
rect 58121 236468 58133 236471
rect 48599 236440 58133 236468
rect 48599 236437 48611 236440
rect 48553 236431 48611 236437
rect 58121 236437 58133 236440
rect 58167 236437 58179 236471
rect 58121 236431 58179 236437
rect 29138 235884 29144 235936
rect 29196 235924 29202 235936
rect 82222 235924 82228 235936
rect 29196 235896 82228 235924
rect 29196 235884 29202 235896
rect 82222 235884 82228 235896
rect 82280 235884 82286 235936
rect 86178 235884 86184 235936
rect 86236 235924 86242 235936
rect 99610 235924 99616 235936
rect 86236 235896 99616 235924
rect 86236 235884 86242 235896
rect 99610 235884 99616 235896
rect 99668 235884 99674 235936
rect 136778 235884 136784 235936
rect 136836 235924 136842 235936
rect 169530 235924 169536 235936
rect 136836 235896 169536 235924
rect 136836 235884 136842 235896
rect 169530 235884 169536 235896
rect 169588 235884 169594 235936
rect 63822 235816 63828 235868
rect 63880 235856 63886 235868
rect 166218 235856 166224 235868
rect 63880 235828 166224 235856
rect 63880 235816 63886 235828
rect 166218 235816 166224 235828
rect 166276 235816 166282 235868
rect 114422 235272 114428 235324
rect 114480 235312 114486 235324
rect 159502 235312 159508 235324
rect 114480 235284 159508 235312
rect 114480 235272 114486 235284
rect 159502 235272 159508 235284
rect 159560 235272 159566 235324
rect 173486 235272 173492 235324
rect 173544 235312 173550 235324
rect 174038 235312 174044 235324
rect 173544 235284 174044 235312
rect 173544 235272 173550 235284
rect 174038 235272 174044 235284
rect 174096 235272 174102 235324
rect 47538 235204 47544 235256
rect 47596 235244 47602 235256
rect 65570 235244 65576 235256
rect 47596 235216 65576 235244
rect 47596 235204 47602 235216
rect 65570 235204 65576 235216
rect 65628 235204 65634 235256
rect 156834 235204 156840 235256
rect 156892 235244 156898 235256
rect 215714 235244 215720 235256
rect 156892 235216 215720 235244
rect 156892 235204 156898 235216
rect 215714 235204 215720 235216
rect 215772 235204 215778 235256
rect 37418 235136 37424 235188
rect 37476 235176 37482 235188
rect 75506 235176 75512 235188
rect 37476 235148 75512 235176
rect 37476 235136 37482 235148
rect 75506 235136 75512 235148
rect 75564 235136 75570 235188
rect 146530 235136 146536 235188
rect 146588 235176 146594 235188
rect 216910 235176 216916 235188
rect 146588 235148 216916 235176
rect 146588 235136 146594 235148
rect 216910 235136 216916 235148
rect 216968 235136 216974 235188
rect 135398 233912 135404 233964
rect 135456 233952 135462 233964
rect 142298 233952 142304 233964
rect 135456 233924 142304 233952
rect 135456 233912 135462 233924
rect 142298 233912 142304 233924
rect 142356 233912 142362 233964
rect 49930 233776 49936 233828
rect 49988 233816 49994 233828
rect 58118 233816 58124 233828
rect 49988 233788 58124 233816
rect 49988 233776 49994 233788
rect 58118 233776 58124 233788
rect 58176 233776 58182 233828
rect 177166 233708 177172 233760
rect 177224 233748 177230 233760
rect 185078 233748 185084 233760
rect 177224 233720 185084 233748
rect 177224 233708 177230 233720
rect 185078 233708 185084 233720
rect 185136 233708 185142 233760
rect 92710 233028 92716 233080
rect 92768 233068 92774 233080
rect 100990 233068 100996 233080
rect 92768 233040 100996 233068
rect 92768 233028 92774 233040
rect 100990 233028 100996 233040
rect 101048 233028 101054 233080
rect 135398 232688 135404 232740
rect 135456 232728 135462 232740
rect 142206 232728 142212 232740
rect 135456 232700 142212 232728
rect 135456 232688 135462 232700
rect 142206 232688 142212 232700
rect 142264 232688 142270 232740
rect 134294 232620 134300 232672
rect 134352 232660 134358 232672
rect 142298 232660 142304 232672
rect 134352 232632 142304 232660
rect 134352 232620 134358 232632
rect 142298 232620 142304 232632
rect 142356 232620 142362 232672
rect 51218 232484 51224 232536
rect 51276 232524 51282 232536
rect 58026 232524 58032 232536
rect 51276 232496 58032 232524
rect 51276 232484 51282 232496
rect 58026 232484 58032 232496
rect 58084 232484 58090 232536
rect 182318 232484 182324 232536
rect 182376 232524 182382 232536
rect 185262 232524 185268 232536
rect 182376 232496 185268 232524
rect 182376 232484 182382 232496
rect 185262 232484 185268 232496
rect 185320 232484 185326 232536
rect 50574 232416 50580 232468
rect 50632 232456 50638 232468
rect 58118 232456 58124 232468
rect 50632 232428 58124 232456
rect 50632 232416 50638 232428
rect 58118 232416 58124 232428
rect 58176 232416 58182 232468
rect 100990 232456 100996 232468
rect 98156 232428 100996 232456
rect 93998 232348 94004 232400
rect 94056 232388 94062 232400
rect 98156 232388 98184 232428
rect 100990 232416 100996 232428
rect 101048 232416 101054 232468
rect 185170 232456 185176 232468
rect 182336 232428 185176 232456
rect 94056 232360 98184 232388
rect 94056 232348 94062 232360
rect 177718 232348 177724 232400
rect 177776 232388 177782 232400
rect 182336 232388 182364 232428
rect 185170 232416 185176 232428
rect 185228 232416 185234 232468
rect 177776 232360 182364 232388
rect 177776 232348 177782 232360
rect 218290 232348 218296 232400
rect 218348 232388 218354 232400
rect 222338 232388 222344 232400
rect 218348 232360 222344 232388
rect 218348 232348 218354 232360
rect 222338 232348 222344 232360
rect 222396 232348 222402 232400
rect 177718 231804 177724 231856
rect 177776 231844 177782 231856
rect 182318 231844 182324 231856
rect 177776 231816 182324 231844
rect 177776 231804 177782 231816
rect 182318 231804 182324 231816
rect 182376 231804 182382 231856
rect 92710 231668 92716 231720
rect 92768 231708 92774 231720
rect 100990 231708 100996 231720
rect 92768 231680 100996 231708
rect 92768 231668 92774 231680
rect 100990 231668 100996 231680
rect 101048 231668 101054 231720
rect 134846 231464 134852 231516
rect 134904 231504 134910 231516
rect 139630 231504 139636 231516
rect 134904 231476 139636 231504
rect 134904 231464 134910 231476
rect 139630 231464 139636 231476
rect 139688 231464 139694 231516
rect 51218 231328 51224 231380
rect 51276 231368 51282 231380
rect 56738 231368 56744 231380
rect 51276 231340 56744 231368
rect 51276 231328 51282 231340
rect 56738 231328 56744 231340
rect 56796 231328 56802 231380
rect 51126 231192 51132 231244
rect 51184 231232 51190 231244
rect 51184 231204 56784 231232
rect 51184 231192 51190 231204
rect 51218 231056 51224 231108
rect 51276 231096 51282 231108
rect 52690 231096 52696 231108
rect 51276 231068 52696 231096
rect 51276 231056 51282 231068
rect 52690 231056 52696 231068
rect 52748 231056 52754 231108
rect 56756 230960 56784 231204
rect 95378 231124 95384 231176
rect 95436 231164 95442 231176
rect 100990 231164 100996 231176
rect 95436 231136 100996 231164
rect 95436 231124 95442 231136
rect 100990 231124 100996 231136
rect 101048 231124 101054 231176
rect 135306 231056 135312 231108
rect 135364 231096 135370 231108
rect 136870 231096 136876 231108
rect 135364 231068 136876 231096
rect 135364 231056 135370 231068
rect 136870 231056 136876 231068
rect 136928 231056 136934 231108
rect 178270 231056 178276 231108
rect 178328 231096 178334 231108
rect 185262 231096 185268 231108
rect 178328 231068 185268 231096
rect 178328 231056 178334 231068
rect 185262 231056 185268 231068
rect 185320 231056 185326 231108
rect 94090 230988 94096 231040
rect 94148 231028 94154 231040
rect 101082 231028 101088 231040
rect 94148 231000 101088 231028
rect 94148 230988 94154 231000
rect 101082 230988 101088 231000
rect 101140 230988 101146 231040
rect 135398 230988 135404 231040
rect 135456 231028 135462 231040
rect 185170 231028 185176 231040
rect 135456 231000 139676 231028
rect 135456 230988 135462 231000
rect 58210 230960 58216 230972
rect 56756 230932 58216 230960
rect 58210 230920 58216 230932
rect 58268 230920 58274 230972
rect 92710 230852 92716 230904
rect 92768 230892 92774 230904
rect 95378 230892 95384 230904
rect 92768 230864 95384 230892
rect 92768 230852 92774 230864
rect 95378 230852 95384 230864
rect 95436 230852 95442 230904
rect 139648 230892 139676 231000
rect 178288 231000 185176 231028
rect 177718 230920 177724 230972
rect 177776 230960 177782 230972
rect 178288 230960 178316 231000
rect 185170 230988 185176 231000
rect 185228 230988 185234 231040
rect 177776 230932 178316 230960
rect 177776 230920 177782 230932
rect 143678 230892 143684 230904
rect 139648 230864 143684 230892
rect 143678 230852 143684 230864
rect 143736 230852 143742 230904
rect 56738 230716 56744 230768
rect 56796 230756 56802 230768
rect 58302 230756 58308 230768
rect 56796 230728 58308 230756
rect 56796 230716 56802 230728
rect 58302 230716 58308 230728
rect 58360 230716 58366 230768
rect 139630 230580 139636 230632
rect 139688 230620 139694 230632
rect 142942 230620 142948 230632
rect 139688 230592 142948 230620
rect 139688 230580 139694 230592
rect 142942 230580 142948 230592
rect 143000 230580 143006 230632
rect 135306 229968 135312 230020
rect 135364 230008 135370 230020
rect 139630 230008 139636 230020
rect 135364 229980 139636 230008
rect 135364 229968 135370 229980
rect 139630 229968 139636 229980
rect 139688 229968 139694 230020
rect 51218 229832 51224 229884
rect 51276 229872 51282 229884
rect 56462 229872 56468 229884
rect 51276 229844 56468 229872
rect 51276 229832 51282 229844
rect 56462 229832 56468 229844
rect 56520 229832 56526 229884
rect 51126 229696 51132 229748
rect 51184 229736 51190 229748
rect 56186 229736 56192 229748
rect 51184 229708 56192 229736
rect 51184 229696 51190 229708
rect 56186 229696 56192 229708
rect 56244 229696 56250 229748
rect 135398 229628 135404 229680
rect 135456 229668 135462 229680
rect 135456 229640 139676 229668
rect 135456 229628 135462 229640
rect 52690 229560 52696 229612
rect 52748 229600 52754 229612
rect 58210 229600 58216 229612
rect 52748 229572 58216 229600
rect 52748 229560 52754 229572
rect 58210 229560 58216 229572
rect 58268 229560 58274 229612
rect 92710 229560 92716 229612
rect 92768 229600 92774 229612
rect 101082 229600 101088 229612
rect 92768 229572 101088 229600
rect 92768 229560 92774 229572
rect 101082 229560 101088 229572
rect 101140 229560 101146 229612
rect 139648 229600 139676 229640
rect 143586 229600 143592 229612
rect 139648 229572 143592 229600
rect 143586 229560 143592 229572
rect 143644 229560 143650 229612
rect 177626 229560 177632 229612
rect 177684 229600 177690 229612
rect 185262 229600 185268 229612
rect 177684 229572 185268 229600
rect 177684 229560 177690 229572
rect 185262 229560 185268 229572
rect 185320 229560 185326 229612
rect 93170 229492 93176 229544
rect 93228 229532 93234 229544
rect 100990 229532 100996 229544
rect 93228 229504 100996 229532
rect 93228 229492 93234 229504
rect 100990 229492 100996 229504
rect 101048 229492 101054 229544
rect 136870 229492 136876 229544
rect 136928 229532 136934 229544
rect 143678 229532 143684 229544
rect 136928 229504 143684 229532
rect 136928 229492 136934 229504
rect 143678 229492 143684 229504
rect 143736 229492 143742 229544
rect 177810 229492 177816 229544
rect 177868 229532 177874 229544
rect 185170 229532 185176 229544
rect 177868 229504 185176 229532
rect 177868 229492 177874 229504
rect 185170 229492 185176 229504
rect 185228 229492 185234 229544
rect 139630 229424 139636 229476
rect 139688 229464 139694 229476
rect 143494 229464 143500 229476
rect 139688 229436 143500 229464
rect 139688 229424 139694 229436
rect 143494 229424 143500 229436
rect 143552 229424 143558 229476
rect 177718 229424 177724 229476
rect 177776 229464 177782 229476
rect 185354 229464 185360 229476
rect 177776 229436 185360 229464
rect 177776 229424 177782 229436
rect 185354 229424 185360 229436
rect 185412 229424 185418 229476
rect 56186 229288 56192 229340
rect 56244 229328 56250 229340
rect 58210 229328 58216 229340
rect 56244 229300 58216 229328
rect 56244 229288 56250 229300
rect 58210 229288 58216 229300
rect 58268 229288 58274 229340
rect 56462 229016 56468 229068
rect 56520 229056 56526 229068
rect 58302 229056 58308 229068
rect 56520 229028 58308 229056
rect 56520 229016 56526 229028
rect 58302 229016 58308 229028
rect 58360 229016 58366 229068
rect 92710 228880 92716 228932
rect 92768 228920 92774 228932
rect 100990 228920 100996 228932
rect 92768 228892 100996 228920
rect 92768 228880 92774 228892
rect 100990 228880 100996 228892
rect 101048 228880 101054 228932
rect 50758 228472 50764 228524
rect 50816 228512 50822 228524
rect 55450 228512 55456 228524
rect 50816 228484 55456 228512
rect 50816 228472 50822 228484
rect 55450 228472 55456 228484
rect 55508 228472 55514 228524
rect 135398 228404 135404 228456
rect 135456 228444 135462 228456
rect 135456 228416 140228 228444
rect 135456 228404 135462 228416
rect 51126 228336 51132 228388
rect 51184 228376 51190 228388
rect 51184 228348 52828 228376
rect 51184 228336 51190 228348
rect 51218 228268 51224 228320
rect 51276 228308 51282 228320
rect 52690 228308 52696 228320
rect 51276 228280 52696 228308
rect 51276 228268 51282 228280
rect 52690 228268 52696 228280
rect 52748 228268 52754 228320
rect 52800 228308 52828 228348
rect 135306 228336 135312 228388
rect 135364 228376 135370 228388
rect 135364 228348 140136 228376
rect 135364 228336 135370 228348
rect 52800 228280 55496 228308
rect 55468 228240 55496 228280
rect 135398 228268 135404 228320
rect 135456 228308 135462 228320
rect 138158 228308 138164 228320
rect 135456 228280 138164 228308
rect 135456 228268 135462 228280
rect 138158 228268 138164 228280
rect 138216 228268 138222 228320
rect 58210 228240 58216 228252
rect 55468 228212 58216 228240
rect 58210 228200 58216 228212
rect 58268 228200 58274 228252
rect 93170 228200 93176 228252
rect 93228 228240 93234 228252
rect 101082 228240 101088 228252
rect 93228 228212 101088 228240
rect 93228 228200 93234 228212
rect 101082 228200 101088 228212
rect 101140 228200 101146 228252
rect 92710 228132 92716 228184
rect 92768 228172 92774 228184
rect 100990 228172 100996 228184
rect 92768 228144 100996 228172
rect 92768 228132 92774 228144
rect 100990 228132 100996 228144
rect 101048 228132 101054 228184
rect 140108 228172 140136 228348
rect 140200 228240 140228 228416
rect 181122 228268 181128 228320
rect 181180 228308 181186 228320
rect 185170 228308 185176 228320
rect 181180 228280 185176 228308
rect 181180 228268 181186 228280
rect 185170 228268 185176 228280
rect 185228 228268 185234 228320
rect 143678 228240 143684 228252
rect 140200 228212 143684 228240
rect 143678 228200 143684 228212
rect 143736 228200 143742 228252
rect 177718 228200 177724 228252
rect 177776 228240 177782 228252
rect 185630 228240 185636 228252
rect 177776 228212 185636 228240
rect 177776 228200 177782 228212
rect 185630 228200 185636 228212
rect 185688 228200 185694 228252
rect 143310 228172 143316 228184
rect 140108 228144 143316 228172
rect 143310 228132 143316 228144
rect 143368 228132 143374 228184
rect 177626 228132 177632 228184
rect 177684 228172 177690 228184
rect 185906 228172 185912 228184
rect 177684 228144 185912 228172
rect 177684 228132 177690 228144
rect 185906 228132 185912 228144
rect 185964 228132 185970 228184
rect 55450 227860 55456 227912
rect 55508 227900 55514 227912
rect 58302 227900 58308 227912
rect 55508 227872 58308 227900
rect 55508 227860 55514 227872
rect 58302 227860 58308 227872
rect 58360 227860 58366 227912
rect 50942 227248 50948 227300
rect 51000 227288 51006 227300
rect 56738 227288 56744 227300
rect 51000 227260 56744 227288
rect 51000 227248 51006 227260
rect 56738 227248 56744 227260
rect 56796 227248 56802 227300
rect 135398 226840 135404 226892
rect 135456 226880 135462 226892
rect 135456 226852 139676 226880
rect 135456 226840 135462 226852
rect 52690 226772 52696 226824
rect 52748 226812 52754 226824
rect 58210 226812 58216 226824
rect 52748 226784 58216 226812
rect 52748 226772 52754 226784
rect 58210 226772 58216 226784
rect 58268 226772 58274 226824
rect 93630 226772 93636 226824
rect 93688 226812 93694 226824
rect 100990 226812 100996 226824
rect 93688 226784 100996 226812
rect 93688 226772 93694 226784
rect 100990 226772 100996 226784
rect 101048 226772 101054 226824
rect 139648 226812 139676 226852
rect 182318 226840 182324 226892
rect 182376 226880 182382 226892
rect 185262 226880 185268 226892
rect 182376 226852 185268 226880
rect 182376 226840 182382 226852
rect 185262 226840 185268 226852
rect 185320 226840 185326 226892
rect 143310 226812 143316 226824
rect 139648 226784 143316 226812
rect 143310 226772 143316 226784
rect 143368 226772 143374 226824
rect 177626 226772 177632 226824
rect 177684 226812 177690 226824
rect 185170 226812 185176 226824
rect 177684 226784 185176 226812
rect 177684 226772 177690 226784
rect 185170 226772 185176 226784
rect 185228 226772 185234 226824
rect 92710 226704 92716 226756
rect 92768 226744 92774 226756
rect 101082 226744 101088 226756
rect 92768 226716 101088 226744
rect 92768 226704 92774 226716
rect 101082 226704 101088 226716
rect 101140 226704 101146 226756
rect 138158 226704 138164 226756
rect 138216 226744 138222 226756
rect 143678 226744 143684 226756
rect 138216 226716 143684 226744
rect 138216 226704 138222 226716
rect 143678 226704 143684 226716
rect 143736 226704 143742 226756
rect 56738 226636 56744 226688
rect 56796 226676 56802 226688
rect 58302 226676 58308 226688
rect 56796 226648 58308 226676
rect 56796 226636 56802 226648
rect 58302 226636 58308 226648
rect 58360 226636 58366 226688
rect 177718 226636 177724 226688
rect 177776 226676 177782 226688
rect 181122 226676 181128 226688
rect 177776 226648 181128 226676
rect 177776 226636 177782 226648
rect 181122 226636 181128 226648
rect 181180 226636 181186 226688
rect 50482 225548 50488 225600
rect 50540 225588 50546 225600
rect 58394 225588 58400 225600
rect 50540 225560 58400 225588
rect 50540 225548 50546 225560
rect 58394 225548 58400 225560
rect 58452 225548 58458 225600
rect 134570 225548 134576 225600
rect 134628 225588 134634 225600
rect 143494 225588 143500 225600
rect 134628 225560 143500 225588
rect 134628 225548 134634 225560
rect 143494 225548 143500 225560
rect 143552 225548 143558 225600
rect 50758 225480 50764 225532
rect 50816 225520 50822 225532
rect 58302 225520 58308 225532
rect 50816 225492 58308 225520
rect 50816 225480 50822 225492
rect 58302 225480 58308 225492
rect 58360 225480 58366 225532
rect 135214 225480 135220 225532
rect 135272 225520 135278 225532
rect 143586 225520 143592 225532
rect 135272 225492 143592 225520
rect 135272 225480 135278 225492
rect 143586 225480 143592 225492
rect 143644 225480 143650 225532
rect 51310 225412 51316 225464
rect 51368 225452 51374 225464
rect 58210 225452 58216 225464
rect 51368 225424 58216 225452
rect 51368 225412 51374 225424
rect 58210 225412 58216 225424
rect 58268 225412 58274 225464
rect 92802 225412 92808 225464
rect 92860 225452 92866 225464
rect 101082 225452 101088 225464
rect 92860 225424 101088 225452
rect 92860 225412 92866 225424
rect 101082 225412 101088 225424
rect 101140 225412 101146 225464
rect 135490 225412 135496 225464
rect 135548 225452 135554 225464
rect 143678 225452 143684 225464
rect 135548 225424 143684 225452
rect 135548 225412 135554 225424
rect 143678 225412 143684 225424
rect 143736 225412 143742 225464
rect 177626 225412 177632 225464
rect 177684 225452 177690 225464
rect 185170 225452 185176 225464
rect 177684 225424 185176 225452
rect 177684 225412 177690 225424
rect 185170 225412 185176 225424
rect 185228 225412 185234 225464
rect 92894 225344 92900 225396
rect 92952 225384 92958 225396
rect 100990 225384 100996 225396
rect 92952 225356 100996 225384
rect 92952 225344 92958 225356
rect 100990 225344 100996 225356
rect 101048 225344 101054 225396
rect 177810 225344 177816 225396
rect 177868 225384 177874 225396
rect 185262 225384 185268 225396
rect 177868 225356 185268 225384
rect 177868 225344 177874 225356
rect 185262 225344 185268 225356
rect 185320 225344 185326 225396
rect 92710 225276 92716 225328
rect 92768 225316 92774 225328
rect 101174 225316 101180 225328
rect 92768 225288 101180 225316
rect 92768 225276 92774 225288
rect 101174 225276 101180 225288
rect 101232 225276 101238 225328
rect 177718 225276 177724 225328
rect 177776 225316 177782 225328
rect 182318 225316 182324 225328
rect 177776 225288 182324 225316
rect 177776 225276 177782 225288
rect 182318 225276 182324 225288
rect 182376 225276 182382 225328
rect 51034 224256 51040 224308
rect 51092 224296 51098 224308
rect 52690 224296 52696 224308
rect 51092 224268 52696 224296
rect 51092 224256 51098 224268
rect 52690 224256 52696 224268
rect 52748 224256 52754 224308
rect 135214 224256 135220 224308
rect 135272 224296 135278 224308
rect 136870 224296 136876 224308
rect 135272 224268 136876 224296
rect 135272 224256 135278 224268
rect 136870 224256 136876 224268
rect 136928 224256 136934 224308
rect 51126 224188 51132 224240
rect 51184 224228 51190 224240
rect 51184 224200 56784 224228
rect 51184 224188 51190 224200
rect 51218 224120 51224 224172
rect 51276 224160 51282 224172
rect 51276 224132 56692 224160
rect 51276 224120 51282 224132
rect 56664 224024 56692 224132
rect 56756 224092 56784 224200
rect 135306 224188 135312 224240
rect 135364 224228 135370 224240
rect 135364 224200 139860 224228
rect 135364 224188 135370 224200
rect 135398 224120 135404 224172
rect 135456 224160 135462 224172
rect 135456 224132 139768 224160
rect 135456 224120 135462 224132
rect 58210 224092 58216 224104
rect 56756 224064 58216 224092
rect 58210 224052 58216 224064
rect 58268 224052 58274 224104
rect 93906 224052 93912 224104
rect 93964 224092 93970 224104
rect 100990 224092 100996 224104
rect 93964 224064 100996 224092
rect 93964 224052 93970 224064
rect 100990 224052 100996 224064
rect 101048 224052 101054 224104
rect 58302 224024 58308 224036
rect 56664 223996 58308 224024
rect 58302 223984 58308 223996
rect 58360 223984 58366 224036
rect 93722 223984 93728 224036
rect 93780 224024 93786 224036
rect 101082 224024 101088 224036
rect 93780 223996 101088 224024
rect 93780 223984 93786 223996
rect 101082 223984 101088 223996
rect 101140 223984 101146 224036
rect 139740 224024 139768 224132
rect 139832 224092 139860 224200
rect 143678 224092 143684 224104
rect 139832 224064 143684 224092
rect 143678 224052 143684 224064
rect 143736 224052 143742 224104
rect 177718 224052 177724 224104
rect 177776 224092 177782 224104
rect 185354 224092 185360 224104
rect 177776 224064 185360 224092
rect 177776 224052 177782 224064
rect 185354 224052 185360 224064
rect 185412 224052 185418 224104
rect 143310 224024 143316 224036
rect 139740 223996 143316 224024
rect 143310 223984 143316 223996
rect 143368 223984 143374 224036
rect 177350 223984 177356 224036
rect 177408 224024 177414 224036
rect 185170 224024 185176 224036
rect 177408 223996 185176 224024
rect 177408 223984 177414 223996
rect 185170 223984 185176 223996
rect 185228 223984 185234 224036
rect 50942 223168 50948 223220
rect 51000 223208 51006 223220
rect 56278 223208 56284 223220
rect 51000 223180 56284 223208
rect 51000 223168 51006 223180
rect 56278 223168 56284 223180
rect 56336 223168 56342 223220
rect 51218 223032 51224 223084
rect 51276 223072 51282 223084
rect 52782 223072 52788 223084
rect 51276 223044 52788 223072
rect 51276 223032 51282 223044
rect 52782 223032 52788 223044
rect 52840 223032 52846 223084
rect 135306 223032 135312 223084
rect 135364 223072 135370 223084
rect 137606 223072 137612 223084
rect 135364 223044 137612 223072
rect 135364 223032 135370 223044
rect 137606 223032 137612 223044
rect 137664 223032 137670 223084
rect 135398 222760 135404 222812
rect 135456 222800 135462 222812
rect 135456 222772 139676 222800
rect 135456 222760 135462 222772
rect 52690 222692 52696 222744
rect 52748 222732 52754 222744
rect 58210 222732 58216 222744
rect 52748 222704 58216 222732
rect 52748 222692 52754 222704
rect 58210 222692 58216 222704
rect 58268 222692 58274 222744
rect 92710 222692 92716 222744
rect 92768 222732 92774 222744
rect 101450 222732 101456 222744
rect 92768 222704 101456 222732
rect 92768 222692 92774 222704
rect 101450 222692 101456 222704
rect 101508 222692 101514 222744
rect 139648 222732 139676 222772
rect 143310 222732 143316 222744
rect 139648 222704 143316 222732
rect 143310 222692 143316 222704
rect 143368 222692 143374 222744
rect 177626 222692 177632 222744
rect 177684 222732 177690 222744
rect 185170 222732 185176 222744
rect 177684 222704 185176 222732
rect 177684 222692 177690 222704
rect 185170 222692 185176 222704
rect 185228 222692 185234 222744
rect 92986 222624 92992 222676
rect 93044 222664 93050 222676
rect 101542 222664 101548 222676
rect 93044 222636 101548 222664
rect 93044 222624 93050 222636
rect 101542 222624 101548 222636
rect 101600 222624 101606 222676
rect 136870 222624 136876 222676
rect 136928 222664 136934 222676
rect 143678 222664 143684 222676
rect 136928 222636 143684 222664
rect 136928 222624 136934 222636
rect 143678 222624 143684 222636
rect 143736 222624 143742 222676
rect 177718 222624 177724 222676
rect 177776 222664 177782 222676
rect 185262 222664 185268 222676
rect 177776 222636 185268 222664
rect 177776 222624 177782 222636
rect 185262 222624 185268 222636
rect 185320 222624 185326 222676
rect 56278 222420 56284 222472
rect 56336 222460 56342 222472
rect 58302 222460 58308 222472
rect 56336 222432 58308 222460
rect 56336 222420 56342 222432
rect 58302 222420 58308 222432
rect 58360 222420 58366 222472
rect 134846 222352 134852 222404
rect 134904 222392 134910 222404
rect 139722 222392 139728 222404
rect 134904 222364 139728 222392
rect 134904 222352 134910 222364
rect 139722 222352 139728 222364
rect 139780 222352 139786 222404
rect 134478 221808 134484 221860
rect 134536 221848 134542 221860
rect 139630 221848 139636 221860
rect 134536 221820 139636 221848
rect 134536 221808 134542 221820
rect 139630 221808 139636 221820
rect 139688 221808 139694 221860
rect 51218 221672 51224 221724
rect 51276 221712 51282 221724
rect 56738 221712 56744 221724
rect 51276 221684 56744 221712
rect 51276 221672 51282 221684
rect 56738 221672 56744 221684
rect 56796 221672 56802 221724
rect 51126 221536 51132 221588
rect 51184 221576 51190 221588
rect 55910 221576 55916 221588
rect 51184 221548 55916 221576
rect 51184 221536 51190 221548
rect 55910 221536 55916 221548
rect 55968 221536 55974 221588
rect 51218 221400 51224 221452
rect 51276 221440 51282 221452
rect 52690 221440 52696 221452
rect 51276 221412 52696 221440
rect 51276 221400 51282 221412
rect 52690 221400 52696 221412
rect 52748 221400 52754 221452
rect 135306 221400 135312 221452
rect 135364 221440 135370 221452
rect 136870 221440 136876 221452
rect 135364 221412 136876 221440
rect 135364 221400 135370 221412
rect 136870 221400 136876 221412
rect 136928 221400 136934 221452
rect 52782 221264 52788 221316
rect 52840 221304 52846 221316
rect 58210 221304 58216 221316
rect 52840 221276 58216 221304
rect 52840 221264 52846 221276
rect 58210 221264 58216 221276
rect 58268 221264 58274 221316
rect 93170 221264 93176 221316
rect 93228 221304 93234 221316
rect 101726 221304 101732 221316
rect 93228 221276 101732 221304
rect 93228 221264 93234 221276
rect 101726 221264 101732 221276
rect 101784 221264 101790 221316
rect 137606 221264 137612 221316
rect 137664 221304 137670 221316
rect 143678 221304 143684 221316
rect 137664 221276 143684 221304
rect 137664 221264 137670 221276
rect 143678 221264 143684 221276
rect 143736 221264 143742 221316
rect 177626 221264 177632 221316
rect 177684 221304 177690 221316
rect 185262 221304 185268 221316
rect 177684 221276 185268 221304
rect 177684 221264 177690 221276
rect 185262 221264 185268 221276
rect 185320 221264 185326 221316
rect 93722 221196 93728 221248
rect 93780 221236 93786 221248
rect 101542 221236 101548 221248
rect 93780 221208 101548 221236
rect 93780 221196 93786 221208
rect 101542 221196 101548 221208
rect 101600 221196 101606 221248
rect 177810 221196 177816 221248
rect 177868 221236 177874 221248
rect 185170 221236 185176 221248
rect 177868 221208 185176 221236
rect 177868 221196 177874 221208
rect 185170 221196 185176 221208
rect 185228 221196 185234 221248
rect 92710 221128 92716 221180
rect 92768 221168 92774 221180
rect 101266 221168 101272 221180
rect 92768 221140 101272 221168
rect 92768 221128 92774 221140
rect 101266 221128 101272 221140
rect 101324 221128 101330 221180
rect 139722 221128 139728 221180
rect 139780 221168 139786 221180
rect 143586 221168 143592 221180
rect 139780 221140 143592 221168
rect 139780 221128 139786 221140
rect 143586 221128 143592 221140
rect 143644 221128 143650 221180
rect 177718 221128 177724 221180
rect 177776 221168 177782 221180
rect 185446 221168 185452 221180
rect 177776 221140 185452 221168
rect 177776 221128 177782 221140
rect 185446 221128 185452 221140
rect 185504 221128 185510 221180
rect 55910 220992 55916 221044
rect 55968 221032 55974 221044
rect 58210 221032 58216 221044
rect 55968 221004 58216 221032
rect 55968 220992 55974 221004
rect 58210 220992 58216 221004
rect 58268 220992 58274 221044
rect 56738 220856 56744 220908
rect 56796 220896 56802 220908
rect 58302 220896 58308 220908
rect 56796 220868 58308 220896
rect 56796 220856 56802 220868
rect 58302 220856 58308 220868
rect 58360 220856 58366 220908
rect 139630 220584 139636 220636
rect 139688 220624 139694 220636
rect 143678 220624 143684 220636
rect 139688 220596 143684 220624
rect 139688 220584 139694 220596
rect 143678 220584 143684 220596
rect 143736 220584 143742 220636
rect 50942 220312 50948 220364
rect 51000 220352 51006 220364
rect 56462 220352 56468 220364
rect 51000 220324 56468 220352
rect 51000 220312 51006 220324
rect 56462 220312 56468 220324
rect 56520 220312 56526 220364
rect 135306 220108 135312 220160
rect 135364 220148 135370 220160
rect 138158 220148 138164 220160
rect 135364 220120 138164 220148
rect 135364 220108 135370 220120
rect 138158 220108 138164 220120
rect 138216 220108 138222 220160
rect 50206 219972 50212 220024
rect 50264 220012 50270 220024
rect 52782 220012 52788 220024
rect 50264 219984 52788 220012
rect 50264 219972 50270 219984
rect 52782 219972 52788 219984
rect 52840 219972 52846 220024
rect 135398 219972 135404 220024
rect 135456 220012 135462 220024
rect 135456 219984 139676 220012
rect 135456 219972 135462 219984
rect 52690 219904 52696 219956
rect 52748 219944 52754 219956
rect 58210 219944 58216 219956
rect 52748 219916 58216 219944
rect 52748 219904 52754 219916
rect 58210 219904 58216 219916
rect 58268 219904 58274 219956
rect 92710 219904 92716 219956
rect 92768 219944 92774 219956
rect 101818 219944 101824 219956
rect 92768 219916 101824 219944
rect 92768 219904 92774 219916
rect 101818 219904 101824 219916
rect 101876 219904 101882 219956
rect 139648 219944 139676 219984
rect 143126 219944 143132 219956
rect 139648 219916 143132 219944
rect 143126 219904 143132 219916
rect 143184 219904 143190 219956
rect 177626 219904 177632 219956
rect 177684 219944 177690 219956
rect 185170 219944 185176 219956
rect 177684 219916 185176 219944
rect 177684 219904 177690 219916
rect 185170 219904 185176 219916
rect 185228 219904 185234 219956
rect 92802 219836 92808 219888
rect 92860 219876 92866 219888
rect 101726 219876 101732 219888
rect 92860 219848 101732 219876
rect 92860 219836 92866 219848
rect 101726 219836 101732 219848
rect 101784 219836 101790 219888
rect 136870 219836 136876 219888
rect 136928 219876 136934 219888
rect 143678 219876 143684 219888
rect 136928 219848 143684 219876
rect 136928 219836 136934 219848
rect 143678 219836 143684 219848
rect 143736 219836 143742 219888
rect 177718 219836 177724 219888
rect 177776 219876 177782 219888
rect 185354 219876 185360 219888
rect 177776 219848 185360 219876
rect 177776 219836 177782 219848
rect 185354 219836 185360 219848
rect 185412 219836 185418 219888
rect 56462 219496 56468 219548
rect 56520 219536 56526 219548
rect 58302 219536 58308 219548
rect 56520 219508 58308 219536
rect 56520 219496 56526 219508
rect 58302 219496 58308 219508
rect 58360 219496 58366 219548
rect 50206 218884 50212 218936
rect 50264 218924 50270 218936
rect 53058 218924 53064 218936
rect 50264 218896 53064 218924
rect 50264 218884 50270 218896
rect 53058 218884 53064 218896
rect 53116 218884 53122 218936
rect 135030 218816 135036 218868
rect 135088 218856 135094 218868
rect 137514 218856 137520 218868
rect 135088 218828 137520 218856
rect 135088 218816 135094 218828
rect 137514 218816 137520 218828
rect 137572 218816 137578 218868
rect 51218 218680 51224 218732
rect 51276 218720 51282 218732
rect 52690 218720 52696 218732
rect 51276 218692 52696 218720
rect 51276 218680 51282 218692
rect 52690 218680 52696 218692
rect 52748 218680 52754 218732
rect 135398 218680 135404 218732
rect 135456 218720 135462 218732
rect 135456 218692 140228 218720
rect 135456 218680 135462 218692
rect 50850 218612 50856 218664
rect 50908 218652 50914 218664
rect 55450 218652 55456 218664
rect 50908 218624 55456 218652
rect 50908 218612 50914 218624
rect 55450 218612 55456 218624
rect 55508 218612 55514 218664
rect 135306 218612 135312 218664
rect 135364 218652 135370 218664
rect 137974 218652 137980 218664
rect 135364 218624 137980 218652
rect 135364 218612 135370 218624
rect 137974 218612 137980 218624
rect 138032 218612 138038 218664
rect 52782 218544 52788 218596
rect 52840 218584 52846 218596
rect 58210 218584 58216 218596
rect 52840 218556 58216 218584
rect 52840 218544 52846 218556
rect 58210 218544 58216 218556
rect 58268 218544 58274 218596
rect 92802 218544 92808 218596
rect 92860 218584 92866 218596
rect 101910 218584 101916 218596
rect 92860 218556 101916 218584
rect 92860 218544 92866 218556
rect 101910 218544 101916 218556
rect 101968 218544 101974 218596
rect 140200 218584 140228 218692
rect 185814 218612 185820 218664
rect 185872 218652 185878 218664
rect 185998 218652 186004 218664
rect 185872 218624 186004 218652
rect 185872 218612 185878 218624
rect 185998 218612 186004 218624
rect 186056 218612 186062 218664
rect 143494 218584 143500 218596
rect 140200 218556 143500 218584
rect 143494 218544 143500 218556
rect 143552 218544 143558 218596
rect 177718 218544 177724 218596
rect 177776 218584 177782 218596
rect 185538 218584 185544 218596
rect 177776 218556 185544 218584
rect 177776 218544 177782 218556
rect 185538 218544 185544 218556
rect 185596 218544 185602 218596
rect 93722 218476 93728 218528
rect 93780 218516 93786 218528
rect 101726 218516 101732 218528
rect 93780 218488 101732 218516
rect 93780 218476 93786 218488
rect 101726 218476 101732 218488
rect 101784 218476 101790 218528
rect 138158 218476 138164 218528
rect 138216 218516 138222 218528
rect 143678 218516 143684 218528
rect 138216 218488 143684 218516
rect 138216 218476 138222 218488
rect 143678 218476 143684 218488
rect 143736 218476 143742 218528
rect 177626 218476 177632 218528
rect 177684 218516 177690 218528
rect 185722 218516 185728 218528
rect 177684 218488 185728 218516
rect 177684 218476 177690 218488
rect 185722 218476 185728 218488
rect 185780 218476 185786 218528
rect 55450 218000 55456 218052
rect 55508 218040 55514 218052
rect 58210 218040 58216 218052
rect 55508 218012 58216 218040
rect 55508 218000 55514 218012
rect 58210 218000 58216 218012
rect 58268 218000 58274 218052
rect 51218 217456 51224 217508
rect 51276 217496 51282 217508
rect 52874 217496 52880 217508
rect 51276 217468 52880 217496
rect 51276 217456 51282 217468
rect 52874 217456 52880 217468
rect 52932 217456 52938 217508
rect 135398 217456 135404 217508
rect 135456 217496 135462 217508
rect 137698 217496 137704 217508
rect 135456 217468 137704 217496
rect 135456 217456 135462 217468
rect 137698 217456 137704 217468
rect 137756 217456 137762 217508
rect 51218 217320 51224 217372
rect 51276 217360 51282 217372
rect 52782 217360 52788 217372
rect 51276 217332 52788 217360
rect 51276 217320 51282 217332
rect 52782 217320 52788 217332
rect 52840 217320 52846 217372
rect 135398 217320 135404 217372
rect 135456 217360 135462 217372
rect 137606 217360 137612 217372
rect 135456 217332 137612 217360
rect 135456 217320 135462 217332
rect 137606 217320 137612 217332
rect 137664 217320 137670 217372
rect 97954 217252 97960 217304
rect 98012 217292 98018 217304
rect 101818 217292 101824 217304
rect 98012 217264 101824 217292
rect 98012 217252 98018 217264
rect 101818 217252 101824 217264
rect 101876 217252 101882 217304
rect 181030 217252 181036 217304
rect 181088 217292 181094 217304
rect 185722 217292 185728 217304
rect 181088 217264 185728 217292
rect 181088 217252 181094 217264
rect 185722 217252 185728 217264
rect 185780 217252 185786 217304
rect 98046 217184 98052 217236
rect 98104 217224 98110 217236
rect 101726 217224 101732 217236
rect 98104 217196 101732 217224
rect 98104 217184 98110 217196
rect 101726 217184 101732 217196
rect 101784 217184 101790 217236
rect 181214 217184 181220 217236
rect 181272 217224 181278 217236
rect 185538 217224 185544 217236
rect 181272 217196 185544 217224
rect 181272 217184 181278 217196
rect 185538 217184 185544 217196
rect 185596 217184 185602 217236
rect 52690 217116 52696 217168
rect 52748 217156 52754 217168
rect 58302 217156 58308 217168
rect 52748 217128 58308 217156
rect 52748 217116 52754 217128
rect 58302 217116 58308 217128
rect 58360 217116 58366 217168
rect 92710 217116 92716 217168
rect 92768 217156 92774 217168
rect 101910 217156 101916 217168
rect 92768 217128 101916 217156
rect 92768 217116 92774 217128
rect 101910 217116 101916 217128
rect 101968 217116 101974 217168
rect 137514 217116 137520 217168
rect 137572 217156 137578 217168
rect 143678 217156 143684 217168
rect 137572 217128 143684 217156
rect 137572 217116 137578 217128
rect 143678 217116 143684 217128
rect 143736 217116 143742 217168
rect 177718 217116 177724 217168
rect 177776 217156 177782 217168
rect 185630 217156 185636 217168
rect 177776 217128 185636 217156
rect 177776 217116 177782 217128
rect 185630 217116 185636 217128
rect 185688 217116 185694 217168
rect 53058 217048 53064 217100
rect 53116 217088 53122 217100
rect 58210 217088 58216 217100
rect 53116 217060 58216 217088
rect 53116 217048 53122 217060
rect 58210 217048 58216 217060
rect 58268 217048 58274 217100
rect 93906 217048 93912 217100
rect 93964 217088 93970 217100
rect 102002 217088 102008 217100
rect 93964 217060 102008 217088
rect 93964 217048 93970 217060
rect 102002 217048 102008 217060
rect 102060 217048 102066 217100
rect 137974 217048 137980 217100
rect 138032 217088 138038 217100
rect 143126 217088 143132 217100
rect 138032 217060 143132 217088
rect 138032 217048 138038 217060
rect 143126 217048 143132 217060
rect 143184 217048 143190 217100
rect 177626 217048 177632 217100
rect 177684 217088 177690 217100
rect 185906 217088 185912 217100
rect 177684 217060 185912 217088
rect 177684 217048 177690 217060
rect 185906 217048 185912 217060
rect 185964 217048 185970 217100
rect 51126 215824 51132 215876
rect 51184 215864 51190 215876
rect 56646 215864 56652 215876
rect 51184 215836 56652 215864
rect 51184 215824 51190 215836
rect 56646 215824 56652 215836
rect 56704 215824 56710 215876
rect 98138 215824 98144 215876
rect 98196 215864 98202 215876
rect 101726 215864 101732 215876
rect 98196 215836 101732 215864
rect 98196 215824 98202 215836
rect 101726 215824 101732 215836
rect 101784 215824 101790 215876
rect 135398 215824 135404 215876
rect 135456 215864 135462 215876
rect 135456 215836 139676 215864
rect 135456 215824 135462 215836
rect 52782 215756 52788 215808
rect 52840 215796 52846 215808
rect 58302 215796 58308 215808
rect 52840 215768 58308 215796
rect 52840 215756 52846 215768
rect 58302 215756 58308 215768
rect 58360 215756 58366 215808
rect 93538 215756 93544 215808
rect 93596 215796 93602 215808
rect 101818 215796 101824 215808
rect 93596 215768 101824 215796
rect 93596 215756 93602 215768
rect 101818 215756 101824 215768
rect 101876 215756 101882 215808
rect 139648 215796 139676 215836
rect 181122 215824 181128 215876
rect 181180 215864 181186 215876
rect 185722 215864 185728 215876
rect 181180 215836 185728 215864
rect 181180 215824 181186 215836
rect 185722 215824 185728 215836
rect 185780 215824 185786 215876
rect 143494 215796 143500 215808
rect 139648 215768 143500 215796
rect 143494 215756 143500 215768
rect 143552 215756 143558 215808
rect 177626 215756 177632 215808
rect 177684 215796 177690 215808
rect 185906 215796 185912 215808
rect 177684 215768 185912 215796
rect 177684 215756 177690 215768
rect 185906 215756 185912 215768
rect 185964 215756 185970 215808
rect 52874 215688 52880 215740
rect 52932 215728 52938 215740
rect 58210 215728 58216 215740
rect 52932 215700 58216 215728
rect 52932 215688 52938 215700
rect 58210 215688 58216 215700
rect 58268 215688 58274 215740
rect 92710 215688 92716 215740
rect 92768 215728 92774 215740
rect 97954 215728 97960 215740
rect 92768 215700 97960 215728
rect 92768 215688 92774 215700
rect 97954 215688 97960 215700
rect 98012 215688 98018 215740
rect 137698 215688 137704 215740
rect 137756 215728 137762 215740
rect 143126 215728 143132 215740
rect 137756 215700 143132 215728
rect 137756 215688 137762 215700
rect 143126 215688 143132 215700
rect 143184 215688 143190 215740
rect 92802 215620 92808 215672
rect 92860 215660 92866 215672
rect 98046 215660 98052 215672
rect 92860 215632 98052 215660
rect 92860 215620 92866 215632
rect 98046 215620 98052 215632
rect 98104 215620 98110 215672
rect 137606 215620 137612 215672
rect 137664 215660 137670 215672
rect 142942 215660 142948 215672
rect 137664 215632 142948 215660
rect 137664 215620 137670 215632
rect 142942 215620 142948 215632
rect 143000 215620 143006 215672
rect 177718 215620 177724 215672
rect 177776 215660 177782 215672
rect 181030 215660 181036 215672
rect 177776 215632 181036 215660
rect 177776 215620 177782 215632
rect 181030 215620 181036 215632
rect 181088 215620 181094 215672
rect 177718 215484 177724 215536
rect 177776 215524 177782 215536
rect 181214 215524 181220 215536
rect 177776 215496 181220 215524
rect 177776 215484 177782 215496
rect 181214 215484 181220 215496
rect 181272 215484 181278 215536
rect 56646 215144 56652 215196
rect 56704 215184 56710 215196
rect 58210 215184 58216 215196
rect 56704 215156 58216 215184
rect 56704 215144 56710 215156
rect 58210 215144 58216 215156
rect 58268 215144 58274 215196
rect 50390 214872 50396 214924
rect 50448 214912 50454 214924
rect 52782 214912 52788 214924
rect 50448 214884 52788 214912
rect 50448 214872 50454 214884
rect 52782 214872 52788 214884
rect 52840 214872 52846 214924
rect 134846 214872 134852 214924
rect 134904 214912 134910 214924
rect 137606 214912 137612 214924
rect 134904 214884 137612 214912
rect 134904 214872 134910 214884
rect 137606 214872 137612 214884
rect 137664 214872 137670 214924
rect 51126 214532 51132 214584
rect 51184 214572 51190 214584
rect 52690 214572 52696 214584
rect 51184 214544 52696 214572
rect 51184 214532 51190 214544
rect 52690 214532 52696 214544
rect 52748 214532 52754 214584
rect 135306 214532 135312 214584
rect 135364 214572 135370 214584
rect 136870 214572 136876 214584
rect 135364 214544 136876 214572
rect 135364 214532 135370 214544
rect 136870 214532 136876 214544
rect 136928 214532 136934 214584
rect 181214 214532 181220 214584
rect 181272 214572 181278 214584
rect 185262 214572 185268 214584
rect 181272 214544 185268 214572
rect 181272 214532 181278 214544
rect 185262 214532 185268 214544
rect 185320 214532 185326 214584
rect 51218 214464 51224 214516
rect 51276 214504 51282 214516
rect 58302 214504 58308 214516
rect 51276 214476 58308 214504
rect 51276 214464 51282 214476
rect 58302 214464 58308 214476
rect 58360 214464 58366 214516
rect 98046 214464 98052 214516
rect 98104 214504 98110 214516
rect 101818 214504 101824 214516
rect 98104 214476 101824 214504
rect 98104 214464 98110 214476
rect 101818 214464 101824 214476
rect 101876 214464 101882 214516
rect 135398 214464 135404 214516
rect 135456 214504 135462 214516
rect 143678 214504 143684 214516
rect 135456 214476 143684 214504
rect 135456 214464 135462 214476
rect 143678 214464 143684 214476
rect 143736 214464 143742 214516
rect 181030 214464 181036 214516
rect 181088 214504 181094 214516
rect 185722 214504 185728 214516
rect 181088 214476 185728 214504
rect 181088 214464 181094 214476
rect 185722 214464 185728 214476
rect 185780 214464 185786 214516
rect 51310 214396 51316 214448
rect 51368 214436 51374 214448
rect 58210 214436 58216 214448
rect 51368 214408 58216 214436
rect 51368 214396 51374 214408
rect 58210 214396 58216 214408
rect 58268 214396 58274 214448
rect 92710 214396 92716 214448
rect 92768 214436 92774 214448
rect 100990 214436 100996 214448
rect 92768 214408 100996 214436
rect 92768 214396 92774 214408
rect 100990 214396 100996 214408
rect 101048 214396 101054 214448
rect 135490 214396 135496 214448
rect 135548 214436 135554 214448
rect 142942 214436 142948 214448
rect 135548 214408 142948 214436
rect 135548 214396 135554 214408
rect 142942 214396 142948 214408
rect 143000 214396 143006 214448
rect 177626 214396 177632 214448
rect 177684 214436 177690 214448
rect 185630 214436 185636 214448
rect 177684 214408 185636 214436
rect 177684 214396 177690 214408
rect 185630 214396 185636 214408
rect 185688 214396 185694 214448
rect 92802 214328 92808 214380
rect 92860 214368 92866 214380
rect 98138 214368 98144 214380
rect 92860 214340 98144 214368
rect 92860 214328 92866 214340
rect 98138 214328 98144 214340
rect 98196 214328 98202 214380
rect 177718 214260 177724 214312
rect 177776 214300 177782 214312
rect 181122 214300 181128 214312
rect 177776 214272 181128 214300
rect 177776 214260 177782 214272
rect 181122 214260 181128 214272
rect 181180 214260 181186 214312
rect 50206 213376 50212 213428
rect 50264 213416 50270 213428
rect 52874 213416 52880 213428
rect 50264 213388 52880 213416
rect 50264 213376 50270 213388
rect 52874 213376 52880 213388
rect 52932 213376 52938 213428
rect 135398 213376 135404 213428
rect 135456 213416 135462 213428
rect 137514 213416 137520 213428
rect 135456 213388 137520 213416
rect 135456 213376 135462 213388
rect 137514 213376 137520 213388
rect 137572 213376 137578 213428
rect 50942 213240 50948 213292
rect 51000 213280 51006 213292
rect 52966 213280 52972 213292
rect 51000 213252 52972 213280
rect 51000 213240 51006 213252
rect 52966 213240 52972 213252
rect 53024 213240 53030 213292
rect 97954 213172 97960 213224
rect 98012 213212 98018 213224
rect 101174 213212 101180 213224
rect 98012 213184 101180 213212
rect 98012 213172 98018 213184
rect 101174 213172 101180 213184
rect 101232 213172 101238 213224
rect 181950 213172 181956 213224
rect 182008 213212 182014 213224
rect 185170 213212 185176 213224
rect 182008 213184 185176 213212
rect 182008 213172 182014 213184
rect 185170 213172 185176 213184
rect 185228 213172 185234 213224
rect 98138 213104 98144 213156
rect 98196 213144 98202 213156
rect 101082 213144 101088 213156
rect 98196 213116 101088 213144
rect 98196 213104 98202 213116
rect 101082 213104 101088 213116
rect 101140 213104 101146 213156
rect 134662 213104 134668 213156
rect 134720 213144 134726 213156
rect 136962 213144 136968 213156
rect 134720 213116 136968 213144
rect 134720 213104 134726 213116
rect 136962 213104 136968 213116
rect 137020 213104 137026 213156
rect 181858 213104 181864 213156
rect 181916 213144 181922 213156
rect 185722 213144 185728 213156
rect 181916 213116 185728 213144
rect 181916 213104 181922 213116
rect 185722 213104 185728 213116
rect 185780 213104 185786 213156
rect 52690 213036 52696 213088
rect 52748 213076 52754 213088
rect 58302 213076 58308 213088
rect 52748 213048 58308 213076
rect 52748 213036 52754 213048
rect 58302 213036 58308 213048
rect 58360 213036 58366 213088
rect 93630 213036 93636 213088
rect 93688 213076 93694 213088
rect 100990 213076 100996 213088
rect 93688 213048 100996 213076
rect 93688 213036 93694 213048
rect 100990 213036 100996 213048
rect 101048 213036 101054 213088
rect 137606 213036 137612 213088
rect 137664 213076 137670 213088
rect 143678 213076 143684 213088
rect 137664 213048 143684 213076
rect 137664 213036 137670 213048
rect 143678 213036 143684 213048
rect 143736 213036 143742 213088
rect 177718 213036 177724 213088
rect 177776 213076 177782 213088
rect 181030 213076 181036 213088
rect 177776 213048 181036 213076
rect 177776 213036 177782 213048
rect 181030 213036 181036 213048
rect 181088 213036 181094 213088
rect 52782 212968 52788 213020
rect 52840 213008 52846 213020
rect 58210 213008 58216 213020
rect 52840 212980 58216 213008
rect 52840 212968 52846 212980
rect 58210 212968 58216 212980
rect 58268 212968 58274 213020
rect 92710 212968 92716 213020
rect 92768 213008 92774 213020
rect 98046 213008 98052 213020
rect 92768 212980 98052 213008
rect 92768 212968 92774 212980
rect 98046 212968 98052 212980
rect 98104 212968 98110 213020
rect 136870 212968 136876 213020
rect 136928 213008 136934 213020
rect 143494 213008 143500 213020
rect 136928 212980 143500 213008
rect 136928 212968 136934 212980
rect 143494 212968 143500 212980
rect 143552 212968 143558 213020
rect 177718 212492 177724 212544
rect 177776 212532 177782 212544
rect 181214 212532 181220 212544
rect 177776 212504 181220 212532
rect 177776 212492 177782 212504
rect 181214 212492 181220 212504
rect 181272 212492 181278 212544
rect 51218 212016 51224 212068
rect 51276 212056 51282 212068
rect 52690 212056 52696 212068
rect 51276 212028 52696 212056
rect 51276 212016 51282 212028
rect 52690 212016 52696 212028
rect 52748 212016 52754 212068
rect 135398 212016 135404 212068
rect 135456 212056 135462 212068
rect 137606 212056 137612 212068
rect 135456 212028 137612 212056
rect 135456 212016 135462 212028
rect 137606 212016 137612 212028
rect 137664 212016 137670 212068
rect 50758 211880 50764 211932
rect 50816 211920 50822 211932
rect 56462 211920 56468 211932
rect 50816 211892 56468 211920
rect 50816 211880 50822 211892
rect 56462 211880 56468 211892
rect 56520 211880 56526 211932
rect 134846 211880 134852 211932
rect 134904 211920 134910 211932
rect 139630 211920 139636 211932
rect 134904 211892 139636 211920
rect 134904 211880 134910 211892
rect 139630 211880 139636 211892
rect 139688 211880 139694 211932
rect 98046 211744 98052 211796
rect 98104 211784 98110 211796
rect 101082 211784 101088 211796
rect 98104 211756 101088 211784
rect 98104 211744 98110 211756
rect 101082 211744 101088 211756
rect 101140 211744 101146 211796
rect 182134 211744 182140 211796
rect 182192 211784 182198 211796
rect 185722 211784 185728 211796
rect 182192 211756 185728 211784
rect 182192 211744 182198 211756
rect 185722 211744 185728 211756
rect 185780 211744 185786 211796
rect 100990 211716 100996 211728
rect 98156 211688 100996 211716
rect 52966 211608 52972 211660
rect 53024 211648 53030 211660
rect 58210 211648 58216 211660
rect 53024 211620 58216 211648
rect 53024 211608 53030 211620
rect 58210 211608 58216 211620
rect 58268 211608 58274 211660
rect 93538 211608 93544 211660
rect 93596 211648 93602 211660
rect 98156 211648 98184 211688
rect 100990 211676 100996 211688
rect 101048 211676 101054 211728
rect 181674 211676 181680 211728
rect 181732 211716 181738 211728
rect 185906 211716 185912 211728
rect 181732 211688 185912 211716
rect 181732 211676 181738 211688
rect 185906 211676 185912 211688
rect 185964 211676 185970 211728
rect 93596 211620 98184 211648
rect 93596 211608 93602 211620
rect 136962 211608 136968 211660
rect 137020 211648 137026 211660
rect 143678 211648 143684 211660
rect 137020 211620 143684 211648
rect 137020 211608 137026 211620
rect 143678 211608 143684 211620
rect 143736 211608 143742 211660
rect 177718 211608 177724 211660
rect 177776 211648 177782 211660
rect 181858 211648 181864 211660
rect 177776 211620 181864 211648
rect 177776 211608 177782 211620
rect 181858 211608 181864 211620
rect 181916 211608 181922 211660
rect 52874 211540 52880 211592
rect 52932 211580 52938 211592
rect 58302 211580 58308 211592
rect 52932 211552 58308 211580
rect 52932 211540 52938 211552
rect 58302 211540 58308 211552
rect 58360 211540 58366 211592
rect 92802 211540 92808 211592
rect 92860 211580 92866 211592
rect 98138 211580 98144 211592
rect 92860 211552 98144 211580
rect 92860 211540 92866 211552
rect 98138 211540 98144 211552
rect 98196 211540 98202 211592
rect 92710 211472 92716 211524
rect 92768 211512 92774 211524
rect 97954 211512 97960 211524
rect 92768 211484 97960 211512
rect 92768 211472 92774 211484
rect 97954 211472 97960 211484
rect 98012 211472 98018 211524
rect 137514 211336 137520 211388
rect 137572 211376 137578 211388
rect 143678 211376 143684 211388
rect 137572 211348 143684 211376
rect 137572 211336 137578 211348
rect 143678 211336 143684 211348
rect 143736 211336 143742 211388
rect 177718 211268 177724 211320
rect 177776 211308 177782 211320
rect 181950 211308 181956 211320
rect 177776 211280 181956 211308
rect 177776 211268 177782 211280
rect 181950 211268 181956 211280
rect 182008 211268 182014 211320
rect 56462 211064 56468 211116
rect 56520 211104 56526 211116
rect 58394 211104 58400 211116
rect 56520 211076 58400 211104
rect 56520 211064 56526 211076
rect 58394 211064 58400 211076
rect 58452 211064 58458 211116
rect 177718 210996 177724 211048
rect 177776 211036 177782 211048
rect 182134 211036 182140 211048
rect 177776 211008 182140 211036
rect 177776 210996 177782 211008
rect 182134 210996 182140 211008
rect 182192 210996 182198 211048
rect 139630 210928 139636 210980
rect 139688 210968 139694 210980
rect 143586 210968 143592 210980
rect 139688 210940 143592 210968
rect 139688 210928 139694 210940
rect 143586 210928 143592 210940
rect 143644 210928 143650 210980
rect 51126 210656 51132 210708
rect 51184 210696 51190 210708
rect 56278 210696 56284 210708
rect 51184 210668 56284 210696
rect 51184 210656 51190 210668
rect 56278 210656 56284 210668
rect 56336 210656 56342 210708
rect 94090 210452 94096 210504
rect 94148 210492 94154 210504
rect 101174 210492 101180 210504
rect 94148 210464 101180 210492
rect 94148 210452 94154 210464
rect 101174 210452 101180 210464
rect 101232 210452 101238 210504
rect 178270 210452 178276 210504
rect 178328 210492 178334 210504
rect 185722 210492 185728 210504
rect 178328 210464 185728 210492
rect 178328 210452 178334 210464
rect 185722 210452 185728 210464
rect 185780 210452 185786 210504
rect 93998 210384 94004 210436
rect 94056 210424 94062 210436
rect 101082 210424 101088 210436
rect 94056 210396 101088 210424
rect 94056 210384 94062 210396
rect 101082 210384 101088 210396
rect 101140 210384 101146 210436
rect 178086 210384 178092 210436
rect 178144 210424 178150 210436
rect 185814 210424 185820 210436
rect 178144 210396 185820 210424
rect 178144 210384 178150 210396
rect 185814 210384 185820 210396
rect 185872 210384 185878 210436
rect 92618 210316 92624 210368
rect 92676 210356 92682 210368
rect 100990 210356 100996 210368
rect 92676 210328 100996 210356
rect 92676 210316 92682 210328
rect 100990 210316 100996 210328
rect 101048 210316 101054 210368
rect 135398 210316 135404 210368
rect 135456 210356 135462 210368
rect 135456 210328 139676 210356
rect 135456 210316 135462 210328
rect 52690 210248 52696 210300
rect 52748 210288 52754 210300
rect 58210 210288 58216 210300
rect 52748 210260 58216 210288
rect 52748 210248 52754 210260
rect 58210 210248 58216 210260
rect 58268 210248 58274 210300
rect 92710 210248 92716 210300
rect 92768 210288 92774 210300
rect 98046 210288 98052 210300
rect 92768 210260 98052 210288
rect 92768 210248 92774 210260
rect 98046 210248 98052 210260
rect 98104 210248 98110 210300
rect 139648 210288 139676 210328
rect 176798 210316 176804 210368
rect 176856 210356 176862 210368
rect 185998 210356 186004 210368
rect 176856 210328 186004 210356
rect 176856 210316 176862 210328
rect 185998 210316 186004 210328
rect 186056 210316 186062 210368
rect 143678 210288 143684 210300
rect 139648 210260 143684 210288
rect 143678 210248 143684 210260
rect 143736 210248 143742 210300
rect 137606 210180 137612 210232
rect 137664 210220 137670 210232
rect 142942 210220 142948 210232
rect 137664 210192 142948 210220
rect 137664 210180 137670 210192
rect 142942 210180 142948 210192
rect 143000 210180 143006 210232
rect 177718 210044 177724 210096
rect 177776 210084 177782 210096
rect 181674 210084 181680 210096
rect 177776 210056 181680 210084
rect 177776 210044 177782 210056
rect 181674 210044 181680 210056
rect 181732 210044 181738 210096
rect 56278 209908 56284 209960
rect 56336 209948 56342 209960
rect 58302 209948 58308 209960
rect 56336 209920 58308 209948
rect 56336 209908 56342 209920
rect 58302 209908 58308 209920
rect 58360 209908 58366 209960
rect 91238 209024 91244 209076
rect 91296 209064 91302 209076
rect 101082 209064 101088 209076
rect 91296 209036 101088 209064
rect 91296 209024 91302 209036
rect 101082 209024 101088 209036
rect 101140 209024 101146 209076
rect 175418 209024 175424 209076
rect 175476 209064 175482 209076
rect 185722 209064 185728 209076
rect 175476 209036 185728 209064
rect 175476 209024 175482 209036
rect 185722 209024 185728 209036
rect 185780 209024 185786 209076
rect 83050 208956 83056 209008
rect 83108 208996 83114 209008
rect 84246 208996 84252 209008
rect 83108 208968 84252 208996
rect 83108 208956 83114 208968
rect 84246 208956 84252 208968
rect 84304 208956 84310 209008
rect 90594 208956 90600 209008
rect 90652 208996 90658 209008
rect 100990 208996 100996 209008
rect 90652 208968 100996 208996
rect 90652 208956 90658 208968
rect 100990 208956 100996 208968
rect 101048 208956 101054 209008
rect 174774 208956 174780 209008
rect 174832 208996 174838 209008
rect 185814 208996 185820 209008
rect 174832 208968 185820 208996
rect 174832 208956 174838 208968
rect 185814 208956 185820 208968
rect 185872 208956 185878 209008
rect 51218 207664 51224 207716
rect 51276 207704 51282 207716
rect 56094 207704 56100 207716
rect 51276 207676 56100 207704
rect 51276 207664 51282 207676
rect 56094 207664 56100 207676
rect 56152 207664 56158 207716
rect 135398 207596 135404 207648
rect 135456 207636 135462 207648
rect 140274 207636 140280 207648
rect 135456 207608 140280 207636
rect 135456 207596 135462 207608
rect 140274 207596 140280 207608
rect 140332 207596 140338 207648
rect 50574 207460 50580 207512
rect 50632 207500 50638 207512
rect 61246 207500 61252 207512
rect 50632 207472 61252 207500
rect 50632 207460 50638 207472
rect 61246 207460 61252 207472
rect 61304 207460 61310 207512
rect 87558 207460 87564 207512
rect 87616 207500 87622 207512
rect 101634 207500 101640 207512
rect 87616 207472 101640 207500
rect 87616 207460 87622 207472
rect 101634 207460 101640 207472
rect 101692 207460 101698 207512
rect 134754 207460 134760 207512
rect 134812 207500 134818 207512
rect 145334 207500 145340 207512
rect 134812 207472 145340 207500
rect 134812 207460 134818 207472
rect 145334 207460 145340 207472
rect 145392 207460 145398 207512
rect 171186 207460 171192 207512
rect 171244 207500 171250 207512
rect 185906 207500 185912 207512
rect 171244 207472 185912 207500
rect 171244 207460 171250 207472
rect 185906 207460 185912 207472
rect 185964 207460 185970 207512
rect 174038 207392 174044 207444
rect 174096 207432 174102 207444
rect 187930 207432 187936 207444
rect 174096 207404 187936 207432
rect 174096 207392 174102 207404
rect 187930 207392 187936 207404
rect 187988 207392 187994 207444
rect 172566 206916 172572 206968
rect 172624 206956 172630 206968
rect 177534 206956 177540 206968
rect 172624 206928 177540 206956
rect 172624 206916 172630 206928
rect 177534 206916 177540 206928
rect 177592 206916 177598 206968
rect 148738 206780 148744 206832
rect 148796 206820 148802 206832
rect 149382 206820 149388 206832
rect 148796 206792 149388 206820
rect 148796 206780 148802 206792
rect 149382 206780 149388 206792
rect 149440 206780 149446 206832
rect 90410 206508 90416 206560
rect 90468 206548 90474 206560
rect 91146 206548 91152 206560
rect 90468 206520 91152 206548
rect 90468 206508 90474 206520
rect 91146 206508 91152 206520
rect 91204 206508 91210 206560
rect 63270 206236 63276 206288
rect 63328 206276 63334 206288
rect 65110 206276 65116 206288
rect 63328 206248 65116 206276
rect 63328 206236 63334 206248
rect 65110 206236 65116 206248
rect 65168 206236 65174 206288
rect 64742 206168 64748 206220
rect 64800 206208 64806 206220
rect 65202 206208 65208 206220
rect 64800 206180 65208 206208
rect 64800 206168 64806 206180
rect 65202 206168 65208 206180
rect 65260 206168 65266 206220
rect 66122 206168 66128 206220
rect 66180 206208 66186 206220
rect 66582 206208 66588 206220
rect 66180 206180 66588 206208
rect 66180 206168 66186 206180
rect 66582 206168 66588 206180
rect 66640 206168 66646 206220
rect 72102 206168 72108 206220
rect 72160 206208 72166 206220
rect 72654 206208 72660 206220
rect 72160 206180 72660 206208
rect 72160 206168 72166 206180
rect 72654 206168 72660 206180
rect 72712 206168 72718 206220
rect 73390 206168 73396 206220
rect 73448 206208 73454 206220
rect 74034 206208 74040 206220
rect 73448 206180 74040 206208
rect 73448 206168 73454 206180
rect 74034 206168 74040 206180
rect 74092 206168 74098 206220
rect 74770 206168 74776 206220
rect 74828 206208 74834 206220
rect 75506 206208 75512 206220
rect 74828 206180 75512 206208
rect 74828 206168 74834 206180
rect 75506 206168 75512 206180
rect 75564 206168 75570 206220
rect 76150 206168 76156 206220
rect 76208 206208 76214 206220
rect 76886 206208 76892 206220
rect 76208 206180 76892 206208
rect 76208 206168 76214 206180
rect 76886 206168 76892 206180
rect 76944 206168 76950 206220
rect 77530 206168 77536 206220
rect 77588 206208 77594 206220
rect 78358 206208 78364 206220
rect 77588 206180 78364 206208
rect 77588 206168 77594 206180
rect 78358 206168 78364 206180
rect 78416 206168 78422 206220
rect 85718 206168 85724 206220
rect 85776 206208 85782 206220
rect 100990 206208 100996 206220
rect 85776 206180 100996 206208
rect 85776 206168 85782 206180
rect 100990 206168 100996 206180
rect 101048 206168 101054 206220
rect 147266 206168 147272 206220
rect 147324 206208 147330 206220
rect 149290 206208 149296 206220
rect 147324 206180 149296 206208
rect 147324 206168 147330 206180
rect 149290 206168 149296 206180
rect 149348 206168 149354 206220
rect 150118 206168 150124 206220
rect 150176 206208 150182 206220
rect 150762 206208 150768 206220
rect 150176 206180 150768 206208
rect 150176 206168 150182 206180
rect 150762 206168 150768 206180
rect 150820 206168 150826 206220
rect 152970 206168 152976 206220
rect 153028 206208 153034 206220
rect 153522 206208 153528 206220
rect 153028 206180 153528 206208
rect 153028 206168 153034 206180
rect 153522 206168 153528 206180
rect 153580 206168 153586 206220
rect 156190 206168 156196 206220
rect 156248 206208 156254 206220
rect 156650 206208 156656 206220
rect 156248 206180 156656 206208
rect 156248 206168 156254 206180
rect 156650 206168 156656 206180
rect 156708 206168 156714 206220
rect 157570 206168 157576 206220
rect 157628 206208 157634 206220
rect 158030 206208 158036 206220
rect 157628 206180 158036 206208
rect 157628 206168 157634 206180
rect 158030 206168 158036 206180
rect 158088 206168 158094 206220
rect 158950 206168 158956 206220
rect 159008 206208 159014 206220
rect 159502 206208 159508 206220
rect 159008 206180 159508 206208
rect 159008 206168 159014 206180
rect 159502 206168 159508 206180
rect 159560 206168 159566 206220
rect 160330 206168 160336 206220
rect 160388 206208 160394 206220
rect 160882 206208 160888 206220
rect 160388 206180 160888 206208
rect 160388 206168 160394 206180
rect 160882 206168 160888 206180
rect 160940 206168 160946 206220
rect 169898 206168 169904 206220
rect 169956 206208 169962 206220
rect 185170 206208 185176 206220
rect 169956 206180 185176 206208
rect 169956 206168 169962 206180
rect 185170 206168 185176 206180
rect 185228 206168 185234 206220
rect 205410 204672 205416 204724
rect 205468 204712 205474 204724
rect 208354 204712 208360 204724
rect 205468 204684 208360 204712
rect 205468 204672 205474 204684
rect 208354 204672 208360 204684
rect 208412 204672 208418 204724
rect 22790 204604 22796 204656
rect 22848 204644 22854 204656
rect 26838 204644 26844 204656
rect 22848 204616 26844 204644
rect 22848 204604 22854 204616
rect 26838 204604 26844 204616
rect 26896 204604 26902 204656
rect 121414 204604 121420 204656
rect 121472 204644 121478 204656
rect 124266 204644 124272 204656
rect 121472 204616 124272 204644
rect 121472 204604 121478 204616
rect 124266 204604 124272 204616
rect 124324 204604 124330 204656
rect 23434 204536 23440 204588
rect 23492 204576 23498 204588
rect 26746 204576 26752 204588
rect 23492 204548 26752 204576
rect 23492 204536 23498 204548
rect 26746 204536 26752 204548
rect 26804 204536 26810 204588
rect 208354 204536 208360 204588
rect 208412 204576 208418 204588
rect 211114 204576 211120 204588
rect 208412 204548 211120 204576
rect 208412 204536 208418 204548
rect 211114 204536 211120 204548
rect 211172 204536 211178 204588
rect 26654 204468 26660 204520
rect 26712 204508 26718 204520
rect 27758 204508 27764 204520
rect 26712 204480 27764 204508
rect 26712 204468 26718 204480
rect 27758 204468 27764 204480
rect 27816 204468 27822 204520
rect 208538 204468 208544 204520
rect 208596 204508 208602 204520
rect 212218 204508 212224 204520
rect 208596 204480 212224 204508
rect 208596 204468 208602 204480
rect 212218 204468 212224 204480
rect 212276 204468 212282 204520
rect 24078 204400 24084 204452
rect 24136 204440 24142 204452
rect 28034 204440 28040 204452
rect 24136 204412 28040 204440
rect 24136 204400 24142 204412
rect 28034 204400 28040 204412
rect 28092 204400 28098 204452
rect 98966 204400 98972 204452
rect 99024 204440 99030 204452
rect 104762 204440 104768 204452
rect 99024 204412 104768 204440
rect 99024 204400 99030 204412
rect 104762 204400 104768 204412
rect 104820 204400 104826 204452
rect 120218 204400 120224 204452
rect 120276 204440 120282 204452
rect 121506 204440 121512 204452
rect 120276 204412 121512 204440
rect 120276 204400 120282 204412
rect 121506 204400 121512 204412
rect 121564 204400 121570 204452
rect 208262 204400 208268 204452
rect 208320 204440 208326 204452
rect 210562 204440 210568 204452
rect 208320 204412 210568 204440
rect 208320 204400 208326 204412
rect 210562 204400 210568 204412
rect 210620 204400 210626 204452
rect 22146 204332 22152 204384
rect 22204 204372 22210 204384
rect 26654 204372 26660 204384
rect 22204 204344 26660 204372
rect 22204 204332 22210 204344
rect 26654 204332 26660 204344
rect 26712 204332 26718 204384
rect 24722 204264 24728 204316
rect 24780 204304 24786 204316
rect 28126 204304 28132 204316
rect 24780 204276 28132 204304
rect 24780 204264 24786 204276
rect 28126 204264 28132 204276
rect 28184 204264 28190 204316
rect 99426 204264 99432 204316
rect 99484 204304 99490 204316
rect 107522 204304 107528 204316
rect 99484 204276 107528 204304
rect 99484 204264 99490 204276
rect 107522 204264 107528 204276
rect 107580 204264 107586 204316
rect 121506 204264 121512 204316
rect 121564 204304 121570 204316
rect 123162 204304 123168 204316
rect 121564 204276 123168 204304
rect 121564 204264 121570 204276
rect 123162 204264 123168 204276
rect 123220 204264 123226 204316
rect 121598 204196 121604 204248
rect 121656 204236 121662 204248
rect 123714 204236 123720 204248
rect 121656 204208 123720 204236
rect 121656 204196 121662 204208
rect 123714 204196 123720 204208
rect 123772 204196 123778 204248
rect 208446 204196 208452 204248
rect 208504 204236 208510 204248
rect 211666 204236 211672 204248
rect 208504 204208 211672 204236
rect 208504 204196 208510 204208
rect 211666 204196 211672 204208
rect 211724 204196 211730 204248
rect 99242 204128 99248 204180
rect 99300 204168 99306 204180
rect 106970 204168 106976 204180
rect 99300 204140 106976 204168
rect 99300 204128 99306 204140
rect 106970 204128 106976 204140
rect 107028 204128 107034 204180
rect 183606 204128 183612 204180
rect 183664 204168 183670 204180
rect 191334 204168 191340 204180
rect 183664 204140 191340 204168
rect 183664 204128 183670 204140
rect 191334 204128 191340 204140
rect 191392 204128 191398 204180
rect 20214 204060 20220 204112
rect 20272 204100 20278 204112
rect 41742 204100 41748 204112
rect 20272 204072 41748 204100
rect 20272 204060 20278 204072
rect 41742 204060 41748 204072
rect 41800 204060 41806 204112
rect 99518 204060 99524 204112
rect 99576 204100 99582 204112
rect 108074 204100 108080 204112
rect 99576 204072 108080 204100
rect 99576 204060 99582 204072
rect 108074 204060 108080 204072
rect 108132 204060 108138 204112
rect 183422 204060 183428 204112
rect 183480 204100 183486 204112
rect 190782 204100 190788 204112
rect 183480 204072 190788 204100
rect 183480 204060 183486 204072
rect 190782 204060 190788 204072
rect 190840 204060 190846 204112
rect 191978 204060 191984 204112
rect 192036 204100 192042 204112
rect 214426 204100 214432 204112
rect 192036 204072 214432 204100
rect 192036 204060 192042 204072
rect 214426 204060 214432 204072
rect 214484 204060 214490 204112
rect 99150 203788 99156 203840
rect 99208 203828 99214 203840
rect 106418 203828 106424 203840
rect 99208 203800 106424 203828
rect 99208 203788 99214 203800
rect 106418 203788 106424 203800
rect 106476 203788 106482 203840
rect 124266 203788 124272 203840
rect 124324 203828 124330 203840
rect 128222 203828 128228 203840
rect 124324 203800 128228 203828
rect 124324 203788 124330 203800
rect 128222 203788 128228 203800
rect 128280 203788 128286 203840
rect 123714 203720 123720 203772
rect 123772 203760 123778 203772
rect 125462 203760 125468 203772
rect 123772 203732 125468 203760
rect 123772 203720 123778 203732
rect 125462 203720 125468 203732
rect 125520 203720 125526 203772
rect 187194 203720 187200 203772
rect 187252 203760 187258 203772
rect 191886 203760 191892 203772
rect 187252 203732 191892 203760
rect 187252 203720 187258 203732
rect 191886 203720 191892 203732
rect 191944 203720 191950 203772
rect 21502 203652 21508 203704
rect 21560 203692 21566 203704
rect 26930 203692 26936 203704
rect 21560 203664 26936 203692
rect 21560 203652 21566 203664
rect 26930 203652 26936 203664
rect 26988 203652 26994 203704
rect 36038 203652 36044 203704
rect 36096 203692 36102 203704
rect 37050 203692 37056 203704
rect 36096 203664 37056 203692
rect 36096 203652 36102 203664
rect 37050 203652 37056 203664
rect 37108 203652 37114 203704
rect 124174 203652 124180 203704
rect 124232 203692 124238 203704
rect 127118 203692 127124 203704
rect 124232 203664 127124 203692
rect 124232 203652 124238 203664
rect 127118 203652 127124 203664
rect 127176 203652 127182 203704
rect 183330 203652 183336 203704
rect 183388 203692 183394 203704
rect 190230 203692 190236 203704
rect 183388 203664 190236 203692
rect 183388 203652 183394 203664
rect 190230 203652 190236 203664
rect 190288 203652 190294 203704
rect 40914 203584 40920 203636
rect 40972 203624 40978 203636
rect 43582 203624 43588 203636
rect 40972 203596 43588 203624
rect 40972 203584 40978 203596
rect 43582 203584 43588 203596
rect 43640 203584 43646 203636
rect 45054 203584 45060 203636
rect 45112 203624 45118 203636
rect 46158 203624 46164 203636
rect 45112 203596 46164 203624
rect 45112 203584 45118 203596
rect 46158 203584 46164 203596
rect 46216 203584 46222 203636
rect 99334 203584 99340 203636
rect 99392 203624 99398 203636
rect 105866 203624 105872 203636
rect 99392 203596 105872 203624
rect 99392 203584 99398 203596
rect 105866 203584 105872 203596
rect 105924 203584 105930 203636
rect 120126 203584 120132 203636
rect 120184 203624 120190 203636
rect 122610 203624 122616 203636
rect 120184 203596 122616 203624
rect 120184 203584 120190 203596
rect 122610 203584 122616 203596
rect 122668 203584 122674 203636
rect 123990 203584 123996 203636
rect 124048 203624 124054 203636
rect 126566 203624 126572 203636
rect 124048 203596 126572 203624
rect 124048 203584 124054 203596
rect 126566 203584 126572 203596
rect 126624 203584 126630 203636
rect 127854 203584 127860 203636
rect 127912 203624 127918 203636
rect 129878 203624 129884 203636
rect 127912 203596 129884 203624
rect 127912 203584 127918 203596
rect 129878 203584 129884 203596
rect 129936 203584 129942 203636
rect 183238 203584 183244 203636
rect 183296 203624 183302 203636
rect 189126 203624 189132 203636
rect 183296 203596 189132 203624
rect 183296 203584 183302 203596
rect 189126 203584 189132 203596
rect 189184 203584 189190 203636
rect 201546 203584 201552 203636
rect 201604 203624 201610 203636
rect 202834 203624 202840 203636
rect 201604 203596 202840 203624
rect 201604 203584 201610 203596
rect 202834 203584 202840 203596
rect 202892 203584 202898 203636
rect 204306 203584 204312 203636
rect 204364 203624 204370 203636
rect 206146 203624 206152 203636
rect 204364 203596 206152 203624
rect 204364 203584 204370 203596
rect 206146 203584 206152 203596
rect 206204 203584 206210 203636
rect 39534 203516 39540 203568
rect 39592 203556 39598 203568
rect 41006 203556 41012 203568
rect 39592 203528 41012 203556
rect 39592 203516 39598 203528
rect 41006 203516 41012 203528
rect 41064 203516 41070 203568
rect 41190 203516 41196 203568
rect 41248 203556 41254 203568
rect 42938 203556 42944 203568
rect 41248 203528 42944 203556
rect 41248 203516 41254 203528
rect 42938 203516 42944 203528
rect 42996 203516 43002 203568
rect 99058 203516 99064 203568
rect 99116 203556 99122 203568
rect 105314 203556 105320 203568
rect 99116 203528 105320 203556
rect 99116 203516 99122 203528
rect 105314 203516 105320 203528
rect 105372 203516 105378 203568
rect 118562 203516 118568 203568
rect 118620 203556 118626 203568
rect 119850 203556 119856 203568
rect 118620 203528 119856 203556
rect 118620 203516 118626 203528
rect 119850 203516 119856 203528
rect 119908 203516 119914 203568
rect 120034 203516 120040 203568
rect 120092 203556 120098 203568
rect 122058 203556 122064 203568
rect 120092 203528 122064 203556
rect 120092 203516 120098 203528
rect 122058 203516 122064 203528
rect 122116 203516 122122 203568
rect 123898 203516 123904 203568
rect 123956 203556 123962 203568
rect 126014 203556 126020 203568
rect 123956 203528 126020 203556
rect 123956 203516 123962 203528
rect 126014 203516 126020 203528
rect 126072 203516 126078 203568
rect 128038 203516 128044 203568
rect 128096 203556 128102 203568
rect 130430 203556 130436 203568
rect 128096 203528 130436 203556
rect 128096 203516 128102 203528
rect 130430 203516 130436 203528
rect 130488 203516 130494 203568
rect 183146 203516 183152 203568
rect 183204 203556 183210 203568
rect 188574 203556 188580 203568
rect 183204 203528 188580 203556
rect 183204 203516 183210 203528
rect 188574 203516 188580 203528
rect 188632 203516 188638 203568
rect 204490 203556 204496 203568
rect 202944 203528 204496 203556
rect 37326 203448 37332 203500
rect 37384 203488 37390 203500
rect 39074 203488 39080 203500
rect 37384 203460 39080 203488
rect 37384 203448 37390 203460
rect 39074 203448 39080 203460
rect 39132 203448 39138 203500
rect 41098 203448 41104 203500
rect 41156 203488 41162 203500
rect 42294 203488 42300 203500
rect 41156 203460 42300 203488
rect 41156 203448 41162 203460
rect 42294 203448 42300 203460
rect 42352 203448 42358 203500
rect 45514 203488 45520 203500
rect 43692 203460 45520 203488
rect 20858 203380 20864 203432
rect 20916 203420 20922 203432
rect 24354 203420 24360 203432
rect 20916 203392 24360 203420
rect 20916 203380 20922 203392
rect 24354 203380 24360 203392
rect 24412 203380 24418 203432
rect 25366 203380 25372 203432
rect 25424 203420 25430 203432
rect 26286 203420 26292 203432
rect 25424 203392 26292 203420
rect 25424 203380 25430 203392
rect 26286 203380 26292 203392
rect 26344 203380 26350 203432
rect 27942 203380 27948 203432
rect 28000 203420 28006 203432
rect 29138 203420 29144 203432
rect 28000 203392 29144 203420
rect 28000 203380 28006 203392
rect 29138 203380 29144 203392
rect 29196 203380 29202 203432
rect 29230 203380 29236 203432
rect 29288 203420 29294 203432
rect 30242 203420 30248 203432
rect 29288 203392 30248 203420
rect 29288 203380 29294 203392
rect 30242 203380 30248 203392
rect 30300 203380 30306 203432
rect 31254 203380 31260 203432
rect 31312 203420 31318 203432
rect 31806 203420 31812 203432
rect 31312 203392 31812 203420
rect 31312 203380 31318 203392
rect 31806 203380 31812 203392
rect 31864 203380 31870 203432
rect 37234 203380 37240 203432
rect 37292 203420 37298 203432
rect 38338 203420 38344 203432
rect 37292 203392 38344 203420
rect 37292 203380 37298 203392
rect 38338 203380 38344 203392
rect 38396 203380 38402 203432
rect 39626 203380 39632 203432
rect 39684 203420 39690 203432
rect 40362 203420 40368 203432
rect 39684 203392 40368 203420
rect 39684 203380 39690 203392
rect 40362 203380 40368 203392
rect 40420 203380 40426 203432
rect 41006 203380 41012 203432
rect 41064 203420 41070 203432
rect 41650 203420 41656 203432
rect 41064 203392 41656 203420
rect 41064 203380 41070 203392
rect 41650 203380 41656 203392
rect 41708 203380 41714 203432
rect 33370 203040 33376 203092
rect 33428 203080 33434 203092
rect 34198 203080 34204 203092
rect 33428 203052 34204 203080
rect 33428 203040 33434 203052
rect 34198 203040 34204 203052
rect 34256 203040 34262 203092
rect 34750 203040 34756 203092
rect 34808 203080 34814 203092
rect 35486 203080 35492 203092
rect 34808 203052 35492 203080
rect 34808 203040 34814 203052
rect 35486 203040 35492 203052
rect 35544 203040 35550 203092
rect 43692 203024 43720 203460
rect 45514 203448 45520 203460
rect 45572 203448 45578 203500
rect 98874 203448 98880 203500
rect 98932 203488 98938 203500
rect 104210 203488 104216 203500
rect 98932 203460 104216 203488
rect 98932 203448 98938 203460
rect 104210 203448 104216 203460
rect 104268 203448 104274 203500
rect 110282 203448 110288 203500
rect 110340 203488 110346 203500
rect 111018 203488 111024 203500
rect 110340 203460 111024 203488
rect 110340 203448 110346 203460
rect 111018 203448 111024 203460
rect 111076 203448 111082 203500
rect 116078 203448 116084 203500
rect 116136 203488 116142 203500
rect 116998 203488 117004 203500
rect 116136 203460 117004 203488
rect 116136 203448 116142 203460
rect 116998 203448 117004 203460
rect 117056 203448 117062 203500
rect 117642 203448 117648 203500
rect 117700 203488 117706 203500
rect 118746 203488 118752 203500
rect 117700 203460 118752 203488
rect 117700 203448 117706 203460
rect 118746 203448 118752 203460
rect 118804 203448 118810 203500
rect 118838 203448 118844 203500
rect 118896 203488 118902 203500
rect 120954 203488 120960 203500
rect 118896 203460 120960 203488
rect 118896 203448 118902 203460
rect 120954 203448 120960 203460
rect 121012 203448 121018 203500
rect 123806 203448 123812 203500
rect 123864 203488 123870 203500
rect 124818 203488 124824 203500
rect 123864 203460 124824 203488
rect 123864 203448 123870 203460
rect 124818 203448 124824 203460
rect 124876 203448 124882 203500
rect 127946 203448 127952 203500
rect 128004 203488 128010 203500
rect 129326 203488 129332 203500
rect 128004 203460 129332 203488
rect 128004 203448 128010 203460
rect 129326 203448 129332 203460
rect 129384 203448 129390 203500
rect 183054 203448 183060 203500
rect 183112 203488 183118 203500
rect 188114 203488 188120 203500
rect 183112 203460 188120 203488
rect 183112 203448 183118 203460
rect 188114 203448 188120 203460
rect 188172 203448 188178 203500
rect 202944 203432 202972 203528
rect 204490 203516 204496 203528
rect 204548 203516 204554 203568
rect 205502 203516 205508 203568
rect 205560 203556 205566 203568
rect 207802 203556 207808 203568
rect 205560 203528 207808 203556
rect 205560 203516 205566 203528
rect 207802 203516 207808 203528
rect 207860 203516 207866 203568
rect 207894 203516 207900 203568
rect 207952 203556 207958 203568
rect 209458 203556 209464 203568
rect 207952 203528 209464 203556
rect 207952 203516 207958 203528
rect 209458 203516 209464 203528
rect 209516 203516 209522 203568
rect 204398 203448 204404 203500
rect 204456 203488 204462 203500
rect 205594 203488 205600 203500
rect 204456 203460 205600 203488
rect 204456 203448 204462 203460
rect 205594 203448 205600 203460
rect 205652 203448 205658 203500
rect 205686 203448 205692 203500
rect 205744 203488 205750 203500
rect 207250 203488 207256 203500
rect 205744 203460 207256 203488
rect 205744 203448 205750 203460
rect 207250 203448 207256 203460
rect 207308 203448 207314 203500
rect 208078 203448 208084 203500
rect 208136 203488 208142 203500
rect 210010 203488 210016 203500
rect 208136 203460 210016 203488
rect 208136 203448 208142 203460
rect 210010 203448 210016 203460
rect 210068 203448 210074 203500
rect 43766 203380 43772 203432
rect 43824 203420 43830 203432
rect 44870 203420 44876 203432
rect 43824 203392 44876 203420
rect 43824 203380 43830 203392
rect 44870 203380 44876 203392
rect 44928 203380 44934 203432
rect 108626 203380 108632 203432
rect 108684 203420 108690 203432
rect 109270 203420 109276 203432
rect 108684 203392 109276 203420
rect 108684 203380 108690 203392
rect 109270 203380 109276 203392
rect 109328 203380 109334 203432
rect 109730 203380 109736 203432
rect 109788 203420 109794 203432
rect 110926 203420 110932 203432
rect 109788 203392 110932 203420
rect 109788 203380 109794 203392
rect 110926 203380 110932 203392
rect 110984 203380 110990 203432
rect 111478 203380 111484 203432
rect 111536 203420 111542 203432
rect 112306 203420 112312 203432
rect 111536 203392 112312 203420
rect 111536 203380 111542 203392
rect 112306 203380 112312 203392
rect 112364 203380 112370 203432
rect 115986 203380 115992 203432
rect 116044 203420 116050 203432
rect 116446 203420 116452 203432
rect 116044 203392 116452 203420
rect 116044 203380 116050 203392
rect 116446 203380 116452 203392
rect 116504 203380 116510 203432
rect 117274 203380 117280 203432
rect 117332 203420 117338 203432
rect 118194 203420 118200 203432
rect 117332 203392 118200 203420
rect 117332 203380 117338 203392
rect 118194 203380 118200 203392
rect 118252 203380 118258 203432
rect 118654 203380 118660 203432
rect 118712 203420 118718 203432
rect 119298 203420 119304 203432
rect 118712 203392 119304 203420
rect 118712 203380 118718 203392
rect 119298 203380 119304 203392
rect 119356 203380 119362 203432
rect 120402 203420 120408 203432
rect 119408 203392 120408 203420
rect 118746 203312 118752 203364
rect 118804 203352 118810 203364
rect 119408 203352 119436 203392
rect 120402 203380 120408 203392
rect 120460 203380 120466 203432
rect 124358 203380 124364 203432
rect 124416 203420 124422 203432
rect 127670 203420 127676 203432
rect 124416 203392 127676 203420
rect 124416 203380 124422 203392
rect 127670 203380 127676 203392
rect 127728 203380 127734 203432
rect 128130 203380 128136 203432
rect 128188 203420 128194 203432
rect 128774 203420 128780 203432
rect 128188 203392 128780 203420
rect 128188 203380 128194 203392
rect 128774 203380 128780 203392
rect 128832 203380 128838 203432
rect 183514 203380 183520 203432
rect 183572 203420 183578 203432
rect 189678 203420 189684 203432
rect 183572 203392 189684 203420
rect 183572 203380 183578 203392
rect 189678 203380 189684 203392
rect 189736 203380 189742 203432
rect 192438 203380 192444 203432
rect 192496 203420 192502 203432
rect 193358 203420 193364 203432
rect 192496 203392 193364 203420
rect 192496 203380 192502 203392
rect 193358 203380 193364 203392
rect 193416 203380 193422 203432
rect 193542 203380 193548 203432
rect 193600 203420 193606 203432
rect 194646 203420 194652 203432
rect 193600 203392 194652 203420
rect 193600 203380 193606 203392
rect 194646 203380 194652 203392
rect 194704 203380 194710 203432
rect 201454 203380 201460 203432
rect 201512 203420 201518 203432
rect 202282 203420 202288 203432
rect 201512 203392 202288 203420
rect 201512 203380 201518 203392
rect 202282 203380 202288 203392
rect 202340 203380 202346 203432
rect 202926 203380 202932 203432
rect 202984 203380 202990 203432
rect 203018 203380 203024 203432
rect 203076 203420 203082 203432
rect 203938 203420 203944 203432
rect 203076 203392 203944 203420
rect 203076 203380 203082 203392
rect 203938 203380 203944 203392
rect 203996 203380 204002 203432
rect 204214 203380 204220 203432
rect 204272 203420 204278 203432
rect 205042 203420 205048 203432
rect 204272 203392 205048 203420
rect 204272 203380 204278 203392
rect 205042 203380 205048 203392
rect 205100 203380 205106 203432
rect 205410 203380 205416 203432
rect 205468 203420 205474 203432
rect 205468 203392 205640 203420
rect 205468 203380 205474 203392
rect 205612 203364 205640 203392
rect 205778 203380 205784 203432
rect 205836 203420 205842 203432
rect 206698 203420 206704 203432
rect 205836 203392 206704 203420
rect 205836 203380 205842 203392
rect 206698 203380 206704 203392
rect 206756 203380 206762 203432
rect 207986 203380 207992 203432
rect 208044 203420 208050 203432
rect 208906 203420 208912 203432
rect 208044 203392 208912 203420
rect 208044 203380 208050 203392
rect 208906 203380 208912 203392
rect 208964 203380 208970 203432
rect 118804 203324 119436 203352
rect 118804 203312 118810 203324
rect 205594 203312 205600 203364
rect 205652 203312 205658 203364
rect 199154 203040 199160 203092
rect 199212 203080 199218 203092
rect 199798 203080 199804 203092
rect 199212 203052 199804 203080
rect 199212 203040 199218 203052
rect 199798 203040 199804 203052
rect 199856 203040 199862 203092
rect 212862 203040 212868 203092
rect 212920 203080 212926 203092
rect 213598 203080 213604 203092
rect 212920 203052 213604 203080
rect 212920 203040 212926 203052
rect 213598 203040 213604 203052
rect 213656 203040 213662 203092
rect 43674 202972 43680 203024
rect 43732 202972 43738 203024
rect 30978 202836 30984 202888
rect 31036 202876 31042 202888
rect 31898 202876 31904 202888
rect 31036 202848 31904 202876
rect 31036 202836 31042 202848
rect 31898 202836 31904 202848
rect 31956 202836 31962 202888
rect 197590 199504 197596 199556
rect 197648 199544 197654 199556
rect 198142 199544 198148 199556
rect 197648 199516 198148 199544
rect 197648 199504 197654 199516
rect 198142 199504 198148 199516
rect 198200 199504 198206 199556
rect 122886 196444 122892 196496
rect 122944 196484 122950 196496
rect 123990 196484 123996 196496
rect 122944 196456 123996 196484
rect 122944 196444 122950 196456
rect 123990 196444 123996 196456
rect 124048 196444 124054 196496
rect 194830 196444 194836 196496
rect 194888 196484 194894 196496
rect 196026 196484 196032 196496
rect 194888 196456 196032 196484
rect 194888 196444 194894 196456
rect 196026 196444 196032 196456
rect 196084 196444 196090 196496
rect 26746 196376 26752 196428
rect 26804 196416 26810 196428
rect 27390 196416 27396 196428
rect 26804 196388 27396 196416
rect 26804 196376 26810 196388
rect 27390 196376 27396 196388
rect 27448 196376 27454 196428
rect 30426 196376 30432 196428
rect 30484 196416 30490 196428
rect 31254 196416 31260 196428
rect 30484 196388 31260 196416
rect 30484 196376 30490 196388
rect 31254 196376 31260 196388
rect 31312 196376 31318 196428
rect 31714 196376 31720 196428
rect 31772 196416 31778 196428
rect 32818 196416 32824 196428
rect 31772 196388 32824 196416
rect 31772 196376 31778 196388
rect 32818 196376 32824 196388
rect 32876 196376 32882 196428
rect 39258 196376 39264 196428
rect 39316 196416 39322 196428
rect 41098 196416 41104 196428
rect 39316 196388 41104 196416
rect 39316 196376 39322 196388
rect 41098 196376 41104 196388
rect 41156 196376 41162 196428
rect 115250 196376 115256 196428
rect 115308 196416 115314 196428
rect 115894 196416 115900 196428
rect 115308 196388 115900 196416
rect 115308 196376 115314 196388
rect 115894 196376 115900 196388
rect 115952 196376 115958 196428
rect 119666 196376 119672 196428
rect 119724 196416 119730 196428
rect 120034 196416 120040 196428
rect 119724 196388 120040 196416
rect 119724 196376 119730 196388
rect 120034 196376 120040 196388
rect 120092 196376 120098 196428
rect 123622 196376 123628 196428
rect 123680 196416 123686 196428
rect 124358 196416 124364 196428
rect 123680 196388 124364 196416
rect 123680 196376 123686 196388
rect 124358 196376 124364 196388
rect 124416 196376 124422 196428
rect 125646 196376 125652 196428
rect 125704 196416 125710 196428
rect 128038 196416 128044 196428
rect 125704 196388 128044 196416
rect 125704 196376 125710 196388
rect 128038 196376 128044 196388
rect 128096 196376 128102 196428
rect 194738 196376 194744 196428
rect 194796 196416 194802 196428
rect 195658 196416 195664 196428
rect 194796 196388 195664 196416
rect 194796 196376 194802 196388
rect 195658 196376 195664 196388
rect 195716 196376 195722 196428
rect 203662 196376 203668 196428
rect 203720 196416 203726 196428
rect 204398 196416 204404 196428
rect 203720 196388 204404 196416
rect 203720 196376 203726 196388
rect 204398 196376 204404 196388
rect 204456 196376 204462 196428
rect 24354 196308 24360 196360
rect 24412 196348 24418 196360
rect 26102 196348 26108 196360
rect 24412 196320 26108 196348
rect 24412 196308 24418 196320
rect 26102 196308 26108 196320
rect 26160 196308 26166 196360
rect 26562 196308 26568 196360
rect 26620 196348 26626 196360
rect 26930 196348 26936 196360
rect 26620 196320 26936 196348
rect 26620 196308 26626 196320
rect 26930 196308 26936 196320
rect 26988 196308 26994 196360
rect 27758 196308 27764 196360
rect 27816 196348 27822 196360
rect 29690 196348 29696 196360
rect 27816 196320 29696 196348
rect 27816 196308 27822 196320
rect 29690 196308 29696 196320
rect 29748 196308 29754 196360
rect 30518 196308 30524 196360
rect 30576 196348 30582 196360
rect 31622 196348 31628 196360
rect 30576 196320 31628 196348
rect 30576 196308 30582 196320
rect 31622 196308 31628 196320
rect 31680 196308 31686 196360
rect 31990 196308 31996 196360
rect 32048 196348 32054 196360
rect 32910 196348 32916 196360
rect 32048 196320 32916 196348
rect 32048 196308 32054 196320
rect 32910 196308 32916 196320
rect 32968 196308 32974 196360
rect 33370 196308 33376 196360
rect 33428 196348 33434 196360
rect 34474 196348 34480 196360
rect 33428 196320 34480 196348
rect 33428 196308 33434 196320
rect 34474 196308 34480 196320
rect 34532 196308 34538 196360
rect 34750 196308 34756 196360
rect 34808 196348 34814 196360
rect 35302 196348 35308 196360
rect 34808 196320 35308 196348
rect 34808 196308 34814 196320
rect 35302 196308 35308 196320
rect 35360 196308 35366 196360
rect 36866 196308 36872 196360
rect 36924 196348 36930 196360
rect 37234 196348 37240 196360
rect 36924 196320 37240 196348
rect 36924 196308 36930 196320
rect 37234 196308 37240 196320
rect 37292 196308 37298 196360
rect 37694 196308 37700 196360
rect 37752 196348 37758 196360
rect 39350 196348 39356 196360
rect 37752 196320 39356 196348
rect 37752 196308 37758 196320
rect 39350 196308 39356 196320
rect 39408 196308 39414 196360
rect 40086 196308 40092 196360
rect 40144 196348 40150 196360
rect 40914 196348 40920 196360
rect 40144 196320 40920 196348
rect 40144 196308 40150 196320
rect 40914 196308 40920 196320
rect 40972 196308 40978 196360
rect 41650 196308 41656 196360
rect 41708 196348 41714 196360
rect 45054 196348 45060 196360
rect 41708 196320 45060 196348
rect 41708 196308 41714 196320
rect 45054 196308 45060 196320
rect 45112 196308 45118 196360
rect 56094 196308 56100 196360
rect 56152 196348 56158 196360
rect 57566 196348 57572 196360
rect 56152 196320 57572 196348
rect 56152 196308 56158 196320
rect 57566 196308 57572 196320
rect 57624 196308 57630 196360
rect 67778 196308 67784 196360
rect 67836 196348 67842 196360
rect 68606 196348 68612 196360
rect 67836 196320 68612 196348
rect 67836 196308 67842 196320
rect 68606 196308 68612 196320
rect 68664 196308 68670 196360
rect 80842 196308 80848 196360
rect 80900 196348 80906 196360
rect 81670 196348 81676 196360
rect 80900 196320 81676 196348
rect 80900 196308 80906 196320
rect 81670 196308 81676 196320
rect 81728 196308 81734 196360
rect 81946 196308 81952 196360
rect 82004 196348 82010 196360
rect 83050 196348 83056 196360
rect 82004 196320 83056 196348
rect 82004 196308 82010 196320
rect 83050 196308 83056 196320
rect 83108 196308 83114 196360
rect 89766 196308 89772 196360
rect 89824 196348 89830 196360
rect 90594 196348 90600 196360
rect 89824 196320 90600 196348
rect 89824 196308 89830 196320
rect 90594 196308 90600 196320
rect 90652 196308 90658 196360
rect 93078 196308 93084 196360
rect 93136 196348 93142 196360
rect 93998 196348 94004 196360
rect 93136 196320 94004 196348
rect 93136 196308 93142 196320
rect 93998 196308 94004 196320
rect 94056 196308 94062 196360
rect 109362 196308 109368 196360
rect 109420 196348 109426 196360
rect 110282 196348 110288 196360
rect 109420 196320 110288 196348
rect 109420 196308 109426 196320
rect 110282 196308 110288 196320
rect 110340 196308 110346 196360
rect 114882 196308 114888 196360
rect 114940 196348 114946 196360
rect 115342 196348 115348 196360
rect 114940 196320 115348 196348
rect 114940 196308 114946 196320
rect 115342 196308 115348 196320
rect 115400 196308 115406 196360
rect 116814 196308 116820 196360
rect 116872 196348 116878 196360
rect 117274 196348 117280 196360
rect 116872 196320 117280 196348
rect 116872 196308 116878 196320
rect 117274 196308 117280 196320
rect 117332 196308 117338 196360
rect 119298 196308 119304 196360
rect 119356 196348 119362 196360
rect 120218 196348 120224 196360
rect 119356 196320 120224 196348
rect 119356 196308 119362 196320
rect 120218 196308 120224 196320
rect 120276 196308 120282 196360
rect 120862 196308 120868 196360
rect 120920 196348 120926 196360
rect 121598 196348 121604 196360
rect 120920 196320 121604 196348
rect 120920 196308 120926 196320
rect 121598 196308 121604 196320
rect 121656 196308 121662 196360
rect 123254 196308 123260 196360
rect 123312 196348 123318 196360
rect 124174 196348 124180 196360
rect 123312 196320 124180 196348
rect 123312 196308 123318 196320
rect 124174 196308 124180 196320
rect 124232 196308 124238 196360
rect 125278 196308 125284 196360
rect 125336 196348 125342 196360
rect 127854 196348 127860 196360
rect 125336 196320 127860 196348
rect 125336 196308 125342 196320
rect 127854 196308 127860 196320
rect 127912 196308 127918 196360
rect 140274 196308 140280 196360
rect 140332 196348 140338 196360
rect 141562 196348 141568 196360
rect 140332 196320 141568 196348
rect 140332 196308 140338 196320
rect 141562 196308 141568 196320
rect 141620 196308 141626 196360
rect 163734 196308 163740 196360
rect 163792 196348 163798 196360
rect 164470 196348 164476 196360
rect 163792 196320 164476 196348
rect 163792 196308 163798 196320
rect 164470 196308 164476 196320
rect 164528 196308 164534 196360
rect 164838 196308 164844 196360
rect 164896 196348 164902 196360
rect 165850 196348 165856 196360
rect 164896 196320 165856 196348
rect 164896 196308 164902 196320
rect 165850 196308 165856 196320
rect 165908 196308 165914 196360
rect 173762 196308 173768 196360
rect 173820 196348 173826 196360
rect 174774 196348 174780 196360
rect 173820 196320 174780 196348
rect 173820 196308 173826 196320
rect 174774 196308 174780 196320
rect 174832 196308 174838 196360
rect 175970 196308 175976 196360
rect 176028 196348 176034 196360
rect 176798 196348 176804 196360
rect 176028 196320 176804 196348
rect 176028 196308 176034 196320
rect 176798 196308 176804 196320
rect 176856 196308 176862 196360
rect 177074 196308 177080 196360
rect 177132 196348 177138 196360
rect 178178 196348 178184 196360
rect 177132 196320 178184 196348
rect 177132 196308 177138 196320
rect 178178 196308 178184 196320
rect 178236 196308 178242 196360
rect 194554 196308 194560 196360
rect 194612 196348 194618 196360
rect 195290 196348 195296 196360
rect 194612 196320 195296 196348
rect 194612 196308 194618 196320
rect 195290 196308 195296 196320
rect 195348 196308 195354 196360
rect 196394 196308 196400 196360
rect 196452 196348 196458 196360
rect 197222 196348 197228 196360
rect 196452 196320 197228 196348
rect 196452 196308 196458 196320
rect 197222 196308 197228 196320
rect 197280 196308 197286 196360
rect 197590 196308 197596 196360
rect 197648 196348 197654 196360
rect 198418 196348 198424 196360
rect 197648 196320 198424 196348
rect 197648 196308 197654 196320
rect 198418 196308 198424 196320
rect 198476 196308 198482 196360
rect 199154 196308 199160 196360
rect 199212 196348 199218 196360
rect 199614 196348 199620 196360
rect 199212 196320 199620 196348
rect 199212 196308 199218 196320
rect 199614 196308 199620 196320
rect 199672 196308 199678 196360
rect 202466 196308 202472 196360
rect 202524 196348 202530 196360
rect 203018 196348 203024 196360
rect 202524 196320 203024 196348
rect 202524 196308 202530 196320
rect 203018 196308 203024 196320
rect 203076 196308 203082 196360
rect 203294 196308 203300 196360
rect 203352 196348 203358 196360
rect 204214 196348 204220 196360
rect 203352 196320 204220 196348
rect 203352 196308 203358 196320
rect 204214 196308 204220 196320
rect 204272 196308 204278 196360
rect 204858 196308 204864 196360
rect 204916 196348 204922 196360
rect 205686 196348 205692 196360
rect 204916 196320 205692 196348
rect 204916 196308 204922 196320
rect 205686 196308 205692 196320
rect 205744 196308 205750 196360
rect 206882 196308 206888 196360
rect 206940 196348 206946 196360
rect 208078 196348 208084 196360
rect 206940 196320 208084 196348
rect 206940 196308 206946 196320
rect 208078 196308 208084 196320
rect 208136 196308 208142 196360
rect 27666 196240 27672 196292
rect 27724 196280 27730 196292
rect 30058 196280 30064 196292
rect 27724 196252 30064 196280
rect 27724 196240 27730 196252
rect 30058 196240 30064 196252
rect 30116 196240 30122 196292
rect 165942 196240 165948 196292
rect 166000 196280 166006 196292
rect 167230 196280 167236 196292
rect 166000 196252 167236 196280
rect 166000 196240 166006 196252
rect 167230 196240 167236 196252
rect 167288 196240 167294 196292
rect 122426 196172 122432 196224
rect 122484 196212 122490 196224
rect 123898 196212 123904 196224
rect 122484 196184 123904 196212
rect 122484 196172 122490 196184
rect 123898 196172 123904 196184
rect 123956 196172 123962 196224
rect 29046 196104 29052 196156
rect 29104 196144 29110 196156
rect 30886 196144 30892 196156
rect 29104 196116 30892 196144
rect 29104 196104 29110 196116
rect 30886 196104 30892 196116
rect 30944 196104 30950 196156
rect 51218 196104 51224 196156
rect 51276 196144 51282 196156
rect 59774 196144 59780 196156
rect 51276 196116 59780 196144
rect 51276 196104 51282 196116
rect 59774 196104 59780 196116
rect 59832 196104 59838 196156
rect 202098 196104 202104 196156
rect 202156 196144 202162 196156
rect 202834 196144 202840 196156
rect 202156 196116 202840 196144
rect 202156 196104 202162 196116
rect 202834 196104 202840 196116
rect 202892 196104 202898 196156
rect 207250 196104 207256 196156
rect 207308 196144 207314 196156
rect 208262 196144 208268 196156
rect 207308 196116 208268 196144
rect 207308 196104 207314 196116
rect 208262 196104 208268 196116
rect 208320 196104 208326 196156
rect 38062 196036 38068 196088
rect 38120 196076 38126 196088
rect 39626 196076 39632 196088
rect 38120 196048 39632 196076
rect 38120 196036 38126 196048
rect 39626 196036 39632 196048
rect 39684 196036 39690 196088
rect 51034 196036 51040 196088
rect 51092 196076 51098 196088
rect 58670 196076 58676 196088
rect 51092 196048 58676 196076
rect 51092 196036 51098 196048
rect 58670 196036 58676 196048
rect 58728 196036 58734 196088
rect 122058 196036 122064 196088
rect 122116 196076 122122 196088
rect 123714 196076 123720 196088
rect 122116 196048 123720 196076
rect 122116 196036 122122 196048
rect 123714 196036 123720 196048
rect 123772 196036 123778 196088
rect 135214 196036 135220 196088
rect 135272 196076 135278 196088
rect 142666 196076 142672 196088
rect 135272 196048 142672 196076
rect 135272 196036 135278 196048
rect 142666 196036 142672 196048
rect 142724 196036 142730 196088
rect 38890 195968 38896 196020
rect 38948 196008 38954 196020
rect 41006 196008 41012 196020
rect 38948 195980 41012 196008
rect 38948 195968 38954 195980
rect 41006 195968 41012 195980
rect 41064 195968 41070 196020
rect 50942 195968 50948 196020
rect 51000 196008 51006 196020
rect 60878 196008 60884 196020
rect 51000 195980 60884 196008
rect 51000 195968 51006 195980
rect 60878 195968 60884 195980
rect 60936 195968 60942 196020
rect 117642 195968 117648 196020
rect 117700 196008 117706 196020
rect 118654 196008 118660 196020
rect 117700 195980 118660 196008
rect 117700 195968 117706 195980
rect 118654 195968 118660 195980
rect 118712 195968 118718 196020
rect 121690 195968 121696 196020
rect 121748 196008 121754 196020
rect 123806 196008 123812 196020
rect 121748 195980 123812 196008
rect 121748 195968 121754 195980
rect 123806 195968 123812 195980
rect 123864 195968 123870 196020
rect 134938 195968 134944 196020
rect 134996 196008 135002 196020
rect 144874 196008 144880 196020
rect 134996 195980 144880 196008
rect 134996 195968 135002 195980
rect 144874 195968 144880 195980
rect 144932 195968 144938 196020
rect 193266 195968 193272 196020
rect 193324 196008 193330 196020
rect 194462 196008 194468 196020
rect 193324 195980 194468 196008
rect 193324 195968 193330 195980
rect 194462 195968 194468 195980
rect 194520 195968 194526 196020
rect 200810 195968 200816 196020
rect 200868 196008 200874 196020
rect 201638 196008 201644 196020
rect 200868 195980 201644 196008
rect 200868 195968 200874 195980
rect 201638 195968 201644 195980
rect 201696 195968 201702 196020
rect 39626 195900 39632 195952
rect 39684 195940 39690 195952
rect 41190 195940 41196 195952
rect 39684 195912 41196 195940
rect 39684 195900 39690 195912
rect 41190 195900 41196 195912
rect 41248 195900 41254 195952
rect 50758 195900 50764 195952
rect 50816 195940 50822 195952
rect 61982 195940 61988 195952
rect 50816 195912 61988 195940
rect 50816 195900 50822 195912
rect 61982 195900 61988 195912
rect 62040 195900 62046 195952
rect 88662 195900 88668 195952
rect 88720 195940 88726 195952
rect 102094 195940 102100 195952
rect 88720 195912 102100 195940
rect 88720 195900 88726 195912
rect 102094 195900 102100 195912
rect 102152 195900 102158 195952
rect 135122 195900 135128 195952
rect 135180 195940 135186 195952
rect 145978 195940 145984 195952
rect 135180 195912 145984 195940
rect 135180 195900 135186 195912
rect 145978 195900 145984 195912
rect 146036 195900 146042 195952
rect 172658 195900 172664 195952
rect 172716 195940 172722 195952
rect 186090 195940 186096 195952
rect 172716 195912 186096 195940
rect 172716 195900 172722 195912
rect 186090 195900 186096 195912
rect 186148 195900 186154 195952
rect 204490 195900 204496 195952
rect 204548 195940 204554 195952
rect 205778 195940 205784 195952
rect 204548 195912 205784 195940
rect 204548 195900 204554 195912
rect 205778 195900 205784 195912
rect 205836 195900 205842 195952
rect 206054 195900 206060 195952
rect 206112 195940 206118 195952
rect 207986 195940 207992 195952
rect 206112 195912 207992 195940
rect 206112 195900 206118 195912
rect 207986 195900 207992 195912
rect 208044 195900 208050 195952
rect 209274 195900 209280 195952
rect 209332 195940 209338 195952
rect 213046 195940 213052 195952
rect 209332 195912 213052 195940
rect 209332 195900 209338 195912
rect 213046 195900 213052 195912
rect 213104 195900 213110 195952
rect 50850 195832 50856 195884
rect 50908 195872 50914 195884
rect 63086 195872 63092 195884
rect 50908 195844 63092 195872
rect 50908 195832 50914 195844
rect 63086 195832 63092 195844
rect 63144 195832 63150 195884
rect 91146 195832 91152 195884
rect 91204 195872 91210 195884
rect 94182 195872 94188 195884
rect 91204 195844 94188 195872
rect 91204 195832 91210 195844
rect 94182 195832 94188 195844
rect 94240 195832 94246 195884
rect 134846 195832 134852 195884
rect 134904 195872 134910 195884
rect 147082 195872 147088 195884
rect 134904 195844 147088 195872
rect 134904 195832 134910 195844
rect 147082 195832 147088 195844
rect 147140 195832 147146 195884
rect 171554 195832 171560 195884
rect 171612 195872 171618 195884
rect 186274 195872 186280 195884
rect 171612 195844 186280 195872
rect 171612 195832 171618 195844
rect 186274 195832 186280 195844
rect 186332 195832 186338 195884
rect 208814 195832 208820 195884
rect 208872 195872 208878 195884
rect 212954 195872 212960 195884
rect 208872 195844 212960 195872
rect 208872 195832 208878 195844
rect 212954 195832 212960 195844
rect 213012 195832 213018 195884
rect 26378 195764 26384 195816
rect 26436 195804 26442 195816
rect 29230 195804 29236 195816
rect 26436 195776 29236 195804
rect 26436 195764 26442 195776
rect 29230 195764 29236 195776
rect 29288 195764 29294 195816
rect 50666 195764 50672 195816
rect 50724 195804 50730 195816
rect 64190 195804 64196 195816
rect 50724 195776 64196 195804
rect 50724 195764 50730 195776
rect 64190 195764 64196 195776
rect 64248 195764 64254 195816
rect 86454 195764 86460 195816
rect 86512 195804 86518 195816
rect 101726 195804 101732 195816
rect 86512 195776 101732 195804
rect 86512 195764 86518 195776
rect 101726 195764 101732 195776
rect 101784 195764 101790 195816
rect 124450 195764 124456 195816
rect 124508 195804 124514 195816
rect 128130 195804 128136 195816
rect 124508 195776 128136 195804
rect 124508 195764 124514 195776
rect 128130 195764 128136 195776
rect 128188 195764 128194 195816
rect 135030 195764 135036 195816
rect 135088 195804 135094 195816
rect 148186 195804 148192 195816
rect 135088 195776 148192 195804
rect 135088 195764 135094 195776
rect 148186 195764 148192 195776
rect 148244 195764 148250 195816
rect 170450 195764 170456 195816
rect 170508 195804 170514 195816
rect 185906 195804 185912 195816
rect 170508 195776 185912 195804
rect 170508 195764 170514 195776
rect 185906 195764 185912 195776
rect 185964 195764 185970 195816
rect 209642 195764 209648 195816
rect 209700 195804 209706 195816
rect 212862 195804 212868 195816
rect 209700 195776 212868 195804
rect 209700 195764 209706 195776
rect 212862 195764 212868 195776
rect 212920 195764 212926 195816
rect 38430 195696 38436 195748
rect 38488 195736 38494 195748
rect 39534 195736 39540 195748
rect 38488 195708 39540 195736
rect 38488 195696 38494 195708
rect 39534 195696 39540 195708
rect 39592 195696 39598 195748
rect 41282 195696 41288 195748
rect 41340 195736 41346 195748
rect 43674 195736 43680 195748
rect 41340 195708 43680 195736
rect 41340 195696 41346 195708
rect 43674 195696 43680 195708
rect 43732 195696 43738 195748
rect 87558 195696 87564 195748
rect 87616 195736 87622 195748
rect 101910 195736 101916 195748
rect 87616 195708 101916 195736
rect 87616 195696 87622 195708
rect 101910 195696 101916 195708
rect 101968 195696 101974 195748
rect 110650 195696 110656 195748
rect 110708 195736 110714 195748
rect 111662 195736 111668 195748
rect 110708 195708 111668 195736
rect 110708 195696 110714 195708
rect 111662 195696 111668 195708
rect 111720 195696 111726 195748
rect 118102 195696 118108 195748
rect 118160 195736 118166 195748
rect 118562 195736 118568 195748
rect 118160 195708 118568 195736
rect 118160 195696 118166 195708
rect 118562 195696 118568 195708
rect 118620 195696 118626 195748
rect 135398 195696 135404 195748
rect 135456 195736 135462 195748
rect 143770 195736 143776 195748
rect 135456 195708 143776 195736
rect 135456 195696 135462 195708
rect 143770 195696 143776 195708
rect 143828 195696 143834 195748
rect 26286 195628 26292 195680
rect 26344 195668 26350 195680
rect 28862 195668 28868 195680
rect 26344 195640 28868 195668
rect 26344 195628 26350 195640
rect 28862 195628 28868 195640
rect 28920 195628 28926 195680
rect 40454 195628 40460 195680
rect 40512 195668 40518 195680
rect 43122 195668 43128 195680
rect 40512 195640 43128 195668
rect 40512 195628 40518 195640
rect 43122 195628 43128 195640
rect 43180 195628 43186 195680
rect 33462 195560 33468 195612
rect 33520 195600 33526 195612
rect 34106 195600 34112 195612
rect 33520 195572 34112 195600
rect 33520 195560 33526 195572
rect 34106 195560 34112 195572
rect 34164 195560 34170 195612
rect 36498 195560 36504 195612
rect 36556 195600 36562 195612
rect 37418 195600 37424 195612
rect 36556 195572 37424 195600
rect 36556 195560 36562 195572
rect 37418 195560 37424 195572
rect 37476 195560 37482 195612
rect 40822 195560 40828 195612
rect 40880 195600 40886 195612
rect 43766 195600 43772 195612
rect 40880 195572 43772 195600
rect 40880 195560 40886 195572
rect 43766 195560 43772 195572
rect 43824 195560 43830 195612
rect 116446 195560 116452 195612
rect 116504 195600 116510 195612
rect 117366 195600 117372 195612
rect 116504 195572 117372 195600
rect 116504 195560 116510 195572
rect 117366 195560 117372 195572
rect 117424 195560 117430 195612
rect 124818 195560 124824 195612
rect 124876 195600 124882 195612
rect 127946 195600 127952 195612
rect 124876 195572 127952 195600
rect 124876 195560 124882 195572
rect 127946 195560 127952 195572
rect 128004 195560 128010 195612
rect 135306 195560 135312 195612
rect 135364 195600 135370 195612
rect 140458 195600 140464 195612
rect 135364 195572 140464 195600
rect 135364 195560 135370 195572
rect 140458 195560 140464 195572
rect 140516 195560 140522 195612
rect 120494 195492 120500 195544
rect 120552 195532 120558 195544
rect 121506 195532 121512 195544
rect 120552 195504 121512 195532
rect 120552 195492 120558 195504
rect 121506 195492 121512 195504
rect 121564 195492 121570 195544
rect 51126 195424 51132 195476
rect 51184 195464 51190 195476
rect 56462 195464 56468 195476
rect 51184 195436 56468 195464
rect 51184 195424 51190 195436
rect 56462 195424 56468 195436
rect 56520 195424 56526 195476
rect 112030 195424 112036 195476
rect 112088 195464 112094 195476
rect 112490 195464 112496 195476
rect 112088 195436 112496 195464
rect 112088 195424 112094 195436
rect 112490 195424 112496 195436
rect 112548 195424 112554 195476
rect 29138 195288 29144 195340
rect 29196 195328 29202 195340
rect 30426 195328 30432 195340
rect 29196 195300 30432 195328
rect 29196 195288 29202 195300
rect 30426 195288 30432 195300
rect 30484 195288 30490 195340
rect 31806 195288 31812 195340
rect 31864 195328 31870 195340
rect 32450 195328 32456 195340
rect 31864 195300 32456 195328
rect 31864 195288 31870 195300
rect 32450 195288 32456 195300
rect 32508 195288 32514 195340
rect 177534 195288 177540 195340
rect 177592 195328 177598 195340
rect 179282 195328 179288 195340
rect 177592 195300 179288 195328
rect 177592 195288 177598 195300
rect 179282 195288 179288 195300
rect 179340 195288 179346 195340
rect 206422 195288 206428 195340
rect 206480 195328 206486 195340
rect 207894 195328 207900 195340
rect 206480 195300 207900 195328
rect 206480 195288 206486 195300
rect 207894 195288 207900 195300
rect 207952 195288 207958 195340
rect 182870 193180 182876 193232
rect 182928 193220 182934 193232
rect 187194 193220 187200 193232
rect 182928 193192 187200 193220
rect 182928 193180 182934 193192
rect 187194 193180 187200 193192
rect 187252 193180 187258 193232
rect 18098 190936 18104 190988
rect 18156 190976 18162 190988
rect 22330 190976 22336 190988
rect 18156 190948 22336 190976
rect 18156 190936 18162 190948
rect 22330 190936 22336 190948
rect 22388 190936 22394 190988
rect 187930 188216 187936 188268
rect 187988 188256 187994 188268
rect 191978 188256 191984 188268
rect 187988 188228 191984 188256
rect 187988 188216 187994 188228
rect 191978 188216 191984 188228
rect 192036 188216 192042 188268
rect 99426 186856 99432 186908
rect 99484 186896 99490 186908
rect 106786 186896 106792 186908
rect 99484 186868 106792 186896
rect 99484 186856 99490 186868
rect 106786 186856 106792 186868
rect 106844 186856 106850 186908
rect 13406 185496 13412 185548
rect 13464 185536 13470 185548
rect 16074 185536 16080 185548
rect 13464 185508 16080 185536
rect 13464 185496 13470 185508
rect 16074 185496 16080 185508
rect 16132 185496 16138 185548
rect 104394 184068 104400 184120
rect 104452 184108 104458 184120
rect 106786 184108 106792 184120
rect 104452 184080 106792 184108
rect 104452 184068 104458 184080
rect 106786 184068 106792 184080
rect 106844 184068 106850 184120
rect 13314 184000 13320 184052
rect 13372 184040 13378 184052
rect 22330 184040 22336 184052
rect 13372 184012 22336 184040
rect 13372 184000 13378 184012
rect 22330 184000 22336 184012
rect 22388 184000 22394 184052
rect 99518 184000 99524 184052
rect 99576 184040 99582 184052
rect 105774 184040 105780 184052
rect 99576 184012 105780 184040
rect 99576 184000 99582 184012
rect 105774 184000 105780 184012
rect 105832 184000 105838 184052
rect 182870 184000 182876 184052
rect 182928 184040 182934 184052
rect 187930 184040 187936 184052
rect 182928 184012 187936 184040
rect 182928 184000 182934 184012
rect 187930 184000 187936 184012
rect 187988 184000 187994 184052
rect 104486 182708 104492 182760
rect 104544 182748 104550 182760
rect 107154 182748 107160 182760
rect 104544 182720 107160 182748
rect 104544 182708 104550 182720
rect 107154 182708 107160 182720
rect 107212 182708 107218 182760
rect 128498 182708 128504 182760
rect 128556 182748 128562 182760
rect 137514 182748 137520 182760
rect 128556 182720 137520 182748
rect 128556 182708 128562 182720
rect 137514 182708 137520 182720
rect 137572 182708 137578 182760
rect 98598 182640 98604 182692
rect 98656 182680 98662 182692
rect 106970 182680 106976 182692
rect 98656 182652 106976 182680
rect 98656 182640 98662 182652
rect 106970 182640 106976 182652
rect 107028 182640 107034 182692
rect 183146 182640 183152 182692
rect 183204 182680 183210 182692
rect 191150 182680 191156 182692
rect 183204 182652 191156 182680
rect 183204 182640 183210 182652
rect 191150 182640 191156 182652
rect 191208 182640 191214 182692
rect 183698 181280 183704 181332
rect 183756 181320 183762 181332
rect 191978 181320 191984 181332
rect 183756 181292 191984 181320
rect 183756 181280 183762 181292
rect 191978 181280 191984 181292
rect 192036 181280 192042 181332
rect 105130 180328 105136 180380
rect 105188 180368 105194 180380
rect 106970 180368 106976 180380
rect 105188 180340 106976 180368
rect 105188 180328 105194 180340
rect 106970 180328 106976 180340
rect 107028 180328 107034 180380
rect 98414 179852 98420 179904
rect 98472 179892 98478 179904
rect 104486 179892 104492 179904
rect 98472 179864 104492 179892
rect 98472 179852 98478 179864
rect 104486 179852 104492 179864
rect 104544 179852 104550 179904
rect 182502 179852 182508 179904
rect 182560 179892 182566 179904
rect 190690 179892 190696 179904
rect 182560 179864 190696 179892
rect 182560 179852 182566 179864
rect 190690 179852 190696 179864
rect 190748 179852 190754 179904
rect 212126 179852 212132 179904
rect 212184 179892 212190 179904
rect 222338 179892 222344 179904
rect 212184 179864 222344 179892
rect 212184 179852 212190 179864
rect 222338 179852 222344 179864
rect 222396 179852 222402 179904
rect 183698 179784 183704 179836
rect 183756 179824 183762 179836
rect 190598 179824 190604 179836
rect 183756 179796 190604 179824
rect 183756 179784 183762 179796
rect 190598 179784 190604 179796
rect 190656 179784 190662 179836
rect 99518 179512 99524 179564
rect 99576 179552 99582 179564
rect 104394 179552 104400 179564
rect 99576 179524 104400 179552
rect 99576 179512 99582 179524
rect 104394 179512 104400 179524
rect 104452 179512 104458 179564
rect 44410 178560 44416 178612
rect 44468 178600 44474 178612
rect 49286 178600 49292 178612
rect 44468 178572 49292 178600
rect 44468 178560 44474 178572
rect 49286 178560 49292 178572
rect 49344 178560 49350 178612
rect 182502 178492 182508 178544
rect 182560 178532 182566 178544
rect 191978 178532 191984 178544
rect 182560 178504 191984 178532
rect 182560 178492 182566 178504
rect 191978 178492 191984 178504
rect 192036 178492 192042 178544
rect 99518 177336 99524 177388
rect 99576 177376 99582 177388
rect 105130 177376 105136 177388
rect 99576 177348 105136 177376
rect 99576 177336 99582 177348
rect 105130 177336 105136 177348
rect 105188 177336 105194 177388
rect 16074 177132 16080 177184
rect 16132 177172 16138 177184
rect 22330 177172 22336 177184
rect 16132 177144 22336 177172
rect 16132 177132 16138 177144
rect 22330 177132 22336 177144
rect 22388 177132 22394 177184
rect 98598 177132 98604 177184
rect 98656 177172 98662 177184
rect 106786 177172 106792 177184
rect 98656 177144 106792 177172
rect 98656 177132 98662 177144
rect 106786 177132 106792 177144
rect 106844 177132 106850 177184
rect 183238 176452 183244 176504
rect 183296 176492 183302 176504
rect 191978 176492 191984 176504
rect 183296 176464 191984 176492
rect 183296 176452 183302 176464
rect 191978 176452 191984 176464
rect 192036 176452 192042 176504
rect 211574 175840 211580 175892
rect 211632 175880 211638 175892
rect 216174 175880 216180 175892
rect 211632 175852 216180 175880
rect 211632 175840 211638 175852
rect 216174 175840 216180 175852
rect 216232 175840 216238 175892
rect 98230 175772 98236 175824
rect 98288 175812 98294 175824
rect 106602 175812 106608 175824
rect 98288 175784 106608 175812
rect 98288 175772 98294 175784
rect 106602 175772 106608 175784
rect 106660 175772 106666 175824
rect 183698 175092 183704 175144
rect 183756 175132 183762 175144
rect 191518 175132 191524 175144
rect 183756 175104 191524 175132
rect 183756 175092 183762 175104
rect 191518 175092 191524 175104
rect 191576 175092 191582 175144
rect 49286 174344 49292 174396
rect 49344 174384 49350 174396
rect 52690 174384 52696 174396
rect 49344 174356 52696 174384
rect 49344 174344 49350 174356
rect 52690 174344 52696 174356
rect 52748 174344 52754 174396
rect 99518 173664 99524 173716
rect 99576 173704 99582 173716
rect 106786 173704 106792 173716
rect 99576 173676 106792 173704
rect 99576 173664 99582 173676
rect 106786 173664 106792 173676
rect 106844 173664 106850 173716
rect 183330 173052 183336 173104
rect 183388 173092 183394 173104
rect 191978 173092 191984 173104
rect 183388 173064 191984 173092
rect 183388 173052 183394 173064
rect 191978 173052 191984 173064
rect 192036 173052 192042 173104
rect 99518 171692 99524 171744
rect 99576 171732 99582 171744
rect 106786 171732 106792 171744
rect 99576 171704 106792 171732
rect 99576 171692 99582 171704
rect 106786 171692 106792 171704
rect 106844 171692 106850 171744
rect 183514 171692 183520 171744
rect 183572 171732 183578 171744
rect 191150 171732 191156 171744
rect 183572 171704 191156 171732
rect 183572 171692 183578 171704
rect 191150 171692 191156 171704
rect 191208 171692 191214 171744
rect 182686 171216 182692 171268
rect 182744 171256 182750 171268
rect 185078 171256 185084 171268
rect 182744 171228 185084 171256
rect 182744 171216 182750 171228
rect 185078 171216 185084 171228
rect 185136 171216 185142 171268
rect 99242 170264 99248 170316
rect 99300 170304 99306 170316
rect 99300 170276 99656 170304
rect 99300 170264 99306 170276
rect 99628 170236 99656 170276
rect 106786 170236 106792 170248
rect 99628 170208 106792 170236
rect 106786 170196 106792 170208
rect 106844 170196 106850 170248
rect 99518 168904 99524 168956
rect 99576 168944 99582 168956
rect 106694 168944 106700 168956
rect 99576 168916 106700 168944
rect 99576 168904 99582 168916
rect 106694 168904 106700 168916
rect 106752 168904 106758 168956
rect 182502 168904 182508 168956
rect 182560 168944 182566 168956
rect 191886 168944 191892 168956
rect 182560 168916 191892 168944
rect 182560 168904 182566 168916
rect 191886 168904 191892 168916
rect 191944 168904 191950 168956
rect 185078 168836 185084 168888
rect 185136 168876 185142 168888
rect 191978 168876 191984 168888
rect 185136 168848 191984 168876
rect 185136 168836 185142 168848
rect 191978 168836 191984 168848
rect 192036 168836 192042 168888
rect 99518 167612 99524 167664
rect 99576 167652 99582 167664
rect 106878 167652 106884 167664
rect 99576 167624 106884 167652
rect 99576 167612 99582 167624
rect 106878 167612 106884 167624
rect 106936 167612 106942 167664
rect 44410 167544 44416 167596
rect 44468 167584 44474 167596
rect 53334 167584 53340 167596
rect 44468 167556 53340 167584
rect 44468 167544 44474 167556
rect 53334 167544 53340 167556
rect 53392 167544 53398 167596
rect 99426 167544 99432 167596
rect 99484 167584 99490 167596
rect 106786 167584 106792 167596
rect 99484 167556 106792 167584
rect 99484 167544 99490 167556
rect 106786 167544 106792 167556
rect 106844 167544 106850 167596
rect 183698 167544 183704 167596
rect 183756 167584 183762 167596
rect 191334 167584 191340 167596
rect 183756 167556 191340 167584
rect 183756 167544 183762 167556
rect 191334 167544 191340 167556
rect 191392 167544 191398 167596
rect 182870 166456 182876 166508
rect 182928 166496 182934 166508
rect 187930 166496 187936 166508
rect 182928 166468 187936 166496
rect 182928 166456 182934 166468
rect 187930 166456 187936 166468
rect 187988 166456 187994 166508
rect 99518 166184 99524 166236
rect 99576 166224 99582 166236
rect 107246 166224 107252 166236
rect 99576 166196 107252 166224
rect 99576 166184 99582 166196
rect 107246 166184 107252 166196
rect 107304 166184 107310 166236
rect 183698 164960 183704 165012
rect 183756 165000 183762 165012
rect 190046 165000 190052 165012
rect 183756 164972 190052 165000
rect 183756 164960 183762 164972
rect 190046 164960 190052 164972
rect 190104 164960 190110 165012
rect 99518 164756 99524 164808
rect 99576 164796 99582 164808
rect 107154 164796 107160 164808
rect 99576 164768 107160 164796
rect 99576 164756 99582 164768
rect 107154 164756 107160 164768
rect 107212 164756 107218 164808
rect 211758 163600 211764 163652
rect 211816 163640 211822 163652
rect 217002 163640 217008 163652
rect 211816 163612 217008 163640
rect 211816 163600 211822 163612
rect 217002 163600 217008 163612
rect 217060 163600 217066 163652
rect 99518 163396 99524 163448
rect 99576 163436 99582 163448
rect 104394 163436 104400 163448
rect 99576 163408 104400 163436
rect 99576 163396 99582 163408
rect 104394 163396 104400 163408
rect 104452 163396 104458 163448
rect 128498 163396 128504 163448
rect 128556 163436 128562 163448
rect 137514 163436 137520 163448
rect 128556 163408 137520 163436
rect 128556 163396 128562 163408
rect 137514 163396 137520 163408
rect 137572 163396 137578 163448
rect 183054 163396 183060 163448
rect 183112 163436 183118 163448
rect 189954 163436 189960 163448
rect 183112 163408 189960 163436
rect 183112 163396 183118 163408
rect 189954 163396 189960 163408
rect 190012 163396 190018 163448
rect 13130 163328 13136 163380
rect 13188 163368 13194 163380
rect 22974 163368 22980 163380
rect 13188 163340 22980 163368
rect 13188 163328 13194 163340
rect 22974 163328 22980 163340
rect 23032 163328 23038 163380
rect 183790 162988 183796 163040
rect 183848 163028 183854 163040
rect 191518 163028 191524 163040
rect 183848 163000 191524 163028
rect 183848 162988 183854 163000
rect 191518 162988 191524 163000
rect 191576 162988 191582 163040
rect 187930 161968 187936 162020
rect 187988 162008 187994 162020
rect 191978 162008 191984 162020
rect 187988 161980 191984 162008
rect 187988 161968 187994 161980
rect 191978 161968 191984 161980
rect 192036 161968 192042 162020
rect 212678 157072 212684 157124
rect 212736 157112 212742 157124
rect 216910 157112 216916 157124
rect 212736 157084 216916 157112
rect 212736 157072 212742 157084
rect 216910 157072 216916 157084
rect 216968 157072 216974 157124
rect 216910 156460 216916 156512
rect 216968 156500 216974 156512
rect 218290 156500 218296 156512
rect 216968 156472 218296 156500
rect 216968 156460 216974 156472
rect 218290 156460 218296 156472
rect 218348 156460 218354 156512
rect 182778 155440 182784 155492
rect 182836 155480 182842 155492
rect 188022 155480 188028 155492
rect 182836 155452 188028 155480
rect 182836 155440 182842 155452
rect 188022 155440 188028 155452
rect 188080 155440 188086 155492
rect 104394 155032 104400 155084
rect 104452 155072 104458 155084
rect 106510 155072 106516 155084
rect 104452 155044 106516 155072
rect 104452 155032 104458 155044
rect 106510 155032 106516 155044
rect 106568 155032 106574 155084
rect 212034 153672 212040 153724
rect 212092 153712 212098 153724
rect 222246 153712 222252 153724
rect 212092 153684 222252 153712
rect 212092 153672 212098 153684
rect 222246 153672 222252 153684
rect 222304 153672 222310 153724
rect 32082 152312 32088 152364
rect 32140 152352 32146 152364
rect 32818 152352 32824 152364
rect 32140 152324 32824 152352
rect 32140 152312 32146 152324
rect 32818 152312 32824 152324
rect 32876 152312 32882 152364
rect 33370 152312 33376 152364
rect 33428 152352 33434 152364
rect 34106 152352 34112 152364
rect 33428 152324 34112 152352
rect 33428 152312 33434 152324
rect 34106 152312 34112 152324
rect 34164 152312 34170 152364
rect 36866 152312 36872 152364
rect 36924 152352 36930 152364
rect 37418 152352 37424 152364
rect 36924 152324 37424 152352
rect 36924 152312 36930 152324
rect 37418 152312 37424 152324
rect 37476 152312 37482 152364
rect 37694 152312 37700 152364
rect 37752 152352 37758 152364
rect 38798 152352 38804 152364
rect 37752 152324 38804 152352
rect 37752 152312 37758 152324
rect 38798 152312 38804 152324
rect 38856 152312 38862 152364
rect 41650 152312 41656 152364
rect 41708 152352 41714 152364
rect 43674 152352 43680 152364
rect 41708 152324 43680 152352
rect 41708 152312 41714 152324
rect 43674 152312 43680 152324
rect 43732 152312 43738 152364
rect 110926 152312 110932 152364
rect 110984 152352 110990 152364
rect 111662 152352 111668 152364
rect 110984 152324 111668 152352
rect 110984 152312 110990 152324
rect 111662 152312 111668 152324
rect 111720 152312 111726 152364
rect 113594 152312 113600 152364
rect 113652 152352 113658 152364
rect 114054 152352 114060 152364
rect 113652 152324 114060 152352
rect 113652 152312 113658 152324
rect 114054 152312 114060 152324
rect 114112 152312 114118 152364
rect 117642 152312 117648 152364
rect 117700 152352 117706 152364
rect 118838 152352 118844 152364
rect 117700 152324 118844 152352
rect 117700 152312 117706 152324
rect 118838 152312 118844 152324
rect 118896 152312 118902 152364
rect 119666 152312 119672 152364
rect 119724 152352 119730 152364
rect 121966 152352 121972 152364
rect 119724 152324 121972 152352
rect 119724 152312 119730 152324
rect 121966 152312 121972 152324
rect 122024 152312 122030 152364
rect 124082 152312 124088 152364
rect 124140 152352 124146 152364
rect 127854 152352 127860 152364
rect 124140 152324 127860 152352
rect 124140 152312 124146 152324
rect 127854 152312 127860 152324
rect 127912 152312 127918 152364
rect 197590 152312 197596 152364
rect 197648 152352 197654 152364
rect 198050 152352 198056 152364
rect 197648 152324 198056 152352
rect 197648 152312 197654 152324
rect 198050 152312 198056 152324
rect 198108 152312 198114 152364
rect 200442 152312 200448 152364
rect 200500 152352 200506 152364
rect 201178 152352 201184 152364
rect 200500 152324 201184 152352
rect 200500 152312 200506 152324
rect 201178 152312 201184 152324
rect 201236 152312 201242 152364
rect 201362 152312 201368 152364
rect 201420 152352 201426 152364
rect 201638 152352 201644 152364
rect 201420 152324 201644 152352
rect 201420 152312 201426 152324
rect 201638 152312 201644 152324
rect 201696 152312 201702 152364
rect 203662 152312 203668 152364
rect 203720 152352 203726 152364
rect 205962 152352 205968 152364
rect 203720 152324 205968 152352
rect 203720 152312 203726 152324
rect 205962 152312 205968 152324
rect 206020 152312 206026 152364
rect 35302 152244 35308 152296
rect 35360 152284 35366 152296
rect 35946 152284 35952 152296
rect 35360 152256 35952 152284
rect 35360 152244 35366 152256
rect 35946 152244 35952 152256
rect 36004 152244 36010 152296
rect 36498 152244 36504 152296
rect 36556 152284 36562 152296
rect 37326 152284 37332 152296
rect 36556 152256 37332 152284
rect 36556 152244 36562 152256
rect 37326 152244 37332 152256
rect 37384 152244 37390 152296
rect 38062 152244 38068 152296
rect 38120 152284 38126 152296
rect 38614 152284 38620 152296
rect 38120 152256 38620 152284
rect 38120 152244 38126 152256
rect 38614 152244 38620 152256
rect 38672 152244 38678 152296
rect 118470 152244 118476 152296
rect 118528 152284 118534 152296
rect 120586 152284 120592 152296
rect 118528 152256 120592 152284
rect 118528 152244 118534 152256
rect 120586 152244 120592 152256
rect 120644 152244 120650 152296
rect 124818 152244 124824 152296
rect 124876 152284 124882 152296
rect 129326 152284 129332 152296
rect 124876 152256 129332 152284
rect 124876 152244 124882 152256
rect 129326 152244 129332 152256
rect 129384 152244 129390 152296
rect 203294 152244 203300 152296
rect 203352 152284 203358 152296
rect 205870 152284 205876 152296
rect 203352 152256 205876 152284
rect 203352 152244 203358 152256
rect 205870 152244 205876 152256
rect 205928 152244 205934 152296
rect 207250 152244 207256 152296
rect 207308 152284 207314 152296
rect 210746 152284 210752 152296
rect 207308 152256 210752 152284
rect 207308 152244 207314 152256
rect 210746 152244 210752 152256
rect 210804 152244 210810 152296
rect 39626 152176 39632 152228
rect 39684 152216 39690 152228
rect 43122 152216 43128 152228
rect 39684 152188 43128 152216
rect 39684 152176 39690 152188
rect 43122 152176 43128 152188
rect 43180 152176 43186 152228
rect 118746 152176 118752 152228
rect 118804 152216 118810 152228
rect 120954 152216 120960 152228
rect 118804 152188 120960 152216
rect 118804 152176 118810 152188
rect 120954 152176 120960 152188
rect 121012 152176 121018 152228
rect 196210 152176 196216 152228
rect 196268 152216 196274 152228
rect 197222 152216 197228 152228
rect 196268 152188 197228 152216
rect 196268 152176 196274 152188
rect 197222 152176 197228 152188
rect 197280 152176 197286 152228
rect 204858 152176 204864 152228
rect 204916 152216 204922 152228
rect 207342 152216 207348 152228
rect 204916 152188 207348 152216
rect 204916 152176 204922 152188
rect 207342 152176 207348 152188
rect 207400 152176 207406 152228
rect 39258 152108 39264 152160
rect 39316 152148 39322 152160
rect 43030 152148 43036 152160
rect 39316 152120 43036 152148
rect 39316 152108 39322 152120
rect 43030 152108 43036 152120
rect 43088 152108 43094 152160
rect 120034 152108 120040 152160
rect 120092 152148 120098 152160
rect 123162 152148 123168 152160
rect 120092 152120 123168 152148
rect 120092 152108 120098 152120
rect 123162 152108 123168 152120
rect 123220 152108 123226 152160
rect 204490 152108 204496 152160
rect 204548 152148 204554 152160
rect 207250 152148 207256 152160
rect 204548 152120 207256 152148
rect 204548 152108 204554 152120
rect 207250 152108 207256 152120
rect 207308 152108 207314 152160
rect 41282 152040 41288 152092
rect 41340 152080 41346 152092
rect 45146 152080 45152 152092
rect 41340 152052 45152 152080
rect 41340 152040 41346 152052
rect 45146 152040 45152 152052
rect 45204 152040 45210 152092
rect 109178 152040 109184 152092
rect 109236 152080 109242 152092
rect 110098 152080 110104 152092
rect 109236 152052 110104 152080
rect 109236 152040 109242 152052
rect 110098 152040 110104 152052
rect 110156 152040 110162 152092
rect 119298 152040 119304 152092
rect 119356 152080 119362 152092
rect 121782 152080 121788 152092
rect 119356 152052 121788 152080
rect 119356 152040 119362 152052
rect 121782 152040 121788 152052
rect 121840 152040 121846 152092
rect 124450 152040 124456 152092
rect 124508 152080 124514 152092
rect 128774 152080 128780 152092
rect 124508 152052 128780 152080
rect 124508 152040 124514 152052
rect 128774 152040 128780 152052
rect 128832 152040 128838 152092
rect 205686 152040 205692 152092
rect 205744 152080 205750 152092
rect 207986 152080 207992 152092
rect 205744 152052 207992 152080
rect 205744 152040 205750 152052
rect 207986 152040 207992 152052
rect 208044 152040 208050 152092
rect 40822 151972 40828 152024
rect 40880 152012 40886 152024
rect 45054 152012 45060 152024
rect 40880 151984 45060 152012
rect 40880 151972 40886 151984
rect 45054 151972 45060 151984
rect 45112 151972 45118 152024
rect 122886 151904 122892 151956
rect 122944 151944 122950 151956
rect 123165 151947 123223 151953
rect 123165 151944 123177 151947
rect 122944 151916 123177 151944
rect 122944 151904 122950 151916
rect 123165 151913 123177 151916
rect 123211 151913 123223 151947
rect 123165 151907 123223 151913
rect 123254 151904 123260 151956
rect 123312 151944 123318 151956
rect 127210 151944 127216 151956
rect 123312 151916 127216 151944
rect 123312 151904 123318 151916
rect 127210 151904 127216 151916
rect 127268 151904 127274 151956
rect 205226 151904 205232 151956
rect 205284 151944 205290 151956
rect 207894 151944 207900 151956
rect 205284 151916 207900 151944
rect 205284 151904 205290 151916
rect 207894 151904 207900 151916
rect 207952 151904 207958 151956
rect 31806 151836 31812 151888
rect 31864 151876 31870 151888
rect 32450 151876 32456 151888
rect 31864 151848 32456 151876
rect 31864 151836 31870 151848
rect 32450 151836 32456 151848
rect 32508 151836 32514 151888
rect 112122 151836 112128 151888
rect 112180 151876 112186 151888
rect 112858 151876 112864 151888
rect 112180 151848 112864 151876
rect 112180 151836 112186 151848
rect 112858 151836 112864 151848
rect 112916 151836 112922 151888
rect 31990 151768 31996 151820
rect 32048 151808 32054 151820
rect 33278 151808 33284 151820
rect 32048 151780 33284 151808
rect 32048 151768 32054 151780
rect 33278 151768 33284 151780
rect 33336 151768 33342 151820
rect 40454 151768 40460 151820
rect 40512 151808 40518 151820
rect 44778 151808 44784 151820
rect 40512 151780 44784 151808
rect 40512 151768 40518 151780
rect 44778 151768 44784 151780
rect 44836 151768 44842 151820
rect 79186 151768 79192 151820
rect 79244 151808 79250 151820
rect 96114 151808 96120 151820
rect 79244 151780 96120 151808
rect 79244 151768 79250 151780
rect 96114 151768 96120 151780
rect 96172 151768 96178 151820
rect 120862 151768 120868 151820
rect 120920 151808 120926 151820
rect 123714 151808 123720 151820
rect 120920 151780 123720 151808
rect 120920 151768 120926 151780
rect 123714 151768 123720 151780
rect 123772 151768 123778 151820
rect 72562 151700 72568 151752
rect 72620 151740 72626 151752
rect 98874 151740 98880 151752
rect 72620 151712 98880 151740
rect 72620 151700 72626 151712
rect 98874 151700 98880 151712
rect 98932 151740 98938 151752
rect 156558 151740 156564 151752
rect 98932 151712 156564 151740
rect 98932 151700 98938 151712
rect 156558 151700 156564 151712
rect 156616 151700 156622 151752
rect 69158 151632 69164 151684
rect 69216 151672 69222 151684
rect 92526 151672 92532 151684
rect 69216 151644 92532 151672
rect 69216 151632 69222 151644
rect 92526 151632 92532 151644
rect 92584 151632 92590 151684
rect 96114 151632 96120 151684
rect 96172 151672 96178 151684
rect 163182 151672 163188 151684
rect 96172 151644 163188 151672
rect 96172 151632 96178 151644
rect 163182 151632 163188 151644
rect 163240 151632 163246 151684
rect 40086 151564 40092 151616
rect 40144 151604 40150 151616
rect 43766 151604 43772 151616
rect 40144 151576 43772 151604
rect 40144 151564 40150 151576
rect 43766 151564 43772 151576
rect 43824 151564 43830 151616
rect 123622 151564 123628 151616
rect 123680 151604 123686 151616
rect 127946 151604 127952 151616
rect 123680 151576 127952 151604
rect 123680 151564 123686 151576
rect 127946 151564 127952 151576
rect 128004 151564 128010 151616
rect 123165 151539 123223 151545
rect 123165 151505 123177 151539
rect 123211 151536 123223 151539
rect 127302 151536 127308 151548
rect 123211 151508 127308 151536
rect 123211 151505 123223 151508
rect 123165 151499 123223 151505
rect 127302 151496 127308 151508
rect 127360 151496 127366 151548
rect 24998 151428 25004 151480
rect 25056 151468 25062 151480
rect 28494 151468 28500 151480
rect 25056 151440 28500 151468
rect 25056 151428 25062 151440
rect 28494 151428 28500 151440
rect 28552 151428 28558 151480
rect 204030 151428 204036 151480
rect 204088 151468 204094 151480
rect 206054 151468 206060 151480
rect 204088 151440 206060 151468
rect 204088 151428 204094 151440
rect 206054 151428 206060 151440
rect 206112 151428 206118 151480
rect 206422 151428 206428 151480
rect 206480 151468 206486 151480
rect 210010 151468 210016 151480
rect 206480 151440 210016 151468
rect 206480 151428 206486 151440
rect 210010 151428 210016 151440
rect 210068 151428 210074 151480
rect 24906 151360 24912 151412
rect 24964 151400 24970 151412
rect 28034 151400 28040 151412
rect 24964 151372 28040 151400
rect 24964 151360 24970 151372
rect 28034 151360 28040 151372
rect 28092 151360 28098 151412
rect 121690 151360 121696 151412
rect 121748 151400 121754 151412
rect 124634 151400 124640 151412
rect 121748 151372 124640 151400
rect 121748 151360 121754 151372
rect 124634 151360 124640 151372
rect 124692 151360 124698 151412
rect 202466 151360 202472 151412
rect 202524 151400 202530 151412
rect 203018 151400 203024 151412
rect 202524 151372 203024 151400
rect 202524 151360 202530 151372
rect 203018 151360 203024 151372
rect 203076 151360 203082 151412
rect 206882 151360 206888 151412
rect 206940 151400 206946 151412
rect 210102 151400 210108 151412
rect 206940 151372 210108 151400
rect 206940 151360 206946 151372
rect 210102 151360 210108 151372
rect 210160 151360 210166 151412
rect 26378 151292 26384 151344
rect 26436 151332 26442 151344
rect 29230 151332 29236 151344
rect 26436 151304 29236 151332
rect 26436 151292 26442 151304
rect 29230 151292 29236 151304
rect 29288 151292 29294 151344
rect 122426 151292 122432 151344
rect 122484 151332 122490 151344
rect 125186 151332 125192 151344
rect 122484 151304 125192 151332
rect 122484 151292 122490 151304
rect 125186 151292 125192 151304
rect 125244 151292 125250 151344
rect 125646 151292 125652 151344
rect 125704 151332 125710 151344
rect 131350 151332 131356 151344
rect 125704 151304 131356 151332
rect 125704 151292 125710 151304
rect 131350 151292 131356 151304
rect 131408 151292 131414 151344
rect 207618 151292 207624 151344
rect 207676 151332 207682 151344
rect 210654 151332 210660 151344
rect 207676 151304 210660 151332
rect 207676 151292 207682 151304
rect 210654 151292 210660 151304
rect 210712 151292 210718 151344
rect 25734 151224 25740 151276
rect 25792 151264 25798 151276
rect 27666 151264 27672 151276
rect 25792 151236 27672 151264
rect 25792 151224 25798 151236
rect 27666 151224 27672 151236
rect 27724 151224 27730 151276
rect 116446 151224 116452 151276
rect 116504 151264 116510 151276
rect 117182 151264 117188 151276
rect 116504 151236 117188 151264
rect 116504 151224 116510 151236
rect 117182 151224 117188 151236
rect 117240 151224 117246 151276
rect 118102 151224 118108 151276
rect 118160 151264 118166 151276
rect 120310 151264 120316 151276
rect 118160 151236 120316 151264
rect 118160 151224 118166 151236
rect 120310 151224 120316 151236
rect 120368 151224 120374 151276
rect 120494 151224 120500 151276
rect 120552 151264 120558 151276
rect 123070 151264 123076 151276
rect 120552 151236 123076 151264
rect 120552 151224 120558 151236
rect 123070 151224 123076 151236
rect 123128 151224 123134 151276
rect 200810 151224 200816 151276
rect 200868 151264 200874 151276
rect 201546 151264 201552 151276
rect 200868 151236 201552 151264
rect 200868 151224 200874 151236
rect 201546 151224 201552 151236
rect 201604 151224 201610 151276
rect 208814 151224 208820 151276
rect 208872 151264 208878 151276
rect 212862 151264 212868 151276
rect 208872 151236 212868 151264
rect 208872 151224 208878 151236
rect 212862 151224 212868 151236
rect 212920 151224 212926 151276
rect 26286 151156 26292 151208
rect 26344 151196 26350 151208
rect 28862 151196 28868 151208
rect 26344 151168 28868 151196
rect 26344 151156 26350 151168
rect 28862 151156 28868 151168
rect 28920 151156 28926 151208
rect 29138 151156 29144 151208
rect 29196 151196 29202 151208
rect 30426 151196 30432 151208
rect 29196 151168 30432 151196
rect 29196 151156 29202 151168
rect 30426 151156 30432 151168
rect 30484 151156 30490 151208
rect 208078 151156 208084 151208
rect 208136 151196 208142 151208
rect 210838 151196 210844 151208
rect 208136 151168 210844 151196
rect 208136 151156 208142 151168
rect 210838 151156 210844 151168
rect 210896 151156 210902 151208
rect 25918 151088 25924 151140
rect 25976 151128 25982 151140
rect 27298 151128 27304 151140
rect 25976 151100 27304 151128
rect 25976 151088 25982 151100
rect 27298 151088 27304 151100
rect 27356 151088 27362 151140
rect 29046 151088 29052 151140
rect 29104 151128 29110 151140
rect 30886 151128 30892 151140
rect 29104 151100 30892 151128
rect 29104 151088 29110 151100
rect 30886 151088 30892 151100
rect 30944 151088 30950 151140
rect 208446 151088 208452 151140
rect 208504 151128 208510 151140
rect 210930 151128 210936 151140
rect 208504 151100 210936 151128
rect 208504 151088 208510 151100
rect 210930 151088 210936 151100
rect 210988 151088 210994 151140
rect 25826 151020 25832 151072
rect 25884 151060 25890 151072
rect 26838 151060 26844 151072
rect 25884 151032 26844 151060
rect 25884 151020 25890 151032
rect 26838 151020 26844 151032
rect 26896 151020 26902 151072
rect 27666 151020 27672 151072
rect 27724 151060 27730 151072
rect 30058 151060 30064 151072
rect 27724 151032 30064 151060
rect 27724 151020 27730 151032
rect 30058 151020 30064 151032
rect 30116 151020 30122 151072
rect 30426 151020 30432 151072
rect 30484 151060 30490 151072
rect 31622 151060 31628 151072
rect 30484 151032 31628 151060
rect 30484 151020 30490 151032
rect 31622 151020 31628 151032
rect 31680 151020 31686 151072
rect 109362 151020 109368 151072
rect 109420 151060 109426 151072
rect 110190 151060 110196 151072
rect 109420 151032 110196 151060
rect 109420 151020 109426 151032
rect 110190 151020 110196 151032
rect 110248 151020 110254 151072
rect 121230 151020 121236 151072
rect 121288 151060 121294 151072
rect 123806 151060 123812 151072
rect 121288 151032 123812 151060
rect 121288 151020 121294 151032
rect 123806 151020 123812 151032
rect 123864 151020 123870 151072
rect 125278 151020 125284 151072
rect 125336 151060 125342 151072
rect 129234 151060 129240 151072
rect 125336 151032 129240 151060
rect 125336 151020 125342 151032
rect 129234 151020 129240 151032
rect 129292 151020 129298 151072
rect 193358 151020 193364 151072
rect 193416 151060 193422 151072
rect 194462 151060 194468 151072
rect 193416 151032 194468 151060
rect 193416 151020 193422 151032
rect 194462 151020 194468 151032
rect 194520 151020 194526 151072
rect 209274 151020 209280 151072
rect 209332 151060 209338 151072
rect 214150 151060 214156 151072
rect 209332 151032 214156 151060
rect 209332 151020 209338 151032
rect 214150 151020 214156 151032
rect 214208 151020 214214 151072
rect 26010 150952 26016 151004
rect 26068 150992 26074 151004
rect 26470 150992 26476 151004
rect 26068 150964 26476 150992
rect 26068 150952 26074 150964
rect 26470 150952 26476 150964
rect 26528 150952 26534 151004
rect 27758 150952 27764 151004
rect 27816 150992 27822 151004
rect 29690 150992 29696 151004
rect 27816 150964 29696 150992
rect 27816 150952 27822 150964
rect 29690 150952 29696 150964
rect 29748 150952 29754 151004
rect 30518 150952 30524 151004
rect 30576 150992 30582 151004
rect 31254 150992 31260 151004
rect 30576 150964 31260 150992
rect 30576 150952 30582 150964
rect 31254 150952 31260 150964
rect 31312 150952 31318 151004
rect 38890 150952 38896 151004
rect 38948 150992 38954 151004
rect 41834 150992 41840 151004
rect 38948 150964 41840 150992
rect 38948 150952 38954 150964
rect 41834 150952 41840 150964
rect 41892 150952 41898 151004
rect 111294 150992 111300 151004
rect 110576 150964 111300 150992
rect 110576 150936 110604 150964
rect 111294 150952 111300 150964
rect 111352 150952 111358 151004
rect 115250 150952 115256 151004
rect 115308 150992 115314 151004
rect 115802 150992 115808 151004
rect 115308 150964 115808 150992
rect 115308 150952 115314 150964
rect 115802 150952 115808 150964
rect 115860 150952 115866 151004
rect 122058 150952 122064 151004
rect 122116 150992 122122 151004
rect 125094 150992 125100 151004
rect 122116 150964 125100 150992
rect 122116 150952 122122 150964
rect 125094 150952 125100 150964
rect 125152 150952 125158 151004
rect 193266 150952 193272 151004
rect 193324 150992 193330 151004
rect 194094 150992 194100 151004
rect 193324 150964 194100 150992
rect 193324 150952 193330 150964
rect 194094 150952 194100 150964
rect 194152 150952 194158 151004
rect 195474 150952 195480 151004
rect 195532 150992 195538 151004
rect 196026 150992 196032 151004
rect 195532 150964 196032 150992
rect 195532 150952 195538 150964
rect 196026 150952 196032 150964
rect 196084 150952 196090 151004
rect 196302 150952 196308 151004
rect 196360 150992 196366 151004
rect 196854 150992 196860 151004
rect 196360 150964 196860 150992
rect 196360 150952 196366 150964
rect 196854 150952 196860 150964
rect 196912 150952 196918 151004
rect 202098 150952 202104 151004
rect 202156 150992 202162 151004
rect 202742 150992 202748 151004
rect 202156 150964 202748 150992
rect 202156 150952 202162 150964
rect 202742 150952 202748 150964
rect 202800 150952 202806 151004
rect 206330 150952 206336 151004
rect 206388 150992 206394 151004
rect 208814 150992 208820 151004
rect 206388 150964 208820 150992
rect 206388 150952 206394 150964
rect 208814 150952 208820 150964
rect 208872 150952 208878 151004
rect 209642 150952 209648 151004
rect 209700 150992 209706 151004
rect 214242 150992 214248 151004
rect 209700 150964 214248 150992
rect 209700 150952 209706 150964
rect 214242 150952 214248 150964
rect 214300 150952 214306 151004
rect 110558 150884 110564 150936
rect 110616 150884 110622 150936
rect 196210 148300 196216 148352
rect 196268 148340 196274 148352
rect 197038 148340 197044 148352
rect 196268 148312 197044 148340
rect 196268 148300 196274 148312
rect 197038 148300 197044 148312
rect 197096 148300 197102 148352
rect 33370 147348 33376 147400
rect 33428 147388 33434 147400
rect 34198 147388 34204 147400
rect 33428 147360 34204 147388
rect 33428 147348 33434 147360
rect 34198 147348 34204 147360
rect 34256 147348 34262 147400
rect 59222 146804 59228 146856
rect 59280 146804 59286 146856
rect 59240 146776 59268 146804
rect 59406 146776 59412 146788
rect 59240 146748 59412 146776
rect 59406 146736 59412 146748
rect 59464 146736 59470 146788
rect 123070 146124 123076 146176
rect 123128 146164 123134 146176
rect 123622 146164 123628 146176
rect 123128 146136 123628 146164
rect 123128 146124 123134 146136
rect 123622 146124 123628 146136
rect 123680 146124 123686 146176
rect 127210 146124 127216 146176
rect 127268 146164 127274 146176
rect 127670 146164 127676 146176
rect 127268 146136 127676 146164
rect 127268 146124 127274 146136
rect 127670 146124 127676 146136
rect 127728 146124 127734 146176
rect 197590 146124 197596 146176
rect 197648 146164 197654 146176
rect 198142 146164 198148 146176
rect 197648 146136 198148 146164
rect 197648 146124 197654 146136
rect 198142 146124 198148 146136
rect 198200 146124 198206 146176
rect 59406 144056 59412 144068
rect 59367 144028 59412 144056
rect 59406 144016 59412 144028
rect 59464 144016 59470 144068
rect 118838 144016 118844 144068
rect 118896 144056 118902 144068
rect 119574 144056 119580 144068
rect 118896 144028 119580 144056
rect 118896 144016 118902 144028
rect 119574 144016 119580 144028
rect 119632 144016 119638 144068
rect 120954 144016 120960 144068
rect 121012 144056 121018 144068
rect 121690 144056 121696 144068
rect 121012 144028 121696 144056
rect 121012 144016 121018 144028
rect 121690 144016 121696 144028
rect 121748 144016 121754 144068
rect 123806 144016 123812 144068
rect 123864 144056 123870 144068
rect 124542 144056 124548 144068
rect 123864 144028 124548 144056
rect 123864 144016 123870 144028
rect 124542 144016 124548 144028
rect 124600 144016 124606 144068
rect 125094 144016 125100 144068
rect 125152 144056 125158 144068
rect 126014 144056 126020 144068
rect 125152 144028 126020 144056
rect 125152 144016 125158 144028
rect 126014 144016 126020 144028
rect 126072 144016 126078 144068
rect 127946 144016 127952 144068
rect 128004 144056 128010 144068
rect 128590 144056 128596 144068
rect 128004 144028 128596 144056
rect 128004 144016 128010 144028
rect 128590 144016 128596 144028
rect 128648 144016 128654 144068
rect 129326 144016 129332 144068
rect 129384 144056 129390 144068
rect 130062 144056 130068 144068
rect 129384 144028 130068 144056
rect 129384 144016 129390 144028
rect 130062 144016 130068 144028
rect 130120 144016 130126 144068
rect 183606 144016 183612 144068
rect 183664 144056 183670 144068
rect 187930 144056 187936 144068
rect 183664 144028 187936 144056
rect 183664 144016 183670 144028
rect 187930 144016 187936 144028
rect 187988 144016 187994 144068
rect 198418 144016 198424 144068
rect 198476 144056 198482 144068
rect 199062 144056 199068 144068
rect 198476 144028 199068 144056
rect 198476 144016 198482 144028
rect 199062 144016 199068 144028
rect 199120 144016 199126 144068
rect 201546 144016 201552 144068
rect 201604 144056 201610 144068
rect 202190 144056 202196 144068
rect 201604 144028 202196 144056
rect 201604 144016 201610 144028
rect 202190 144016 202196 144028
rect 202248 144016 202254 144068
rect 203018 144016 203024 144068
rect 203076 144056 203082 144068
rect 204490 144056 204496 144068
rect 203076 144028 204496 144056
rect 203076 144016 203082 144028
rect 204490 144016 204496 144028
rect 204548 144016 204554 144068
rect 207986 144016 207992 144068
rect 208044 144056 208050 144068
rect 208722 144056 208728 144068
rect 208044 144028 208728 144056
rect 208044 144016 208050 144028
rect 208722 144016 208728 144028
rect 208780 144016 208786 144068
rect 210746 144016 210752 144068
rect 210804 144056 210810 144068
rect 211390 144056 211396 144068
rect 210804 144028 211396 144056
rect 210804 144016 210810 144028
rect 211390 144016 211396 144028
rect 211448 144016 211454 144068
rect 21778 143948 21784 144000
rect 21836 143988 21842 144000
rect 26010 143988 26016 144000
rect 21836 143960 26016 143988
rect 21836 143948 21842 143960
rect 26010 143948 26016 143960
rect 26068 143948 26074 144000
rect 41834 143948 41840 144000
rect 41892 143988 41898 144000
rect 42294 143988 42300 144000
rect 41892 143960 42300 143988
rect 41892 143948 41898 143960
rect 42294 143948 42300 143960
rect 42352 143948 42358 144000
rect 123714 143948 123720 144000
rect 123772 143988 123778 144000
rect 124450 143988 124456 144000
rect 123772 143960 124456 143988
rect 123772 143948 123778 143960
rect 124450 143948 124456 143960
rect 124508 143948 124514 144000
rect 125186 143948 125192 144000
rect 125244 143988 125250 144000
rect 126566 143988 126572 144000
rect 125244 143960 126572 143988
rect 125244 143948 125250 143960
rect 126566 143948 126572 143960
rect 126624 143948 126630 144000
rect 127854 143948 127860 144000
rect 127912 143988 127918 144000
rect 128682 143988 128688 144000
rect 127912 143960 128688 143988
rect 127912 143948 127918 143960
rect 128682 143948 128688 143960
rect 128740 143948 128746 144000
rect 129234 143948 129240 144000
rect 129292 143988 129298 144000
rect 130614 143988 130620 144000
rect 129292 143960 130620 143988
rect 129292 143948 129298 143960
rect 130614 143948 130620 143960
rect 130672 143948 130678 144000
rect 183422 143948 183428 144000
rect 183480 143988 183486 144000
rect 189402 143988 189408 144000
rect 183480 143960 189408 143988
rect 183480 143948 183486 143960
rect 189402 143948 189408 143960
rect 189460 143948 189466 144000
rect 198878 143948 198884 144000
rect 198936 143988 198942 144000
rect 199246 143988 199252 144000
rect 198936 143960 199252 143988
rect 198936 143948 198942 143960
rect 199246 143948 199252 143960
rect 199304 143948 199310 144000
rect 201178 143948 201184 144000
rect 201236 143988 201242 144000
rect 201730 143988 201736 144000
rect 201236 143960 201736 143988
rect 201236 143948 201242 143960
rect 201730 143948 201736 143960
rect 201788 143948 201794 144000
rect 202742 143948 202748 144000
rect 202800 143988 202806 144000
rect 203846 143988 203852 144000
rect 202800 143960 203852 143988
rect 202800 143948 202806 143960
rect 203846 143948 203852 143960
rect 203904 143948 203910 144000
rect 207894 143948 207900 144000
rect 207952 143988 207958 144000
rect 208630 143988 208636 144000
rect 207952 143960 208636 143988
rect 207952 143948 207958 143960
rect 208630 143948 208636 143960
rect 208688 143948 208694 144000
rect 210838 143948 210844 144000
rect 210896 143988 210902 144000
rect 212310 143988 212316 144000
rect 210896 143960 212316 143988
rect 210896 143948 210902 143960
rect 212310 143948 212316 143960
rect 212368 143948 212374 144000
rect 117458 143880 117464 143932
rect 117516 143920 117522 143932
rect 119022 143920 119028 143932
rect 117516 143892 119028 143920
rect 117516 143880 117522 143892
rect 119022 143880 119028 143892
rect 119080 143880 119086 143932
rect 183514 143880 183520 143932
rect 183572 143920 183578 143932
rect 190046 143920 190052 143932
rect 183572 143892 190052 143920
rect 183572 143880 183578 143892
rect 190046 143880 190052 143892
rect 190104 143880 190110 143932
rect 202834 143880 202840 143932
rect 202892 143920 202898 143932
rect 204950 143920 204956 143932
rect 202892 143892 204956 143920
rect 202892 143880 202898 143892
rect 204950 143880 204956 143892
rect 205008 143880 205014 143932
rect 210654 143880 210660 143932
rect 210712 143920 210718 143932
rect 211758 143920 211764 143932
rect 210712 143892 211764 143920
rect 210712 143880 210718 143892
rect 211758 143880 211764 143892
rect 211816 143880 211822 143932
rect 38706 143812 38712 143864
rect 38764 143852 38770 143864
rect 41834 143852 41840 143864
rect 38764 143824 41840 143852
rect 38764 143812 38770 143824
rect 41834 143812 41840 143824
rect 41892 143812 41898 143864
rect 183330 143812 183336 143864
rect 183388 143852 183394 143864
rect 189494 143852 189500 143864
rect 183388 143824 189500 143852
rect 183388 143812 183394 143824
rect 189494 143812 189500 143824
rect 189552 143812 189558 143864
rect 201454 143812 201460 143864
rect 201512 143852 201518 143864
rect 202742 143852 202748 143864
rect 201512 143824 202748 143852
rect 201512 143812 201518 143824
rect 202742 143812 202748 143824
rect 202800 143812 202806 143864
rect 210930 143812 210936 143864
rect 210988 143852 210994 143864
rect 212954 143852 212960 143864
rect 210988 143824 212960 143852
rect 210988 143812 210994 143824
rect 212954 143812 212960 143824
rect 213012 143812 213018 143864
rect 201362 143744 201368 143796
rect 201420 143784 201426 143796
rect 203294 143784 203300 143796
rect 201420 143756 203300 143784
rect 201420 143744 201426 143756
rect 203294 143744 203300 143756
rect 203352 143744 203358 143796
rect 24446 143676 24452 143728
rect 24504 143716 24510 143728
rect 24906 143716 24912 143728
rect 24504 143688 24912 143716
rect 24504 143676 24510 143688
rect 24906 143676 24912 143688
rect 24964 143676 24970 143728
rect 23526 143608 23532 143660
rect 23584 143648 23590 143660
rect 25734 143648 25740 143660
rect 23584 143620 25740 143648
rect 23584 143608 23590 143620
rect 25734 143608 25740 143620
rect 25792 143608 25798 143660
rect 26010 143608 26016 143660
rect 26068 143648 26074 143660
rect 26286 143648 26292 143660
rect 26068 143620 26292 143648
rect 26068 143608 26074 143620
rect 26286 143608 26292 143620
rect 26344 143608 26350 143660
rect 27298 143608 27304 143660
rect 27356 143648 27362 143660
rect 27758 143648 27764 143660
rect 27356 143620 27764 143648
rect 27356 143608 27362 143620
rect 27758 143608 27764 143620
rect 27816 143608 27822 143660
rect 28586 143608 28592 143660
rect 28644 143648 28650 143660
rect 29138 143648 29144 143660
rect 28644 143620 29144 143648
rect 28644 143608 28650 143620
rect 29138 143608 29144 143620
rect 29196 143608 29202 143660
rect 30058 143608 30064 143660
rect 30116 143648 30122 143660
rect 30518 143648 30524 143660
rect 30116 143620 30524 143648
rect 30116 143608 30122 143620
rect 30518 143608 30524 143620
rect 30576 143608 30582 143660
rect 31990 143608 31996 143660
rect 32048 143648 32054 143660
rect 32726 143648 32732 143660
rect 32048 143620 32732 143648
rect 32048 143608 32054 143620
rect 32726 143608 32732 143620
rect 32784 143608 32790 143660
rect 34474 143608 34480 143660
rect 34532 143648 34538 143660
rect 34934 143648 34940 143660
rect 34532 143620 34940 143648
rect 34532 143608 34538 143620
rect 34934 143608 34940 143620
rect 34992 143608 34998 143660
rect 35946 143608 35952 143660
rect 36004 143648 36010 143660
rect 36222 143648 36228 143660
rect 36004 143620 36228 143648
rect 36004 143608 36010 143620
rect 36222 143608 36228 143620
rect 36280 143608 36286 143660
rect 37418 143608 37424 143660
rect 37476 143648 37482 143660
rect 38982 143648 38988 143660
rect 37476 143620 38988 143648
rect 37476 143608 37482 143620
rect 38982 143608 38988 143620
rect 39040 143608 39046 143660
rect 43766 143608 43772 143660
rect 43824 143648 43830 143660
rect 44410 143648 44416 143660
rect 43824 143620 44416 143648
rect 43824 143608 43830 143620
rect 44410 143608 44416 143620
rect 44468 143608 44474 143660
rect 110190 143608 110196 143660
rect 110248 143648 110254 143660
rect 110466 143648 110472 143660
rect 110248 143620 110472 143648
rect 110248 143608 110254 143620
rect 110466 143608 110472 143620
rect 110524 143608 110530 143660
rect 112122 143608 112128 143660
rect 112180 143648 112186 143660
rect 112582 143648 112588 143660
rect 112180 143620 112588 143648
rect 112180 143608 112186 143620
rect 112582 143608 112588 143620
rect 112640 143608 112646 143660
rect 114422 143608 114428 143660
rect 114480 143648 114486 143660
rect 114974 143648 114980 143660
rect 114480 143620 114980 143648
rect 114480 143608 114486 143620
rect 114974 143608 114980 143620
rect 115032 143608 115038 143660
rect 115894 143608 115900 143660
rect 115952 143648 115958 143660
rect 116630 143648 116636 143660
rect 115952 143620 116636 143648
rect 115952 143608 115958 143620
rect 116630 143608 116636 143620
rect 116688 143608 116694 143660
rect 192990 143608 192996 143660
rect 193048 143648 193054 143660
rect 193266 143648 193272 143660
rect 193048 143620 193272 143648
rect 193048 143608 193054 143620
rect 193266 143608 193272 143620
rect 193324 143608 193330 143660
rect 194186 143608 194192 143660
rect 194244 143648 194250 143660
rect 194646 143648 194652 143660
rect 194244 143620 194652 143648
rect 194244 143608 194250 143620
rect 194646 143608 194652 143620
rect 194704 143608 194710 143660
rect 20766 143540 20772 143592
rect 20824 143580 20830 143592
rect 25090 143580 25096 143592
rect 20824 143552 25096 143580
rect 20824 143540 20830 143552
rect 25090 143540 25096 143552
rect 25148 143540 25154 143592
rect 34842 143540 34848 143592
rect 34900 143580 34906 143592
rect 35486 143580 35492 143592
rect 34900 143552 35492 143580
rect 34900 143540 34906 143552
rect 35486 143540 35492 143552
rect 35544 143540 35550 143592
rect 35854 143540 35860 143592
rect 35912 143580 35918 143592
rect 37510 143580 37516 143592
rect 35912 143552 37516 143580
rect 35912 143540 35918 143552
rect 37510 143540 37516 143552
rect 37568 143540 37574 143592
rect 43674 143540 43680 143592
rect 43732 143580 43738 143592
rect 47170 143580 47176 143592
rect 43732 143552 47176 143580
rect 43732 143540 43738 143552
rect 47170 143540 47176 143552
rect 47228 143540 47234 143592
rect 99150 143540 99156 143592
rect 99208 143580 99214 143592
rect 106694 143580 106700 143592
rect 99208 143552 106700 143580
rect 99208 143540 99214 143552
rect 106694 143540 106700 143552
rect 106752 143540 106758 143592
rect 114882 143540 114888 143592
rect 114940 143580 114946 143592
rect 115526 143580 115532 143592
rect 114940 143552 115532 143580
rect 114940 143540 114946 143552
rect 115526 143540 115532 143552
rect 115584 143540 115590 143592
rect 116078 143540 116084 143592
rect 116136 143580 116142 143592
rect 117642 143580 117648 143592
rect 116136 143552 117648 143580
rect 116136 143540 116142 143552
rect 117642 143540 117648 143552
rect 117700 143540 117706 143592
rect 99426 143472 99432 143524
rect 99484 143512 99490 143524
rect 106602 143512 106608 143524
rect 99484 143484 106608 143512
rect 99484 143472 99490 143484
rect 106602 143472 106608 143484
rect 106660 143472 106666 143524
rect 113594 143472 113600 143524
rect 113652 143512 113658 143524
rect 114422 143512 114428 143524
rect 113652 143484 114428 143512
rect 113652 143472 113658 143484
rect 114422 143472 114428 143484
rect 114480 143472 114486 143524
rect 183238 143472 183244 143524
rect 183296 143512 183302 143524
rect 190782 143512 190788 143524
rect 183296 143484 190788 143512
rect 183296 143472 183302 143484
rect 190782 143472 190788 143484
rect 190840 143472 190846 143524
rect 38798 143404 38804 143456
rect 38856 143444 38862 143456
rect 40270 143444 40276 143456
rect 38856 143416 40276 143444
rect 38856 143404 38862 143416
rect 40270 143404 40276 143416
rect 40328 143404 40334 143456
rect 99058 143404 99064 143456
rect 99116 143444 99122 143456
rect 107430 143444 107436 143456
rect 99116 143416 107436 143444
rect 99116 143404 99122 143416
rect 107430 143404 107436 143416
rect 107488 143404 107494 143456
rect 183054 143404 183060 143456
rect 183112 143444 183118 143456
rect 192070 143444 192076 143456
rect 183112 143416 192076 143444
rect 183112 143404 183118 143416
rect 192070 143404 192076 143416
rect 192128 143404 192134 143456
rect 22146 143336 22152 143388
rect 22204 143376 22210 143388
rect 25826 143376 25832 143388
rect 22204 143348 25832 143376
rect 22204 143336 22210 143348
rect 25826 143336 25832 143348
rect 25884 143336 25890 143388
rect 44502 143376 44508 143388
rect 25936 143348 44508 143376
rect 20490 143268 20496 143320
rect 20548 143308 20554 143320
rect 25936 143308 25964 143348
rect 44502 143336 44508 143348
rect 44560 143336 44566 143388
rect 98966 143336 98972 143388
rect 99024 143376 99030 143388
rect 107982 143376 107988 143388
rect 99024 143348 107988 143376
rect 99024 143336 99030 143348
rect 107982 143336 107988 143348
rect 108040 143336 108046 143388
rect 183146 143336 183152 143388
rect 183204 143376 183210 143388
rect 191334 143376 191340 143388
rect 183204 143348 191340 143376
rect 183204 143336 183210 143348
rect 191334 143336 191340 143348
rect 191392 143336 191398 143388
rect 191978 143336 191984 143388
rect 192036 143376 192042 143388
rect 215622 143376 215628 143388
rect 192036 143348 215628 143376
rect 192036 143336 192042 143348
rect 215622 143336 215628 143348
rect 215680 143336 215686 143388
rect 20548 143280 25964 143308
rect 20548 143268 20554 143280
rect 37234 143200 37240 143252
rect 37292 143240 37298 143252
rect 39718 143240 39724 143252
rect 37292 143212 39724 143240
rect 37292 143200 37298 143212
rect 39718 143200 39724 143212
rect 39776 143200 39782 143252
rect 45146 143200 45152 143252
rect 45204 143240 45210 143252
rect 46526 143240 46532 143252
rect 45204 143212 46532 143240
rect 45204 143200 45210 143212
rect 46526 143200 46532 143212
rect 46584 143200 46590 143252
rect 35670 143064 35676 143116
rect 35728 143104 35734 143116
rect 36958 143104 36964 143116
rect 35728 143076 36964 143104
rect 35728 143064 35734 143076
rect 36958 143064 36964 143076
rect 37016 143064 37022 143116
rect 117366 143064 117372 143116
rect 117424 143104 117430 143116
rect 118470 143104 118476 143116
rect 117424 143076 118476 143104
rect 117424 143064 117430 143076
rect 118470 143064 118476 143076
rect 118528 143064 118534 143116
rect 31346 142928 31352 142980
rect 31404 142968 31410 142980
rect 31898 142968 31904 142980
rect 31404 142940 31904 142968
rect 31404 142928 31410 142940
rect 31898 142928 31904 142940
rect 31956 142928 31962 142980
rect 38614 142928 38620 142980
rect 38672 142968 38678 142980
rect 41006 142968 41012 142980
rect 38672 142940 41012 142968
rect 38672 142928 38678 142940
rect 41006 142928 41012 142940
rect 41064 142928 41070 142980
rect 45054 142928 45060 142980
rect 45112 142968 45118 142980
rect 45790 142968 45796 142980
rect 45112 142940 45796 142968
rect 45112 142928 45118 142940
rect 45790 142928 45796 142940
rect 45848 142928 45854 142980
rect 98782 142928 98788 142980
rect 98840 142968 98846 142980
rect 103934 142968 103940 142980
rect 98840 142940 103940 142968
rect 98840 142928 98846 142940
rect 103934 142928 103940 142940
rect 103992 142928 103998 142980
rect 117182 142928 117188 142980
rect 117240 142968 117246 142980
rect 117918 142968 117924 142980
rect 117240 142940 117924 142968
rect 117240 142928 117246 142940
rect 117918 142928 117924 142940
rect 117976 142928 117982 142980
rect 99242 142860 99248 142912
rect 99300 142900 99306 142912
rect 105590 142900 105596 142912
rect 99300 142872 105596 142900
rect 99300 142860 99306 142872
rect 105590 142860 105596 142872
rect 105648 142860 105654 142912
rect 23250 142792 23256 142844
rect 23308 142832 23314 142844
rect 25918 142832 25924 142844
rect 23308 142804 25924 142832
rect 23308 142792 23314 142804
rect 25918 142792 25924 142804
rect 25976 142792 25982 142844
rect 37326 142792 37332 142844
rect 37384 142832 37390 142844
rect 38246 142832 38252 142844
rect 37384 142804 38252 142832
rect 37384 142792 37390 142804
rect 38246 142792 38252 142804
rect 38304 142792 38310 142844
rect 99334 142792 99340 142844
rect 99392 142832 99398 142844
rect 105130 142832 105136 142844
rect 99392 142804 105136 142832
rect 99392 142792 99398 142804
rect 105130 142792 105136 142804
rect 105188 142792 105194 142844
rect 200258 142792 200264 142844
rect 200316 142832 200322 142844
rect 200902 142832 200908 142844
rect 200316 142804 200908 142832
rect 200316 142792 200322 142804
rect 200902 142792 200908 142804
rect 200960 142792 200966 142844
rect 99518 142724 99524 142776
rect 99576 142764 99582 142776
rect 104486 142764 104492 142776
rect 99576 142736 104492 142764
rect 99576 142724 99582 142736
rect 104486 142724 104492 142736
rect 104544 142724 104550 142776
rect 68698 142656 68704 142708
rect 68756 142696 68762 142708
rect 69158 142696 69164 142708
rect 68756 142668 69164 142696
rect 68756 142656 68762 142668
rect 69158 142656 69164 142668
rect 69216 142656 69222 142708
rect 167690 142452 167696 142504
rect 167748 142492 167754 142504
rect 169898 142492 169904 142504
rect 167748 142464 169904 142492
rect 167748 142452 167754 142464
rect 169898 142452 169904 142464
rect 169956 142452 169962 142504
rect 49930 140412 49936 140464
rect 49988 140452 49994 140464
rect 53334 140452 53340 140464
rect 49988 140424 53340 140452
rect 49988 140412 49994 140424
rect 53334 140412 53340 140424
rect 53392 140412 53398 140464
rect 134846 140004 134852 140056
rect 134904 140044 134910 140056
rect 143586 140044 143592 140056
rect 134904 140016 143592 140044
rect 134904 140004 134910 140016
rect 143586 140004 143592 140016
rect 143644 140004 143650 140056
rect 49930 139936 49936 139988
rect 49988 139976 49994 139988
rect 58486 139976 58492 139988
rect 49988 139948 58492 139976
rect 49988 139936 49994 139948
rect 58486 139936 58492 139948
rect 58544 139936 58550 139988
rect 135398 139936 135404 139988
rect 135456 139976 135462 139988
rect 143310 139976 143316 139988
rect 135456 139948 143316 139976
rect 135456 139936 135462 139948
rect 143310 139936 143316 139948
rect 143368 139936 143374 139988
rect 135398 138712 135404 138764
rect 135456 138752 135462 138764
rect 139814 138752 139820 138764
rect 135456 138724 139820 138752
rect 135456 138712 135462 138724
rect 139814 138712 139820 138724
rect 139872 138712 139878 138764
rect 49930 138576 49936 138628
rect 49988 138616 49994 138628
rect 58394 138616 58400 138628
rect 49988 138588 58400 138616
rect 49988 138576 49994 138588
rect 58394 138576 58400 138588
rect 58452 138576 58458 138628
rect 134662 138576 134668 138628
rect 134720 138616 134726 138628
rect 139630 138616 139636 138628
rect 134720 138588 139636 138616
rect 134720 138576 134726 138588
rect 139630 138576 139636 138588
rect 139688 138576 139694 138628
rect 92710 138508 92716 138560
rect 92768 138548 92774 138560
rect 100806 138548 100812 138560
rect 92768 138520 100812 138548
rect 92768 138508 92774 138520
rect 100806 138508 100812 138520
rect 100864 138508 100870 138560
rect 177626 138508 177632 138560
rect 177684 138548 177690 138560
rect 185078 138548 185084 138560
rect 177684 138520 185084 138548
rect 177684 138508 177690 138520
rect 185078 138508 185084 138520
rect 185136 138508 185142 138560
rect 49654 138440 49660 138492
rect 49712 138480 49718 138492
rect 58946 138480 58952 138492
rect 49712 138452 58952 138480
rect 49712 138440 49718 138452
rect 58946 138440 58952 138452
rect 59004 138440 59010 138492
rect 92802 138440 92808 138492
rect 92860 138480 92866 138492
rect 100898 138480 100904 138492
rect 92860 138452 100904 138480
rect 92860 138440 92866 138452
rect 100898 138440 100904 138452
rect 100956 138440 100962 138492
rect 177718 138440 177724 138492
rect 177776 138480 177782 138492
rect 184986 138480 184992 138492
rect 177776 138452 184992 138480
rect 177776 138440 177782 138452
rect 184986 138440 184992 138452
rect 185044 138440 185050 138492
rect 97402 137420 97408 137472
rect 97460 137460 97466 137472
rect 101818 137460 101824 137472
rect 97460 137432 101824 137460
rect 97460 137420 97466 137432
rect 101818 137420 101824 137432
rect 101876 137420 101882 137472
rect 134662 137352 134668 137404
rect 134720 137392 134726 137404
rect 139722 137392 139728 137404
rect 134720 137364 139728 137392
rect 134720 137352 134726 137364
rect 139722 137352 139728 137364
rect 139780 137352 139786 137404
rect 49930 137216 49936 137268
rect 49988 137256 49994 137268
rect 58302 137256 58308 137268
rect 49988 137228 58308 137256
rect 49988 137216 49994 137228
rect 58302 137216 58308 137228
rect 58360 137216 58366 137268
rect 98046 137216 98052 137268
rect 98104 137256 98110 137268
rect 101266 137256 101272 137268
rect 98104 137228 101272 137256
rect 98104 137216 98110 137228
rect 101266 137216 101272 137228
rect 101324 137216 101330 137268
rect 181582 137216 181588 137268
rect 181640 137256 181646 137268
rect 185170 137256 185176 137268
rect 181640 137228 185176 137256
rect 181640 137216 181646 137228
rect 185170 137216 185176 137228
rect 185228 137216 185234 137268
rect 50022 137148 50028 137200
rect 50080 137188 50086 137200
rect 58210 137188 58216 137200
rect 50080 137160 58216 137188
rect 50080 137148 50086 137160
rect 58210 137148 58216 137160
rect 58268 137148 58274 137200
rect 135398 137148 135404 137200
rect 135456 137188 135462 137200
rect 143402 137188 143408 137200
rect 135456 137160 143408 137188
rect 135456 137148 135462 137160
rect 143402 137148 143408 137160
rect 143460 137148 143466 137200
rect 182226 137148 182232 137200
rect 182284 137188 182290 137200
rect 185446 137188 185452 137200
rect 182284 137160 185452 137188
rect 182284 137148 182290 137160
rect 185446 137148 185452 137160
rect 185504 137148 185510 137200
rect 92710 137080 92716 137132
rect 92768 137120 92774 137132
rect 101174 137120 101180 137132
rect 92768 137092 101180 137120
rect 92768 137080 92774 137092
rect 101174 137080 101180 137092
rect 101232 137080 101238 137132
rect 177718 137080 177724 137132
rect 177776 137120 177782 137132
rect 185354 137120 185360 137132
rect 177776 137092 185360 137120
rect 177776 137080 177782 137092
rect 185354 137080 185360 137092
rect 185412 137080 185418 137132
rect 92802 137012 92808 137064
rect 92860 137052 92866 137064
rect 101082 137052 101088 137064
rect 92860 137024 101088 137052
rect 92860 137012 92866 137024
rect 101082 137012 101088 137024
rect 101140 137012 101146 137064
rect 139630 137012 139636 137064
rect 139688 137052 139694 137064
rect 143586 137052 143592 137064
rect 139688 137024 143592 137052
rect 139688 137012 139694 137024
rect 143586 137012 143592 137024
rect 143644 137012 143650 137064
rect 177626 137012 177632 137064
rect 177684 137052 177690 137064
rect 185262 137052 185268 137064
rect 177684 137024 185268 137052
rect 177684 137012 177690 137024
rect 185262 137012 185268 137024
rect 185320 137012 185326 137064
rect 92710 136944 92716 136996
rect 92768 136984 92774 136996
rect 97402 136984 97408 136996
rect 92768 136956 97408 136984
rect 92768 136944 92774 136956
rect 97402 136944 97408 136956
rect 97460 136944 97466 136996
rect 139814 136944 139820 136996
rect 139872 136984 139878 136996
rect 143126 136984 143132 136996
rect 139872 136956 143132 136984
rect 139872 136944 139878 136956
rect 143126 136944 143132 136956
rect 143184 136944 143190 136996
rect 139722 136604 139728 136656
rect 139780 136644 139786 136656
rect 143494 136644 143500 136656
rect 139780 136616 143500 136644
rect 139780 136604 139786 136616
rect 143494 136604 143500 136616
rect 143552 136604 143558 136656
rect 177718 136604 177724 136656
rect 177776 136644 177782 136656
rect 181582 136644 181588 136656
rect 177776 136616 181588 136644
rect 177776 136604 177782 136616
rect 181582 136604 181588 136616
rect 181640 136604 181646 136656
rect 51218 135924 51224 135976
rect 51276 135964 51282 135976
rect 56646 135964 56652 135976
rect 51276 135936 56652 135964
rect 51276 135924 51282 135936
rect 56646 135924 56652 135936
rect 56704 135924 56710 135976
rect 135030 135924 135036 135976
rect 135088 135964 135094 135976
rect 143310 135964 143316 135976
rect 135088 135936 143316 135964
rect 135088 135924 135094 135936
rect 143310 135924 143316 135936
rect 143368 135924 143374 135976
rect 51126 135856 51132 135908
rect 51184 135896 51190 135908
rect 56738 135896 56744 135908
rect 51184 135868 56744 135896
rect 51184 135856 51190 135868
rect 56738 135856 56744 135868
rect 56796 135856 56802 135908
rect 97954 135856 97960 135908
rect 98012 135896 98018 135908
rect 101266 135896 101272 135908
rect 98012 135868 101272 135896
rect 98012 135856 98018 135868
rect 101266 135856 101272 135868
rect 101324 135856 101330 135908
rect 135306 135856 135312 135908
rect 135364 135896 135370 135908
rect 143586 135896 143592 135908
rect 135364 135868 143592 135896
rect 135364 135856 135370 135868
rect 143586 135856 143592 135868
rect 143644 135856 143650 135908
rect 182318 135856 182324 135908
rect 182376 135896 182382 135908
rect 185354 135896 185360 135908
rect 182376 135868 185360 135896
rect 182376 135856 182382 135868
rect 185354 135856 185360 135868
rect 185412 135856 185418 135908
rect 51034 135788 51040 135840
rect 51092 135828 51098 135840
rect 56554 135828 56560 135840
rect 51092 135800 56560 135828
rect 51092 135788 51098 135800
rect 56554 135788 56560 135800
rect 56612 135788 56618 135840
rect 98138 135788 98144 135840
rect 98196 135828 98202 135840
rect 101726 135828 101732 135840
rect 98196 135800 101732 135828
rect 98196 135788 98202 135800
rect 101726 135788 101732 135800
rect 101784 135788 101790 135840
rect 135398 135788 135404 135840
rect 135456 135828 135462 135840
rect 143218 135828 143224 135840
rect 135456 135800 143224 135828
rect 135456 135788 135462 135800
rect 143218 135788 143224 135800
rect 143276 135788 143282 135840
rect 181950 135788 181956 135840
rect 182008 135828 182014 135840
rect 185262 135828 185268 135840
rect 182008 135800 185268 135828
rect 182008 135788 182014 135800
rect 185262 135788 185268 135800
rect 185320 135788 185326 135840
rect 92802 135720 92808 135772
rect 92860 135760 92866 135772
rect 101174 135760 101180 135772
rect 92860 135732 101180 135760
rect 92860 135720 92866 135732
rect 101174 135720 101180 135732
rect 101232 135720 101238 135772
rect 177626 135720 177632 135772
rect 177684 135760 177690 135772
rect 185170 135760 185176 135772
rect 177684 135732 185176 135760
rect 177684 135720 177690 135732
rect 185170 135720 185176 135732
rect 185228 135720 185234 135772
rect 92710 135652 92716 135704
rect 92768 135692 92774 135704
rect 98046 135692 98052 135704
rect 92768 135664 98052 135692
rect 92768 135652 92774 135664
rect 98046 135652 98052 135664
rect 98104 135652 98110 135704
rect 177718 135652 177724 135704
rect 177776 135692 177782 135704
rect 182226 135692 182232 135704
rect 177776 135664 182232 135692
rect 177776 135652 177782 135664
rect 182226 135652 182232 135664
rect 182284 135652 182290 135704
rect 56554 135584 56560 135636
rect 56612 135624 56618 135636
rect 58210 135624 58216 135636
rect 56612 135596 58216 135624
rect 56612 135584 56618 135596
rect 58210 135584 58216 135596
rect 58268 135584 58274 135636
rect 56738 135312 56744 135364
rect 56796 135352 56802 135364
rect 58302 135352 58308 135364
rect 56796 135324 58308 135352
rect 56796 135312 56802 135324
rect 58302 135312 58308 135324
rect 58360 135312 58366 135364
rect 134478 134632 134484 134684
rect 134536 134672 134542 134684
rect 136870 134672 136876 134684
rect 134536 134644 136876 134672
rect 134536 134632 134542 134644
rect 136870 134632 136876 134644
rect 136928 134632 136934 134684
rect 51126 134496 51132 134548
rect 51184 134536 51190 134548
rect 59406 134536 59412 134548
rect 51184 134508 56784 134536
rect 59367 134508 59412 134536
rect 51184 134496 51190 134508
rect 51218 134428 51224 134480
rect 51276 134468 51282 134480
rect 56094 134468 56100 134480
rect 51276 134440 56100 134468
rect 51276 134428 51282 134440
rect 56094 134428 56100 134440
rect 56152 134428 56158 134480
rect 56756 134400 56784 134508
rect 59406 134496 59412 134508
rect 59464 134496 59470 134548
rect 134846 134496 134852 134548
rect 134904 134536 134910 134548
rect 139630 134536 139636 134548
rect 134904 134508 139636 134536
rect 134904 134496 134910 134508
rect 139630 134496 139636 134508
rect 139688 134496 139694 134548
rect 58210 134400 58216 134412
rect 56756 134372 58216 134400
rect 58210 134360 58216 134372
rect 58268 134360 58274 134412
rect 92894 134360 92900 134412
rect 92952 134400 92958 134412
rect 101818 134400 101824 134412
rect 92952 134372 101824 134400
rect 92952 134360 92958 134372
rect 101818 134360 101824 134372
rect 101876 134360 101882 134412
rect 177626 134360 177632 134412
rect 177684 134400 177690 134412
rect 185170 134400 185176 134412
rect 177684 134372 185176 134400
rect 177684 134360 177690 134372
rect 185170 134360 185176 134372
rect 185228 134360 185234 134412
rect 92802 134292 92808 134344
rect 92860 134332 92866 134344
rect 98138 134332 98144 134344
rect 92860 134304 98144 134332
rect 92860 134292 92866 134304
rect 98138 134292 98144 134304
rect 98196 134292 98202 134344
rect 177718 134292 177724 134344
rect 177776 134332 177782 134344
rect 181950 134332 181956 134344
rect 177776 134304 181956 134332
rect 177776 134292 177782 134304
rect 181950 134292 181956 134304
rect 182008 134292 182014 134344
rect 56646 134224 56652 134276
rect 56704 134264 56710 134276
rect 58394 134264 58400 134276
rect 56704 134236 58400 134264
rect 56704 134224 56710 134236
rect 58394 134224 58400 134236
rect 58452 134224 58458 134276
rect 92710 134224 92716 134276
rect 92768 134264 92774 134276
rect 97954 134264 97960 134276
rect 92768 134236 97960 134264
rect 92768 134224 92774 134236
rect 97954 134224 97960 134236
rect 98012 134224 98018 134276
rect 177718 134020 177724 134072
rect 177776 134060 177782 134072
rect 182318 134060 182324 134072
rect 177776 134032 182324 134060
rect 177776 134020 177782 134032
rect 182318 134020 182324 134032
rect 182376 134020 182382 134072
rect 139630 133748 139636 133800
rect 139688 133788 139694 133800
rect 142942 133788 142948 133800
rect 139688 133760 142948 133788
rect 139688 133748 139694 133760
rect 142942 133748 142948 133760
rect 143000 133748 143006 133800
rect 56094 133680 56100 133732
rect 56152 133720 56158 133732
rect 58302 133720 58308 133732
rect 56152 133692 58308 133720
rect 56152 133680 56158 133692
rect 58302 133680 58308 133692
rect 58360 133680 58366 133732
rect 50390 133272 50396 133324
rect 50448 133312 50454 133324
rect 56738 133312 56744 133324
rect 50448 133284 56744 133312
rect 50448 133272 50454 133284
rect 56738 133272 56744 133284
rect 56796 133272 56802 133324
rect 51218 133068 51224 133120
rect 51276 133108 51282 133120
rect 55542 133108 55548 133120
rect 51276 133080 55548 133108
rect 51276 133068 51282 133080
rect 55542 133068 55548 133080
rect 55600 133068 55606 133120
rect 135030 133068 135036 133120
rect 135088 133108 135094 133120
rect 138158 133108 138164 133120
rect 135088 133080 138164 133108
rect 135088 133068 135094 133080
rect 138158 133068 138164 133080
rect 138216 133068 138222 133120
rect 51126 133000 51132 133052
rect 51184 133040 51190 133052
rect 51184 133012 56784 133040
rect 51184 133000 51190 133012
rect 56756 132972 56784 133012
rect 135398 133000 135404 133052
rect 135456 133040 135462 133052
rect 135456 133012 139676 133040
rect 135456 133000 135462 133012
rect 58210 132972 58216 132984
rect 56756 132944 58216 132972
rect 58210 132932 58216 132944
rect 58268 132932 58274 132984
rect 59317 132975 59375 132981
rect 59317 132941 59329 132975
rect 59363 132972 59375 132975
rect 59406 132972 59412 132984
rect 59363 132944 59412 132972
rect 59363 132941 59375 132944
rect 59317 132935 59375 132941
rect 59406 132932 59412 132944
rect 59464 132932 59470 132984
rect 92802 132932 92808 132984
rect 92860 132972 92866 132984
rect 101358 132972 101364 132984
rect 92860 132944 101364 132972
rect 92860 132932 92866 132944
rect 101358 132932 101364 132944
rect 101416 132932 101422 132984
rect 139648 132972 139676 133012
rect 143218 132972 143224 132984
rect 139648 132944 143224 132972
rect 143218 132932 143224 132944
rect 143276 132932 143282 132984
rect 177626 132932 177632 132984
rect 177684 132972 177690 132984
rect 185170 132972 185176 132984
rect 177684 132944 185176 132972
rect 177684 132932 177690 132944
rect 185170 132932 185176 132944
rect 185228 132932 185234 132984
rect 56738 132864 56744 132916
rect 56796 132904 56802 132916
rect 58302 132904 58308 132916
rect 56796 132876 58308 132904
rect 56796 132864 56802 132876
rect 58302 132864 58308 132876
rect 58360 132864 58366 132916
rect 92710 132864 92716 132916
rect 92768 132904 92774 132916
rect 100898 132904 100904 132916
rect 92768 132876 100904 132904
rect 92768 132864 92774 132876
rect 100898 132864 100904 132876
rect 100956 132864 100962 132916
rect 177718 132864 177724 132916
rect 177776 132904 177782 132916
rect 185078 132904 185084 132916
rect 177776 132876 185084 132904
rect 177776 132864 177782 132876
rect 185078 132864 185084 132876
rect 185136 132864 185142 132916
rect 136870 132796 136876 132848
rect 136928 132836 136934 132848
rect 143586 132836 143592 132848
rect 136928 132808 143592 132836
rect 136928 132796 136934 132808
rect 143586 132796 143592 132808
rect 143644 132796 143650 132848
rect 135398 131980 135404 132032
rect 135456 132020 135462 132032
rect 138066 132020 138072 132032
rect 135456 131992 138072 132020
rect 135456 131980 135462 131992
rect 138066 131980 138072 131992
rect 138124 131980 138130 132032
rect 135030 131776 135036 131828
rect 135088 131816 135094 131828
rect 137330 131816 137336 131828
rect 135088 131788 137336 131816
rect 135088 131776 135094 131788
rect 137330 131776 137336 131788
rect 137388 131776 137394 131828
rect 51126 131708 51132 131760
rect 51184 131748 51190 131760
rect 55450 131748 55456 131760
rect 51184 131720 55456 131748
rect 51184 131708 51190 131720
rect 55450 131708 55456 131720
rect 55508 131708 55514 131760
rect 51218 131640 51224 131692
rect 51276 131680 51282 131692
rect 58486 131680 58492 131692
rect 51276 131652 58492 131680
rect 51276 131640 51282 131652
rect 58486 131640 58492 131652
rect 58544 131640 58550 131692
rect 135306 131640 135312 131692
rect 135364 131680 135370 131692
rect 135364 131652 140228 131680
rect 135364 131640 135370 131652
rect 92802 131572 92808 131624
rect 92860 131612 92866 131624
rect 101818 131612 101824 131624
rect 92860 131584 101824 131612
rect 92860 131572 92866 131584
rect 101818 131572 101824 131584
rect 101876 131572 101882 131624
rect 140200 131612 140228 131652
rect 142482 131612 142488 131624
rect 140200 131584 142488 131612
rect 142482 131572 142488 131584
rect 142540 131572 142546 131624
rect 177626 131572 177632 131624
rect 177684 131612 177690 131624
rect 185446 131612 185452 131624
rect 177684 131584 185452 131612
rect 177684 131572 177690 131584
rect 185446 131572 185452 131584
rect 185504 131572 185510 131624
rect 92710 131504 92716 131556
rect 92768 131544 92774 131556
rect 101726 131544 101732 131556
rect 92768 131516 101732 131544
rect 92768 131504 92774 131516
rect 101726 131504 101732 131516
rect 101784 131504 101790 131556
rect 138158 131504 138164 131556
rect 138216 131544 138222 131556
rect 143586 131544 143592 131556
rect 138216 131516 143592 131544
rect 138216 131504 138222 131516
rect 143586 131504 143592 131516
rect 143644 131504 143650 131556
rect 177718 131504 177724 131556
rect 177776 131544 177782 131556
rect 185814 131544 185820 131556
rect 177776 131516 185820 131544
rect 177776 131504 177782 131516
rect 185814 131504 185820 131516
rect 185872 131504 185878 131556
rect 55542 131368 55548 131420
rect 55600 131408 55606 131420
rect 58210 131408 58216 131420
rect 55600 131380 58216 131408
rect 55600 131368 55606 131380
rect 58210 131368 58216 131380
rect 58268 131368 58274 131420
rect 55450 131096 55456 131148
rect 55508 131136 55514 131148
rect 58302 131136 58308 131148
rect 55508 131108 58308 131136
rect 55508 131096 55514 131108
rect 58302 131096 58308 131108
rect 58360 131096 58366 131148
rect 135398 130552 135404 130604
rect 135456 130592 135462 130604
rect 137606 130592 137612 130604
rect 135456 130564 137612 130592
rect 135456 130552 135462 130564
rect 137606 130552 137612 130564
rect 137664 130552 137670 130604
rect 51126 130416 51132 130468
rect 51184 130456 51190 130468
rect 56738 130456 56744 130468
rect 51184 130428 56744 130456
rect 51184 130416 51190 130428
rect 56738 130416 56744 130428
rect 56796 130416 56802 130468
rect 51218 130348 51224 130400
rect 51276 130388 51282 130400
rect 56554 130388 56560 130400
rect 51276 130360 56560 130388
rect 51276 130348 51282 130360
rect 56554 130348 56560 130360
rect 56612 130348 56618 130400
rect 50206 130280 50212 130332
rect 50264 130320 50270 130332
rect 50264 130292 56784 130320
rect 50264 130280 50270 130292
rect 56756 130184 56784 130292
rect 135030 130280 135036 130332
rect 135088 130320 135094 130332
rect 137330 130320 137336 130332
rect 135088 130292 137336 130320
rect 135088 130280 135094 130292
rect 137330 130280 137336 130292
rect 137388 130280 137394 130332
rect 92802 130212 92808 130264
rect 92860 130252 92866 130264
rect 101634 130252 101640 130264
rect 92860 130224 101640 130252
rect 92860 130212 92866 130224
rect 101634 130212 101640 130224
rect 101692 130212 101698 130264
rect 138066 130212 138072 130264
rect 138124 130252 138130 130264
rect 143586 130252 143592 130264
rect 138124 130224 143592 130252
rect 138124 130212 138130 130224
rect 143586 130212 143592 130224
rect 143644 130212 143650 130264
rect 177626 130212 177632 130264
rect 177684 130252 177690 130264
rect 185538 130252 185544 130264
rect 177684 130224 185544 130252
rect 177684 130212 177690 130224
rect 185538 130212 185544 130224
rect 185596 130212 185602 130264
rect 58210 130184 58216 130196
rect 56756 130156 58216 130184
rect 58210 130144 58216 130156
rect 58268 130144 58274 130196
rect 92710 130144 92716 130196
rect 92768 130184 92774 130196
rect 101450 130184 101456 130196
rect 92768 130156 101456 130184
rect 92768 130144 92774 130156
rect 101450 130144 101456 130156
rect 101508 130144 101514 130196
rect 137238 130144 137244 130196
rect 137296 130184 137302 130196
rect 143034 130184 143040 130196
rect 137296 130156 143040 130184
rect 137296 130144 137302 130156
rect 143034 130144 143040 130156
rect 143092 130144 143098 130196
rect 177718 130144 177724 130196
rect 177776 130184 177782 130196
rect 185722 130184 185728 130196
rect 177776 130156 185728 130184
rect 177776 130144 177782 130156
rect 185722 130144 185728 130156
rect 185780 130144 185786 130196
rect 135306 129328 135312 129380
rect 135364 129368 135370 129380
rect 137698 129368 137704 129380
rect 135364 129340 137704 129368
rect 135364 129328 135370 129340
rect 137698 129328 137704 129340
rect 137756 129328 137762 129380
rect 51218 128988 51224 129040
rect 51276 129028 51282 129040
rect 56646 129028 56652 129040
rect 51276 129000 56652 129028
rect 51276 128988 51282 129000
rect 56646 128988 56652 129000
rect 56704 128988 56710 129040
rect 51126 128920 51132 128972
rect 51184 128960 51190 128972
rect 56370 128960 56376 128972
rect 51184 128932 56376 128960
rect 51184 128920 51190 128932
rect 56370 128920 56376 128932
rect 56428 128920 56434 128972
rect 135398 128920 135404 128972
rect 135456 128960 135462 128972
rect 135456 128932 139676 128960
rect 135456 128920 135462 128932
rect 92894 128852 92900 128904
rect 92952 128892 92958 128904
rect 101358 128892 101364 128904
rect 92952 128864 101364 128892
rect 92952 128852 92958 128864
rect 101358 128852 101364 128864
rect 101416 128852 101422 128904
rect 139648 128892 139676 128932
rect 143126 128892 143132 128904
rect 139648 128864 143132 128892
rect 143126 128852 143132 128864
rect 143184 128852 143190 128904
rect 177718 128852 177724 128904
rect 177776 128892 177782 128904
rect 185262 128892 185268 128904
rect 177776 128864 185268 128892
rect 177776 128852 177782 128864
rect 185262 128852 185268 128864
rect 185320 128852 185326 128904
rect 56738 128784 56744 128836
rect 56796 128824 56802 128836
rect 58210 128824 58216 128836
rect 56796 128796 58216 128824
rect 56796 128784 56802 128796
rect 58210 128784 58216 128796
rect 58268 128784 58274 128836
rect 92802 128784 92808 128836
rect 92860 128824 92866 128836
rect 101818 128824 101824 128836
rect 92860 128796 101824 128824
rect 92860 128784 92866 128796
rect 101818 128784 101824 128796
rect 101876 128784 101882 128836
rect 137330 128784 137336 128836
rect 137388 128824 137394 128836
rect 142758 128824 142764 128836
rect 137388 128796 142764 128824
rect 137388 128784 137394 128796
rect 142758 128784 142764 128796
rect 142816 128784 142822 128836
rect 177810 128784 177816 128836
rect 177868 128824 177874 128836
rect 185170 128824 185176 128836
rect 177868 128796 185176 128824
rect 177868 128784 177874 128796
rect 185170 128784 185176 128796
rect 185228 128784 185234 128836
rect 56554 128716 56560 128768
rect 56612 128756 56618 128768
rect 58394 128756 58400 128768
rect 56612 128728 58400 128756
rect 56612 128716 56618 128728
rect 58394 128716 58400 128728
rect 58452 128716 58458 128768
rect 92710 128716 92716 128768
rect 92768 128756 92774 128768
rect 101726 128756 101732 128768
rect 92768 128728 101732 128756
rect 92768 128716 92774 128728
rect 101726 128716 101732 128728
rect 101784 128716 101790 128768
rect 137606 128716 137612 128768
rect 137664 128756 137670 128768
rect 143586 128756 143592 128768
rect 137664 128728 143592 128756
rect 137664 128716 137670 128728
rect 143586 128716 143592 128728
rect 143644 128716 143650 128768
rect 177626 128716 177632 128768
rect 177684 128756 177690 128768
rect 185354 128756 185360 128768
rect 177684 128728 185360 128756
rect 177684 128716 177690 128728
rect 185354 128716 185360 128728
rect 185412 128716 185418 128768
rect 56370 128512 56376 128564
rect 56428 128552 56434 128564
rect 58302 128552 58308 128564
rect 56428 128524 58308 128552
rect 56428 128512 56434 128524
rect 58302 128512 58308 128524
rect 58360 128512 58366 128564
rect 135306 127696 135312 127748
rect 135364 127736 135370 127748
rect 137606 127736 137612 127748
rect 135364 127708 137612 127736
rect 135364 127696 135370 127708
rect 137606 127696 137612 127708
rect 137664 127696 137670 127748
rect 50758 127560 50764 127612
rect 50816 127600 50822 127612
rect 58210 127600 58216 127612
rect 50816 127572 58216 127600
rect 50816 127560 50822 127572
rect 58210 127560 58216 127572
rect 58268 127560 58274 127612
rect 134662 127560 134668 127612
rect 134720 127600 134726 127612
rect 137422 127600 137428 127612
rect 134720 127572 137428 127600
rect 134720 127560 134726 127572
rect 137422 127560 137428 127572
rect 137480 127560 137486 127612
rect 51218 127492 51224 127544
rect 51276 127532 51282 127544
rect 58302 127532 58308 127544
rect 51276 127504 58308 127532
rect 51276 127492 51282 127504
rect 58302 127492 58308 127504
rect 58360 127492 58366 127544
rect 135398 127492 135404 127544
rect 135456 127532 135462 127544
rect 135456 127504 139676 127532
rect 135456 127492 135462 127504
rect 56646 127424 56652 127476
rect 56704 127464 56710 127476
rect 58394 127464 58400 127476
rect 56704 127436 58400 127464
rect 56704 127424 56710 127436
rect 58394 127424 58400 127436
rect 58452 127424 58458 127476
rect 92802 127424 92808 127476
rect 92860 127464 92866 127476
rect 100990 127464 100996 127476
rect 92860 127436 100996 127464
rect 92860 127424 92866 127436
rect 100990 127424 100996 127436
rect 101048 127424 101054 127476
rect 139648 127464 139676 127504
rect 143310 127464 143316 127476
rect 139648 127436 143316 127464
rect 143310 127424 143316 127436
rect 143368 127424 143374 127476
rect 177718 127424 177724 127476
rect 177776 127464 177782 127476
rect 185170 127464 185176 127476
rect 177776 127436 185176 127464
rect 177776 127424 177782 127436
rect 185170 127424 185176 127436
rect 185228 127424 185234 127476
rect 216174 127424 216180 127476
rect 216232 127464 216238 127476
rect 222338 127464 222344 127476
rect 216232 127436 222344 127464
rect 216232 127424 216238 127436
rect 222338 127424 222344 127436
rect 222396 127424 222402 127476
rect 92710 127356 92716 127408
rect 92768 127396 92774 127408
rect 101266 127396 101272 127408
rect 92768 127368 101272 127396
rect 92768 127356 92774 127368
rect 101266 127356 101272 127368
rect 101324 127356 101330 127408
rect 137698 127356 137704 127408
rect 137756 127396 137762 127408
rect 142482 127396 142488 127408
rect 137756 127368 142488 127396
rect 137756 127356 137762 127368
rect 142482 127356 142488 127368
rect 142540 127356 142546 127408
rect 177166 127356 177172 127408
rect 177224 127396 177230 127408
rect 185446 127396 185452 127408
rect 177224 127368 185452 127396
rect 177224 127356 177230 127368
rect 185446 127356 185452 127368
rect 185504 127356 185510 127408
rect 50390 126336 50396 126388
rect 50448 126376 50454 126388
rect 56738 126376 56744 126388
rect 50448 126348 56744 126376
rect 50448 126336 50454 126348
rect 56738 126336 56744 126348
rect 56796 126336 56802 126388
rect 51218 126200 51224 126252
rect 51276 126240 51282 126252
rect 56094 126240 56100 126252
rect 51276 126212 56100 126240
rect 51276 126200 51282 126212
rect 56094 126200 56100 126212
rect 56152 126200 56158 126252
rect 98046 126200 98052 126252
rect 98104 126240 98110 126252
rect 101266 126240 101272 126252
rect 98104 126212 101272 126240
rect 98104 126200 98110 126212
rect 101266 126200 101272 126212
rect 101324 126200 101330 126252
rect 182226 126200 182232 126252
rect 182284 126240 182290 126252
rect 185446 126240 185452 126252
rect 182284 126212 185452 126240
rect 182284 126200 182290 126212
rect 185446 126200 185452 126212
rect 185504 126200 185510 126252
rect 50206 126132 50212 126184
rect 50264 126172 50270 126184
rect 58210 126172 58216 126184
rect 50264 126144 58216 126172
rect 50264 126132 50270 126144
rect 58210 126132 58216 126144
rect 58268 126132 58274 126184
rect 98138 126132 98144 126184
rect 98196 126172 98202 126184
rect 100990 126172 100996 126184
rect 98196 126144 100996 126172
rect 98196 126132 98202 126144
rect 100990 126132 100996 126144
rect 101048 126132 101054 126184
rect 182318 126132 182324 126184
rect 182376 126172 182382 126184
rect 185170 126172 185176 126184
rect 182376 126144 185176 126172
rect 182376 126132 182382 126144
rect 185170 126132 185176 126144
rect 185228 126132 185234 126184
rect 92710 126064 92716 126116
rect 92768 126104 92774 126116
rect 101174 126104 101180 126116
rect 92768 126076 101180 126104
rect 92768 126064 92774 126076
rect 101174 126064 101180 126076
rect 101232 126064 101238 126116
rect 137606 126064 137612 126116
rect 137664 126104 137670 126116
rect 143494 126104 143500 126116
rect 137664 126076 143500 126104
rect 137664 126064 137670 126076
rect 143494 126064 143500 126076
rect 143552 126064 143558 126116
rect 177718 126064 177724 126116
rect 177776 126104 177782 126116
rect 185354 126104 185360 126116
rect 177776 126076 185360 126104
rect 177776 126064 177782 126076
rect 185354 126064 185360 126076
rect 185412 126064 185418 126116
rect 92802 125996 92808 126048
rect 92860 126036 92866 126048
rect 101082 126036 101088 126048
rect 92860 126008 101088 126036
rect 92860 125996 92866 126008
rect 101082 125996 101088 126008
rect 101140 125996 101146 126048
rect 137422 125996 137428 126048
rect 137480 126036 137486 126048
rect 143586 126036 143592 126048
rect 137480 126008 143592 126036
rect 137480 125996 137486 126008
rect 143586 125996 143592 126008
rect 143644 125996 143650 126048
rect 177626 125996 177632 126048
rect 177684 126036 177690 126048
rect 185262 126036 185268 126048
rect 177684 126008 185268 126036
rect 177684 125996 177690 126008
rect 185262 125996 185268 126008
rect 185320 125996 185326 126048
rect 135398 125384 135404 125436
rect 135456 125424 135462 125436
rect 137606 125424 137612 125436
rect 135456 125396 137612 125424
rect 135456 125384 135462 125396
rect 137606 125384 137612 125396
rect 137664 125384 137670 125436
rect 51126 124840 51132 124892
rect 51184 124880 51190 124892
rect 55450 124880 55456 124892
rect 51184 124852 55456 124880
rect 51184 124840 51190 124852
rect 55450 124840 55456 124852
rect 55508 124840 55514 124892
rect 135398 124840 135404 124892
rect 135456 124880 135462 124892
rect 136870 124880 136876 124892
rect 135456 124852 136876 124880
rect 135456 124840 135462 124852
rect 136870 124840 136876 124852
rect 136928 124840 136934 124892
rect 51218 124772 51224 124824
rect 51276 124812 51282 124824
rect 58394 124812 58400 124824
rect 51276 124784 58400 124812
rect 51276 124772 51282 124784
rect 58394 124772 58400 124784
rect 58452 124772 58458 124824
rect 135214 124772 135220 124824
rect 135272 124812 135278 124824
rect 142758 124812 142764 124824
rect 135272 124784 142764 124812
rect 135272 124772 135278 124784
rect 142758 124772 142764 124784
rect 142816 124772 142822 124824
rect 55450 124704 55456 124756
rect 55508 124744 55514 124756
rect 58210 124744 58216 124756
rect 55508 124716 58216 124744
rect 55508 124704 55514 124716
rect 58210 124704 58216 124716
rect 58268 124704 58274 124756
rect 92894 124704 92900 124756
rect 92952 124744 92958 124756
rect 100990 124744 100996 124756
rect 92952 124716 100996 124744
rect 92952 124704 92958 124716
rect 100990 124704 100996 124716
rect 101048 124704 101054 124756
rect 135582 124704 135588 124756
rect 135640 124744 135646 124756
rect 143586 124744 143592 124756
rect 135640 124716 143592 124744
rect 135640 124704 135646 124716
rect 143586 124704 143592 124716
rect 143644 124704 143650 124756
rect 177626 124704 177632 124756
rect 177684 124744 177690 124756
rect 185170 124744 185176 124756
rect 177684 124716 185176 124744
rect 177684 124704 177690 124716
rect 185170 124704 185176 124716
rect 185228 124704 185234 124756
rect 56738 124636 56744 124688
rect 56796 124676 56802 124688
rect 58302 124676 58308 124688
rect 56796 124648 58308 124676
rect 56796 124636 56802 124648
rect 58302 124636 58308 124648
rect 58360 124636 58366 124688
rect 92710 124636 92716 124688
rect 92768 124676 92774 124688
rect 98046 124676 98052 124688
rect 92768 124648 98052 124676
rect 92768 124636 92774 124648
rect 98046 124636 98052 124648
rect 98104 124636 98110 124688
rect 177718 124636 177724 124688
rect 177776 124676 177782 124688
rect 182226 124676 182232 124688
rect 177776 124648 182232 124676
rect 177776 124636 177782 124648
rect 182226 124636 182232 124648
rect 182284 124636 182290 124688
rect 56094 124568 56100 124620
rect 56152 124608 56158 124620
rect 58486 124608 58492 124620
rect 56152 124580 58492 124608
rect 56152 124568 56158 124580
rect 58486 124568 58492 124580
rect 58544 124568 58550 124620
rect 92802 124568 92808 124620
rect 92860 124608 92866 124620
rect 98138 124608 98144 124620
rect 92860 124580 98144 124608
rect 92860 124568 92866 124580
rect 98138 124568 98144 124580
rect 98196 124568 98202 124620
rect 135490 124364 135496 124416
rect 135548 124404 135554 124416
rect 142482 124404 142488 124416
rect 135548 124376 142488 124404
rect 135548 124364 135554 124376
rect 142482 124364 142488 124376
rect 142540 124364 142546 124416
rect 177166 124364 177172 124416
rect 177224 124404 177230 124416
rect 182318 124404 182324 124416
rect 177224 124376 182324 124404
rect 177224 124364 177230 124376
rect 182318 124364 182324 124376
rect 182376 124364 182382 124416
rect 51218 123616 51224 123668
rect 51276 123656 51282 123668
rect 55542 123656 55548 123668
rect 51276 123628 55548 123656
rect 51276 123616 51282 123628
rect 55542 123616 55548 123628
rect 55600 123616 55606 123668
rect 135030 123616 135036 123668
rect 135088 123656 135094 123668
rect 137422 123656 137428 123668
rect 135088 123628 137428 123656
rect 135088 123616 135094 123628
rect 137422 123616 137428 123628
rect 137480 123616 137486 123668
rect 51218 123480 51224 123532
rect 51276 123520 51282 123532
rect 55450 123520 55456 123532
rect 51276 123492 55456 123520
rect 51276 123480 51282 123492
rect 55450 123480 55456 123492
rect 55508 123480 55514 123532
rect 50206 123344 50212 123396
rect 50264 123384 50270 123396
rect 50264 123356 56784 123384
rect 50264 123344 50270 123356
rect 56756 123248 56784 123356
rect 134110 123344 134116 123396
rect 134168 123384 134174 123396
rect 138158 123384 138164 123396
rect 134168 123356 138164 123384
rect 134168 123344 134174 123356
rect 138158 123344 138164 123356
rect 138216 123344 138222 123396
rect 92802 123276 92808 123328
rect 92860 123316 92866 123328
rect 101082 123316 101088 123328
rect 92860 123288 101088 123316
rect 92860 123276 92866 123288
rect 101082 123276 101088 123288
rect 101140 123276 101146 123328
rect 137606 123276 137612 123328
rect 137664 123316 137670 123328
rect 143586 123316 143592 123328
rect 137664 123288 143592 123316
rect 137664 123276 137670 123288
rect 143586 123276 143592 123288
rect 143644 123276 143650 123328
rect 177626 123276 177632 123328
rect 177684 123316 177690 123328
rect 185354 123316 185360 123328
rect 177684 123288 185360 123316
rect 177684 123276 177690 123288
rect 185354 123276 185360 123288
rect 185412 123276 185418 123328
rect 58210 123248 58216 123260
rect 56756 123220 58216 123248
rect 58210 123208 58216 123220
rect 58268 123208 58274 123260
rect 92710 123208 92716 123260
rect 92768 123248 92774 123260
rect 101266 123248 101272 123260
rect 92768 123220 101272 123248
rect 92768 123208 92774 123220
rect 101266 123208 101272 123220
rect 101324 123208 101330 123260
rect 177718 123208 177724 123260
rect 177776 123248 177782 123260
rect 185446 123248 185452 123260
rect 177776 123220 185452 123248
rect 177776 123208 177782 123220
rect 185446 123208 185452 123220
rect 185504 123208 185510 123260
rect 136870 122800 136876 122852
rect 136928 122840 136934 122852
rect 143586 122840 143592 122852
rect 136928 122812 143592 122840
rect 136928 122800 136934 122812
rect 143586 122800 143592 122812
rect 143644 122800 143650 122852
rect 135214 122528 135220 122580
rect 135272 122568 135278 122580
rect 137882 122568 137888 122580
rect 135272 122540 137888 122568
rect 135272 122528 135278 122540
rect 137882 122528 137888 122540
rect 137940 122528 137946 122580
rect 135214 122188 135220 122240
rect 135272 122228 135278 122240
rect 137790 122228 137796 122240
rect 135272 122200 137796 122228
rect 135272 122188 135278 122200
rect 137790 122188 137796 122200
rect 137848 122188 137854 122240
rect 51218 122120 51224 122172
rect 51276 122160 51282 122172
rect 55726 122160 55732 122172
rect 51276 122132 55732 122160
rect 51276 122120 51282 122132
rect 55726 122120 55732 122132
rect 55784 122120 55790 122172
rect 51126 121984 51132 122036
rect 51184 122024 51190 122036
rect 55634 122024 55640 122036
rect 51184 121996 55640 122024
rect 51184 121984 51190 121996
rect 55634 121984 55640 121996
rect 55692 121984 55698 122036
rect 92802 121916 92808 121968
rect 92860 121956 92866 121968
rect 100990 121956 100996 121968
rect 92860 121928 100996 121956
rect 92860 121916 92866 121928
rect 100990 121916 100996 121928
rect 101048 121916 101054 121968
rect 137422 121916 137428 121968
rect 137480 121956 137486 121968
rect 142758 121956 142764 121968
rect 137480 121928 142764 121956
rect 137480 121916 137486 121928
rect 142758 121916 142764 121928
rect 142816 121916 142822 121968
rect 177718 121916 177724 121968
rect 177776 121956 177782 121968
rect 185814 121956 185820 121968
rect 177776 121928 185820 121956
rect 177776 121916 177782 121928
rect 185814 121916 185820 121928
rect 185872 121916 185878 121968
rect 92710 121848 92716 121900
rect 92768 121888 92774 121900
rect 101174 121888 101180 121900
rect 92768 121860 101180 121888
rect 92768 121848 92774 121860
rect 101174 121848 101180 121860
rect 101232 121848 101238 121900
rect 138158 121848 138164 121900
rect 138216 121888 138222 121900
rect 143034 121888 143040 121900
rect 138216 121860 143040 121888
rect 138216 121848 138222 121860
rect 143034 121848 143040 121860
rect 143092 121848 143098 121900
rect 177350 121848 177356 121900
rect 177408 121888 177414 121900
rect 185262 121888 185268 121900
rect 177408 121860 185268 121888
rect 177408 121848 177414 121860
rect 185262 121848 185268 121860
rect 185320 121848 185326 121900
rect 55542 121780 55548 121832
rect 55600 121820 55606 121832
rect 58210 121820 58216 121832
rect 55600 121792 58216 121820
rect 55600 121780 55606 121792
rect 58210 121780 58216 121792
rect 58268 121780 58274 121832
rect 55450 121508 55456 121560
rect 55508 121548 55514 121560
rect 58210 121548 58216 121560
rect 55508 121520 58216 121548
rect 55508 121508 55514 121520
rect 58210 121508 58216 121520
rect 58268 121508 58274 121560
rect 97494 120760 97500 120812
rect 97552 120800 97558 120812
rect 100990 120800 100996 120812
rect 97552 120772 100996 120800
rect 97552 120760 97558 120772
rect 100990 120760 100996 120772
rect 101048 120760 101054 120812
rect 134846 120760 134852 120812
rect 134904 120800 134910 120812
rect 137330 120800 137336 120812
rect 134904 120772 137336 120800
rect 134904 120760 134910 120772
rect 137330 120760 137336 120772
rect 137388 120760 137394 120812
rect 182042 120760 182048 120812
rect 182100 120800 182106 120812
rect 185354 120800 185360 120812
rect 182100 120772 185360 120800
rect 182100 120760 182106 120772
rect 185354 120760 185360 120772
rect 185412 120760 185418 120812
rect 51218 120692 51224 120744
rect 51276 120732 51282 120744
rect 58486 120732 58492 120744
rect 51276 120704 58492 120732
rect 51276 120692 51282 120704
rect 58486 120692 58492 120704
rect 58544 120692 58550 120744
rect 97954 120692 97960 120744
rect 98012 120732 98018 120744
rect 101174 120732 101180 120744
rect 98012 120704 101180 120732
rect 98012 120692 98018 120704
rect 101174 120692 101180 120704
rect 101232 120692 101238 120744
rect 134662 120692 134668 120744
rect 134720 120732 134726 120744
rect 137606 120732 137612 120744
rect 134720 120704 137612 120732
rect 134720 120692 134726 120704
rect 137606 120692 137612 120704
rect 137664 120692 137670 120744
rect 182318 120692 182324 120744
rect 182376 120732 182382 120744
rect 185262 120732 185268 120744
rect 182376 120704 185268 120732
rect 182376 120692 182382 120704
rect 185262 120692 185268 120704
rect 185320 120692 185326 120744
rect 51126 120624 51132 120676
rect 51184 120664 51190 120676
rect 58302 120664 58308 120676
rect 51184 120636 58308 120664
rect 51184 120624 51190 120636
rect 58302 120624 58308 120636
rect 58360 120624 58366 120676
rect 98138 120624 98144 120676
rect 98196 120664 98202 120676
rect 100990 120664 100996 120676
rect 98196 120636 100996 120664
rect 98196 120624 98202 120636
rect 100990 120624 100996 120636
rect 101048 120624 101054 120676
rect 135398 120624 135404 120676
rect 135456 120664 135462 120676
rect 136870 120664 136876 120676
rect 135456 120636 136876 120664
rect 135456 120624 135462 120636
rect 136870 120624 136876 120636
rect 136928 120624 136934 120676
rect 181582 120624 181588 120676
rect 181640 120664 181646 120676
rect 185170 120664 185176 120676
rect 181640 120636 185176 120664
rect 181640 120624 181646 120636
rect 185170 120624 185176 120636
rect 185228 120624 185234 120676
rect 55634 120556 55640 120608
rect 55692 120596 55698 120608
rect 58210 120596 58216 120608
rect 55692 120568 58216 120596
rect 55692 120556 55698 120568
rect 58210 120556 58216 120568
rect 58268 120556 58274 120608
rect 92802 120556 92808 120608
rect 92860 120596 92866 120608
rect 101082 120596 101088 120608
rect 92860 120568 101088 120596
rect 92860 120556 92866 120568
rect 101082 120556 101088 120568
rect 101140 120556 101146 120608
rect 137882 120556 137888 120608
rect 137940 120596 137946 120608
rect 142942 120596 142948 120608
rect 137940 120568 142948 120596
rect 137940 120556 137946 120568
rect 142942 120556 142948 120568
rect 143000 120556 143006 120608
rect 177626 120556 177632 120608
rect 177684 120596 177690 120608
rect 185906 120596 185912 120608
rect 177684 120568 185912 120596
rect 177684 120556 177690 120568
rect 185906 120556 185912 120568
rect 185964 120556 185970 120608
rect 55726 120488 55732 120540
rect 55784 120528 55790 120540
rect 58394 120528 58400 120540
rect 55784 120500 58400 120528
rect 55784 120488 55790 120500
rect 58394 120488 58400 120500
rect 58452 120488 58458 120540
rect 92710 120488 92716 120540
rect 92768 120528 92774 120540
rect 101266 120528 101272 120540
rect 92768 120500 101272 120528
rect 92768 120488 92774 120500
rect 101266 120488 101272 120500
rect 101324 120488 101330 120540
rect 137790 120488 137796 120540
rect 137848 120528 137854 120540
rect 143586 120528 143592 120540
rect 137848 120500 143592 120528
rect 137848 120488 137854 120500
rect 143586 120488 143592 120500
rect 143644 120488 143650 120540
rect 177718 120488 177724 120540
rect 177776 120528 177782 120540
rect 185630 120528 185636 120540
rect 177776 120500 185636 120528
rect 177776 120488 177782 120500
rect 185630 120488 185636 120500
rect 185688 120488 185694 120540
rect 134294 120080 134300 120132
rect 134352 120120 134358 120132
rect 136962 120120 136968 120132
rect 134352 120092 136968 120120
rect 134352 120080 134358 120092
rect 136962 120080 136968 120092
rect 137020 120080 137026 120132
rect 51218 119536 51224 119588
rect 51276 119576 51282 119588
rect 56738 119576 56744 119588
rect 51276 119548 56744 119576
rect 51276 119536 51282 119548
rect 56738 119536 56744 119548
rect 56796 119536 56802 119588
rect 135398 119536 135404 119588
rect 135456 119576 135462 119588
rect 137698 119576 137704 119588
rect 135456 119548 137704 119576
rect 135456 119536 135462 119548
rect 137698 119536 137704 119548
rect 137756 119536 137762 119588
rect 51218 119400 51224 119452
rect 51276 119440 51282 119452
rect 56278 119440 56284 119452
rect 51276 119412 56284 119440
rect 51276 119400 51282 119412
rect 56278 119400 56284 119412
rect 56336 119400 56342 119452
rect 97862 119332 97868 119384
rect 97920 119372 97926 119384
rect 101082 119372 101088 119384
rect 97920 119344 101088 119372
rect 97920 119332 97926 119344
rect 101082 119332 101088 119344
rect 101140 119332 101146 119384
rect 182134 119332 182140 119384
rect 182192 119372 182198 119384
rect 185262 119372 185268 119384
rect 182192 119344 185268 119372
rect 182192 119332 182198 119344
rect 185262 119332 185268 119344
rect 185320 119332 185326 119384
rect 50206 119264 50212 119316
rect 50264 119304 50270 119316
rect 50264 119276 56784 119304
rect 50264 119264 50270 119276
rect 56756 119168 56784 119276
rect 98046 119264 98052 119316
rect 98104 119304 98110 119316
rect 100990 119304 100996 119316
rect 98104 119276 100996 119304
rect 98104 119264 98110 119276
rect 100990 119264 100996 119276
rect 101048 119264 101054 119316
rect 182226 119264 182232 119316
rect 182284 119304 182290 119316
rect 185170 119304 185176 119316
rect 182284 119276 185176 119304
rect 182284 119264 182290 119276
rect 185170 119264 185176 119276
rect 185228 119264 185234 119316
rect 92894 119196 92900 119248
rect 92952 119236 92958 119248
rect 98138 119236 98144 119248
rect 92952 119208 98144 119236
rect 92952 119196 92958 119208
rect 98138 119196 98144 119208
rect 98196 119196 98202 119248
rect 137330 119196 137336 119248
rect 137388 119236 137394 119248
rect 143586 119236 143592 119248
rect 137388 119208 143592 119236
rect 137388 119196 137394 119208
rect 143586 119196 143592 119208
rect 143644 119196 143650 119248
rect 58210 119168 58216 119180
rect 56756 119140 58216 119168
rect 58210 119128 58216 119140
rect 58268 119128 58274 119180
rect 92802 119128 92808 119180
rect 92860 119168 92866 119180
rect 97954 119168 97960 119180
rect 92860 119140 97960 119168
rect 92860 119128 92866 119140
rect 97954 119128 97960 119140
rect 98012 119128 98018 119180
rect 137606 119128 137612 119180
rect 137664 119168 137670 119180
rect 143034 119168 143040 119180
rect 137664 119140 143040 119168
rect 137664 119128 137670 119140
rect 143034 119128 143040 119140
rect 143092 119128 143098 119180
rect 92710 119060 92716 119112
rect 92768 119100 92774 119112
rect 97494 119100 97500 119112
rect 92768 119072 97500 119100
rect 92768 119060 92774 119072
rect 97494 119060 97500 119072
rect 97552 119060 97558 119112
rect 136870 119060 136876 119112
rect 136928 119100 136934 119112
rect 143310 119100 143316 119112
rect 136928 119072 143316 119100
rect 136928 119060 136934 119072
rect 143310 119060 143316 119072
rect 143368 119060 143374 119112
rect 177718 119060 177724 119112
rect 177776 119100 177782 119112
rect 182042 119100 182048 119112
rect 177776 119072 182048 119100
rect 177776 119060 177782 119072
rect 182042 119060 182048 119072
rect 182100 119060 182106 119112
rect 177718 118924 177724 118976
rect 177776 118964 177782 118976
rect 181582 118964 181588 118976
rect 177776 118936 181588 118964
rect 177776 118924 177782 118936
rect 181582 118924 181588 118936
rect 181640 118924 181646 118976
rect 177626 118788 177632 118840
rect 177684 118828 177690 118840
rect 182318 118828 182324 118840
rect 177684 118800 182324 118828
rect 177684 118788 177690 118800
rect 182318 118788 182324 118800
rect 182376 118788 182382 118840
rect 134478 118176 134484 118228
rect 134536 118216 134542 118228
rect 137606 118216 137612 118228
rect 134536 118188 137612 118216
rect 134536 118176 134542 118188
rect 137606 118176 137612 118188
rect 137664 118176 137670 118228
rect 51218 118040 51224 118092
rect 51276 118080 51282 118092
rect 56554 118080 56560 118092
rect 51276 118052 56560 118080
rect 51276 118040 51282 118052
rect 56554 118040 56560 118052
rect 56612 118040 56618 118092
rect 50574 117904 50580 117956
rect 50632 117944 50638 117956
rect 55542 117944 55548 117956
rect 50632 117916 55548 117944
rect 50632 117904 50638 117916
rect 55542 117904 55548 117916
rect 55600 117904 55606 117956
rect 97954 117904 97960 117956
rect 98012 117944 98018 117956
rect 101082 117944 101088 117956
rect 98012 117916 101088 117944
rect 98012 117904 98018 117916
rect 101082 117904 101088 117916
rect 101140 117904 101146 117956
rect 134846 117904 134852 117956
rect 134904 117944 134910 117956
rect 137422 117944 137428 117956
rect 134904 117916 137428 117944
rect 134904 117904 134910 117916
rect 137422 117904 137428 117916
rect 137480 117904 137486 117956
rect 182042 117904 182048 117956
rect 182100 117944 182106 117956
rect 185262 117944 185268 117956
rect 182100 117916 185268 117944
rect 182100 117904 182106 117916
rect 185262 117904 185268 117916
rect 185320 117904 185326 117956
rect 98138 117836 98144 117888
rect 98196 117876 98202 117888
rect 100990 117876 100996 117888
rect 98196 117848 100996 117876
rect 98196 117836 98202 117848
rect 100990 117836 100996 117848
rect 101048 117836 101054 117888
rect 182318 117836 182324 117888
rect 182376 117876 182382 117888
rect 185170 117876 185176 117888
rect 182376 117848 185176 117876
rect 182376 117836 182382 117848
rect 185170 117836 185176 117848
rect 185228 117836 185234 117888
rect 56738 117768 56744 117820
rect 56796 117808 56802 117820
rect 58210 117808 58216 117820
rect 56796 117780 58216 117808
rect 56796 117768 56802 117780
rect 58210 117768 58216 117780
rect 58268 117768 58274 117820
rect 92802 117768 92808 117820
rect 92860 117808 92866 117820
rect 98046 117808 98052 117820
rect 92860 117780 98052 117808
rect 92860 117768 92866 117780
rect 98046 117768 98052 117780
rect 98104 117768 98110 117820
rect 136962 117768 136968 117820
rect 137020 117808 137026 117820
rect 142574 117808 142580 117820
rect 137020 117780 142580 117808
rect 137020 117768 137026 117780
rect 142574 117768 142580 117780
rect 142632 117768 142638 117820
rect 56278 117700 56284 117752
rect 56336 117740 56342 117752
rect 58302 117740 58308 117752
rect 56336 117712 58308 117740
rect 56336 117700 56342 117712
rect 58302 117700 58308 117712
rect 58360 117700 58366 117752
rect 92710 117700 92716 117752
rect 92768 117740 92774 117752
rect 97862 117740 97868 117752
rect 92768 117712 97868 117740
rect 92768 117700 92774 117712
rect 97862 117700 97868 117712
rect 97920 117700 97926 117752
rect 137698 117700 137704 117752
rect 137756 117740 137762 117752
rect 143218 117740 143224 117752
rect 137756 117712 143224 117740
rect 137756 117700 137762 117712
rect 143218 117700 143224 117712
rect 143276 117700 143282 117752
rect 177718 117700 177724 117752
rect 177776 117740 177782 117752
rect 182134 117740 182140 117752
rect 177776 117712 182140 117740
rect 177776 117700 177782 117712
rect 182134 117700 182140 117712
rect 182192 117700 182198 117752
rect 177166 117428 177172 117480
rect 177224 117468 177230 117480
rect 182226 117468 182232 117480
rect 177224 117440 182232 117468
rect 177224 117428 177230 117440
rect 182226 117428 182232 117440
rect 182284 117428 182290 117480
rect 93998 116544 94004 116596
rect 94056 116584 94062 116596
rect 101082 116584 101088 116596
rect 94056 116556 101088 116584
rect 94056 116544 94062 116556
rect 101082 116544 101088 116556
rect 101140 116544 101146 116596
rect 178178 116544 178184 116596
rect 178236 116584 178242 116596
rect 185262 116584 185268 116596
rect 178236 116556 185268 116584
rect 178236 116544 178242 116556
rect 185262 116544 185268 116556
rect 185320 116544 185326 116596
rect 50022 116476 50028 116528
rect 50080 116516 50086 116528
rect 58210 116516 58216 116528
rect 50080 116488 58216 116516
rect 50080 116476 50086 116488
rect 58210 116476 58216 116488
rect 58268 116476 58274 116528
rect 92618 116476 92624 116528
rect 92676 116516 92682 116528
rect 100990 116516 100996 116528
rect 92676 116488 100996 116516
rect 92676 116476 92682 116488
rect 100990 116476 100996 116488
rect 101048 116476 101054 116528
rect 134846 116476 134852 116528
rect 134904 116516 134910 116528
rect 134904 116488 139676 116516
rect 134904 116476 134910 116488
rect 55542 116408 55548 116460
rect 55600 116448 55606 116460
rect 58302 116448 58308 116460
rect 55600 116420 58308 116448
rect 55600 116408 55606 116420
rect 58302 116408 58308 116420
rect 58360 116408 58366 116460
rect 92894 116408 92900 116460
rect 92952 116448 92958 116460
rect 101174 116448 101180 116460
rect 92952 116420 101180 116448
rect 92952 116408 92958 116420
rect 101174 116408 101180 116420
rect 101232 116408 101238 116460
rect 139648 116448 139676 116488
rect 176798 116476 176804 116528
rect 176856 116516 176862 116528
rect 185170 116516 185176 116528
rect 176856 116488 185176 116516
rect 176856 116476 176862 116488
rect 185170 116476 185176 116488
rect 185228 116476 185234 116528
rect 142758 116448 142764 116460
rect 139648 116420 142764 116448
rect 142758 116408 142764 116420
rect 142816 116408 142822 116460
rect 177074 116408 177080 116460
rect 177132 116448 177138 116460
rect 185354 116448 185360 116460
rect 177132 116420 185360 116448
rect 177132 116408 177138 116420
rect 185354 116408 185360 116420
rect 185412 116408 185418 116460
rect 56554 116340 56560 116392
rect 56612 116380 56618 116392
rect 58394 116380 58400 116392
rect 56612 116352 58400 116380
rect 56612 116340 56618 116352
rect 58394 116340 58400 116352
rect 58452 116340 58458 116392
rect 92802 116340 92808 116392
rect 92860 116380 92866 116392
rect 98138 116380 98144 116392
rect 92860 116352 98144 116380
rect 92860 116340 92866 116352
rect 98138 116340 98144 116352
rect 98196 116340 98202 116392
rect 137422 116340 137428 116392
rect 137480 116380 137486 116392
rect 142942 116380 142948 116392
rect 137480 116352 142948 116380
rect 137480 116340 137486 116352
rect 142942 116340 142948 116352
rect 143000 116340 143006 116392
rect 177718 116340 177724 116392
rect 177776 116380 177782 116392
rect 182042 116380 182048 116392
rect 177776 116352 182048 116380
rect 177776 116340 177782 116352
rect 182042 116340 182048 116352
rect 182100 116340 182106 116392
rect 92710 116272 92716 116324
rect 92768 116312 92774 116324
rect 97954 116312 97960 116324
rect 92768 116284 97960 116312
rect 92768 116272 92774 116284
rect 97954 116272 97960 116284
rect 98012 116272 98018 116324
rect 137606 116272 137612 116324
rect 137664 116312 137670 116324
rect 143586 116312 143592 116324
rect 137664 116284 143592 116312
rect 137664 116272 137670 116284
rect 143586 116272 143592 116284
rect 143644 116272 143650 116324
rect 177718 116068 177724 116120
rect 177776 116108 177782 116120
rect 182318 116108 182324 116120
rect 177776 116080 182324 116108
rect 177776 116068 177782 116080
rect 182318 116068 182324 116080
rect 182376 116068 182382 116120
rect 91238 115184 91244 115236
rect 91296 115224 91302 115236
rect 101082 115224 101088 115236
rect 91296 115196 101088 115224
rect 91296 115184 91302 115196
rect 101082 115184 101088 115196
rect 101140 115184 101146 115236
rect 175418 115184 175424 115236
rect 175476 115224 175482 115236
rect 185262 115224 185268 115236
rect 175476 115196 185268 115224
rect 175476 115184 175482 115196
rect 185262 115184 185268 115196
rect 185320 115184 185326 115236
rect 59314 115156 59320 115168
rect 59275 115128 59320 115156
rect 59314 115116 59320 115128
rect 59372 115116 59378 115168
rect 90594 115116 90600 115168
rect 90652 115156 90658 115168
rect 100990 115156 100996 115168
rect 90652 115128 100996 115156
rect 90652 115116 90658 115128
rect 100990 115116 100996 115128
rect 101048 115116 101054 115168
rect 174774 115116 174780 115168
rect 174832 115156 174838 115168
rect 185170 115156 185176 115168
rect 174832 115128 185176 115156
rect 174832 115116 174838 115128
rect 185170 115116 185176 115128
rect 185228 115116 185234 115168
rect 135398 113688 135404 113740
rect 135456 113728 135462 113740
rect 141562 113728 141568 113740
rect 135456 113700 141568 113728
rect 135456 113688 135462 113700
rect 141562 113688 141568 113700
rect 141620 113688 141626 113740
rect 18006 113280 18012 113332
rect 18064 113320 18070 113332
rect 64098 113320 64104 113332
rect 18064 113292 64104 113320
rect 18064 113280 18070 113292
rect 64098 113280 64104 113292
rect 64156 113280 64162 113332
rect 147266 113280 147272 113332
rect 147324 113320 147330 113332
rect 218382 113320 218388 113332
rect 147324 113292 218388 113320
rect 147324 113280 147330 113292
rect 218382 113280 218388 113292
rect 218440 113280 218446 113332
rect 51218 112736 51224 112788
rect 51276 112776 51282 112788
rect 54714 112776 54720 112788
rect 51276 112748 54720 112776
rect 51276 112736 51282 112748
rect 54714 112736 54720 112748
rect 54772 112736 54778 112788
rect 85718 112328 85724 112380
rect 85776 112368 85782 112380
rect 100990 112368 100996 112380
rect 85776 112340 100996 112368
rect 85776 112328 85782 112340
rect 100990 112328 100996 112340
rect 101048 112328 101054 112380
rect 169898 112328 169904 112380
rect 169956 112368 169962 112380
rect 185170 112368 185176 112380
rect 169956 112340 185176 112368
rect 169956 112328 169962 112340
rect 185170 112328 185176 112340
rect 185228 112328 185234 112380
rect 90410 112192 90416 112244
rect 90468 112232 90474 112244
rect 93354 112232 93360 112244
rect 90468 112204 93360 112232
rect 90468 112192 90474 112204
rect 93354 112192 93360 112204
rect 93412 112192 93418 112244
rect 82314 111580 82320 111632
rect 82372 111620 82378 111632
rect 85442 111620 85448 111632
rect 82372 111592 85448 111620
rect 82372 111580 82378 111592
rect 85442 111580 85448 111592
rect 85500 111580 85506 111632
rect 129970 111580 129976 111632
rect 130028 111620 130034 111632
rect 148094 111620 148100 111632
rect 130028 111592 148100 111620
rect 130028 111580 130034 111592
rect 148094 111580 148100 111592
rect 148152 111580 148158 111632
rect 83694 111512 83700 111564
rect 83752 111552 83758 111564
rect 87190 111552 87196 111564
rect 83752 111524 87196 111552
rect 83752 111512 83758 111524
rect 87190 111512 87196 111524
rect 87248 111512 87254 111564
rect 80934 111444 80940 111496
rect 80992 111484 80998 111496
rect 84062 111484 84068 111496
rect 80992 111456 84068 111484
rect 80992 111444 80998 111456
rect 84062 111444 84068 111456
rect 84120 111444 84126 111496
rect 79554 111104 79560 111156
rect 79612 111144 79618 111156
rect 82590 111144 82596 111156
rect 79612 111116 82596 111144
rect 79612 111104 79618 111116
rect 82590 111104 82596 111116
rect 82648 111104 82654 111156
rect 163826 111104 163832 111156
rect 163884 111144 163890 111156
rect 166586 111144 166592 111156
rect 163884 111116 166592 111144
rect 163884 111104 163890 111116
rect 166586 111104 166592 111116
rect 166644 111104 166650 111156
rect 167874 111104 167880 111156
rect 167932 111144 167938 111156
rect 170910 111144 170916 111156
rect 167932 111116 170916 111144
rect 167932 111104 167938 111116
rect 170910 111104 170916 111116
rect 170968 111104 170974 111156
rect 74034 111036 74040 111088
rect 74092 111076 74098 111088
rect 75506 111076 75512 111088
rect 74092 111048 75512 111076
rect 74092 111036 74098 111048
rect 75506 111036 75512 111048
rect 75564 111036 75570 111088
rect 77438 111036 77444 111088
rect 77496 111076 77502 111088
rect 79738 111076 79744 111088
rect 77496 111048 79744 111076
rect 77496 111036 77502 111048
rect 79738 111036 79744 111048
rect 79796 111036 79802 111088
rect 158858 111036 158864 111088
rect 158916 111076 158922 111088
rect 160882 111076 160888 111088
rect 158916 111048 160888 111076
rect 158916 111036 158922 111048
rect 160882 111036 160888 111048
rect 160940 111036 160946 111088
rect 166494 111036 166500 111088
rect 166552 111076 166558 111088
rect 169438 111076 169444 111088
rect 166552 111048 169444 111076
rect 166552 111036 166558 111048
rect 169438 111036 169444 111048
rect 169496 111036 169502 111088
rect 74678 110968 74684 111020
rect 74736 111008 74742 111020
rect 76886 111008 76892 111020
rect 74736 110980 76892 111008
rect 74736 110968 74742 110980
rect 76886 110968 76892 110980
rect 76944 110968 76950 111020
rect 79646 110968 79652 111020
rect 79704 111008 79710 111020
rect 81210 111008 81216 111020
rect 79704 110980 81216 111008
rect 79704 110968 79710 110980
rect 81210 110968 81216 110980
rect 81268 110968 81274 111020
rect 156834 110968 156840 111020
rect 156892 111008 156898 111020
rect 158030 111008 158036 111020
rect 156892 110980 158036 111008
rect 156892 110968 156898 110980
rect 158030 110968 158036 110980
rect 158088 110968 158094 111020
rect 158306 110968 158312 111020
rect 158364 111008 158370 111020
rect 159502 111008 159508 111020
rect 158364 110980 159508 111008
rect 158364 110968 158370 110980
rect 159502 110968 159508 110980
rect 159560 110968 159566 111020
rect 161618 110968 161624 111020
rect 161676 111008 161682 111020
rect 163734 111008 163740 111020
rect 161676 110980 163740 111008
rect 161676 110968 161682 110980
rect 163734 110968 163740 110980
rect 163792 110968 163798 111020
rect 165114 110968 165120 111020
rect 165172 111008 165178 111020
rect 168058 111008 168064 111020
rect 165172 110980 168064 111008
rect 165172 110968 165178 110980
rect 168058 110968 168064 110980
rect 168116 110968 168122 111020
rect 172658 110968 172664 111020
rect 172716 111008 172722 111020
rect 176154 111008 176160 111020
rect 172716 110980 176160 111008
rect 172716 110968 172722 110980
rect 176154 110968 176160 110980
rect 176212 110968 176218 111020
rect 61430 110900 61436 110952
rect 61488 110940 61494 110952
rect 108442 110940 108448 110952
rect 61488 110912 108448 110940
rect 61488 110900 61494 110912
rect 108442 110900 108448 110912
rect 108500 110900 108506 110952
rect 108994 110900 109000 110952
rect 109052 110940 109058 110952
rect 129970 110940 129976 110952
rect 109052 110912 129976 110940
rect 109052 110900 109058 110912
rect 129970 110900 129976 110912
rect 130028 110900 130034 110952
rect 137514 110900 137520 110952
rect 137572 110940 137578 110952
rect 145334 110940 145340 110952
rect 137572 110912 145340 110940
rect 137572 110900 137578 110912
rect 145334 110900 145340 110912
rect 145392 110900 145398 110952
rect 63270 110832 63276 110884
rect 63328 110872 63334 110884
rect 109546 110872 109552 110884
rect 63328 110844 109552 110872
rect 63328 110832 63334 110844
rect 109546 110832 109552 110844
rect 109604 110832 109610 110884
rect 113134 110492 113140 110544
rect 113192 110532 113198 110544
rect 114514 110532 114520 110544
rect 113192 110504 114520 110532
rect 113192 110492 113198 110504
rect 114514 110492 114520 110504
rect 114572 110492 114578 110544
rect 114606 110492 114612 110544
rect 114664 110532 114670 110544
rect 115618 110532 115624 110544
rect 114664 110504 115624 110532
rect 114664 110492 114670 110504
rect 115618 110492 115624 110504
rect 115676 110492 115682 110544
rect 115986 110492 115992 110544
rect 116044 110532 116050 110544
rect 117274 110532 117280 110544
rect 116044 110504 117280 110532
rect 116044 110492 116050 110504
rect 117274 110492 117280 110504
rect 117332 110492 117338 110544
rect 117458 110492 117464 110544
rect 117516 110532 117522 110544
rect 118838 110532 118844 110544
rect 117516 110504 118844 110532
rect 117516 110492 117522 110504
rect 118838 110492 118844 110504
rect 118896 110492 118902 110544
rect 99518 110424 99524 110476
rect 99576 110464 99582 110476
rect 107338 110464 107344 110476
rect 99576 110436 107344 110464
rect 99576 110424 99582 110436
rect 107338 110424 107344 110436
rect 107396 110424 107402 110476
rect 183606 110356 183612 110408
rect 183664 110396 183670 110408
rect 191610 110396 191616 110408
rect 183664 110368 191616 110396
rect 183664 110356 183670 110368
rect 191610 110356 191616 110368
rect 191668 110356 191674 110408
rect 99426 110288 99432 110340
rect 99484 110328 99490 110340
rect 106786 110328 106792 110340
rect 99484 110300 106792 110328
rect 99484 110288 99490 110300
rect 106786 110288 106792 110300
rect 106844 110288 106850 110340
rect 183698 110288 183704 110340
rect 183756 110328 183762 110340
rect 192162 110328 192168 110340
rect 183756 110300 192168 110328
rect 183756 110288 183762 110300
rect 192162 110288 192168 110300
rect 192220 110288 192226 110340
rect 208262 110288 208268 110340
rect 208320 110328 208326 110340
rect 213230 110328 213236 110340
rect 208320 110300 213236 110328
rect 208320 110288 208326 110300
rect 213230 110288 213236 110300
rect 213288 110288 213294 110340
rect 20214 110220 20220 110272
rect 20272 110260 20278 110272
rect 41742 110260 41748 110272
rect 20272 110232 41748 110260
rect 20272 110220 20278 110232
rect 41742 110220 41748 110232
rect 41800 110220 41806 110272
rect 53334 110220 53340 110272
rect 53392 110260 53398 110272
rect 61430 110260 61436 110272
rect 53392 110232 61436 110260
rect 53392 110220 53398 110232
rect 61430 110220 61436 110232
rect 61488 110220 61494 110272
rect 98782 110220 98788 110272
rect 98840 110260 98846 110272
rect 107890 110260 107896 110272
rect 98840 110232 107896 110260
rect 98840 110220 98846 110232
rect 107890 110220 107896 110232
rect 107948 110220 107954 110272
rect 108442 110220 108448 110272
rect 108500 110260 108506 110272
rect 133374 110260 133380 110272
rect 108500 110232 133380 110260
rect 108500 110220 108506 110232
rect 133374 110220 133380 110232
rect 133432 110260 133438 110272
rect 137514 110260 137520 110272
rect 133432 110232 137520 110260
rect 133432 110220 133438 110232
rect 137514 110220 137520 110232
rect 137572 110220 137578 110272
rect 183514 110220 183520 110272
rect 183572 110260 183578 110272
rect 191058 110260 191064 110272
rect 183572 110232 191064 110260
rect 183572 110220 183578 110232
rect 191058 110220 191064 110232
rect 191116 110220 191122 110272
rect 191978 110220 191984 110272
rect 192036 110260 192042 110272
rect 215530 110260 215536 110272
rect 192036 110232 215536 110260
rect 192036 110220 192042 110232
rect 215530 110220 215536 110232
rect 215588 110220 215594 110272
rect 113042 110152 113048 110204
rect 113100 110192 113106 110204
rect 113962 110192 113968 110204
rect 113100 110164 113968 110192
rect 113100 110152 113106 110164
rect 113962 110152 113968 110164
rect 114020 110152 114026 110204
rect 115710 110152 115716 110204
rect 115768 110192 115774 110204
rect 116722 110192 116728 110204
rect 115768 110164 116728 110192
rect 115768 110152 115774 110164
rect 116722 110152 116728 110164
rect 116780 110152 116786 110204
rect 115802 110016 115808 110068
rect 115860 110056 115866 110068
rect 118286 110056 118292 110068
rect 115860 110028 118292 110056
rect 115860 110016 115866 110028
rect 118286 110016 118292 110028
rect 118344 110016 118350 110068
rect 25918 109948 25924 110000
rect 25976 109988 25982 110000
rect 26286 109988 26292 110000
rect 25976 109960 26292 109988
rect 25976 109948 25982 109960
rect 26286 109948 26292 109960
rect 26344 109948 26350 110000
rect 29046 109948 29052 110000
rect 29104 109988 29110 110000
rect 30886 109988 30892 110000
rect 29104 109960 30892 109988
rect 29104 109948 29110 109960
rect 30886 109948 30892 109960
rect 30944 109948 30950 110000
rect 24906 109880 24912 109932
rect 24964 109920 24970 109932
rect 24964 109892 27528 109920
rect 24964 109880 24970 109892
rect 22882 109812 22888 109864
rect 22940 109852 22946 109864
rect 27298 109852 27304 109864
rect 22940 109824 27304 109852
rect 22940 109812 22946 109824
rect 27298 109812 27304 109824
rect 27356 109812 27362 109864
rect 27500 109852 27528 109892
rect 27666 109880 27672 109932
rect 27724 109920 27730 109932
rect 30058 109920 30064 109932
rect 27724 109892 30064 109920
rect 27724 109880 27730 109892
rect 30058 109880 30064 109892
rect 30116 109880 30122 109932
rect 28494 109852 28500 109864
rect 27500 109824 28500 109852
rect 28494 109812 28500 109824
rect 28552 109812 28558 109864
rect 99242 109812 99248 109864
rect 99300 109852 99306 109864
rect 106234 109852 106240 109864
rect 99300 109824 106240 109852
rect 99300 109812 99306 109824
rect 106234 109812 106240 109824
rect 106292 109812 106298 109864
rect 119758 109812 119764 109864
rect 119816 109852 119822 109864
rect 121598 109852 121604 109864
rect 119816 109824 121604 109852
rect 119816 109812 119822 109824
rect 121598 109812 121604 109824
rect 121656 109812 121662 109864
rect 183330 109812 183336 109864
rect 183388 109852 183394 109864
rect 190414 109852 190420 109864
rect 183388 109824 190420 109852
rect 183388 109812 183394 109824
rect 190414 109812 190420 109824
rect 190472 109812 190478 109864
rect 203754 109812 203760 109864
rect 203812 109852 203818 109864
rect 205318 109852 205324 109864
rect 203812 109824 205324 109852
rect 203812 109812 203818 109824
rect 205318 109812 205324 109824
rect 205376 109812 205382 109864
rect 23618 109744 23624 109796
rect 23676 109784 23682 109796
rect 27666 109784 27672 109796
rect 23676 109756 27672 109784
rect 23676 109744 23682 109756
rect 27666 109744 27672 109756
rect 27724 109744 27730 109796
rect 99150 109744 99156 109796
rect 99208 109784 99214 109796
rect 105682 109784 105688 109796
rect 99208 109756 105688 109784
rect 99208 109744 99214 109756
rect 105682 109744 105688 109756
rect 105740 109744 105746 109796
rect 118930 109744 118936 109796
rect 118988 109784 118994 109796
rect 119942 109784 119948 109796
rect 118988 109756 119948 109784
rect 118988 109744 118994 109756
rect 119942 109744 119948 109756
rect 120000 109744 120006 109796
rect 126658 109744 126664 109796
rect 126716 109784 126722 109796
rect 129326 109784 129332 109796
rect 126716 109756 129332 109784
rect 126716 109744 126722 109756
rect 129326 109744 129332 109756
rect 129384 109744 129390 109796
rect 183238 109744 183244 109796
rect 183296 109784 183302 109796
rect 189862 109784 189868 109796
rect 183296 109756 189868 109784
rect 183296 109744 183302 109756
rect 189862 109744 189868 109756
rect 189920 109744 189926 109796
rect 21502 109676 21508 109728
rect 21560 109716 21566 109728
rect 26470 109716 26476 109728
rect 21560 109688 26476 109716
rect 21560 109676 21566 109688
rect 26470 109676 26476 109688
rect 26528 109676 26534 109728
rect 42938 109676 42944 109728
rect 42996 109716 43002 109728
rect 47446 109716 47452 109728
rect 42996 109688 47452 109716
rect 42996 109676 43002 109688
rect 47446 109676 47452 109688
rect 47504 109676 47510 109728
rect 99058 109676 99064 109728
rect 99116 109716 99122 109728
rect 104578 109716 104584 109728
rect 99116 109688 104584 109716
rect 99116 109676 99122 109688
rect 104578 109676 104584 109688
rect 104636 109676 104642 109728
rect 115894 109676 115900 109728
rect 115952 109716 115958 109728
rect 117826 109716 117832 109728
rect 115952 109688 117832 109716
rect 115952 109676 115958 109688
rect 117826 109676 117832 109688
rect 117884 109676 117890 109728
rect 119574 109676 119580 109728
rect 119632 109716 119638 109728
rect 121046 109716 121052 109728
rect 119632 109688 121052 109716
rect 119632 109676 119638 109688
rect 121046 109676 121052 109688
rect 121104 109676 121110 109728
rect 183146 109676 183152 109728
rect 183204 109716 183210 109728
rect 188758 109716 188764 109728
rect 183204 109688 188764 109716
rect 183204 109676 183210 109688
rect 188758 109676 188764 109688
rect 188816 109676 188822 109728
rect 205318 109676 205324 109728
rect 205376 109716 205382 109728
rect 206422 109716 206428 109728
rect 205376 109688 206428 109716
rect 205376 109676 205382 109688
rect 206422 109676 206428 109688
rect 206480 109676 206486 109728
rect 208170 109676 208176 109728
rect 208228 109716 208234 109728
rect 212126 109716 212132 109728
rect 208228 109688 212132 109716
rect 208228 109676 208234 109688
rect 212126 109676 212132 109688
rect 212184 109676 212190 109728
rect 22238 109608 22244 109660
rect 22296 109648 22302 109660
rect 26562 109648 26568 109660
rect 22296 109620 26568 109648
rect 22296 109608 22302 109620
rect 26562 109608 26568 109620
rect 26620 109608 26626 109660
rect 27022 109608 27028 109660
rect 27080 109648 27086 109660
rect 29690 109648 29696 109660
rect 27080 109620 29696 109648
rect 27080 109608 27086 109620
rect 29690 109608 29696 109620
rect 29748 109608 29754 109660
rect 38246 109608 38252 109660
rect 38304 109648 38310 109660
rect 39994 109648 40000 109660
rect 38304 109620 40000 109648
rect 38304 109608 38310 109620
rect 39994 109608 40000 109620
rect 40052 109608 40058 109660
rect 45054 109608 45060 109660
rect 45112 109648 45118 109660
rect 46802 109648 46808 109660
rect 45112 109620 46808 109648
rect 45112 109608 45118 109620
rect 46802 109608 46808 109620
rect 46860 109608 46866 109660
rect 98966 109608 98972 109660
rect 99024 109648 99030 109660
rect 104118 109648 104124 109660
rect 99024 109620 104124 109648
rect 99024 109608 99030 109620
rect 104118 109608 104124 109620
rect 104176 109608 104182 109660
rect 119942 109608 119948 109660
rect 120000 109648 120006 109660
rect 122150 109648 122156 109660
rect 120000 109620 122156 109648
rect 120000 109608 120006 109620
rect 122150 109608 122156 109620
rect 122208 109608 122214 109660
rect 126566 109608 126572 109660
rect 126624 109648 126630 109660
rect 128774 109648 128780 109660
rect 126624 109620 128780 109648
rect 126624 109608 126630 109620
rect 128774 109608 128780 109620
rect 128832 109608 128838 109660
rect 129326 109608 129332 109660
rect 129384 109648 129390 109660
rect 130982 109648 130988 109660
rect 129384 109620 130988 109648
rect 129384 109608 129390 109620
rect 130982 109608 130988 109620
rect 131040 109608 131046 109660
rect 183054 109608 183060 109660
rect 183112 109648 183118 109660
rect 188206 109648 188212 109660
rect 183112 109620 188212 109648
rect 183112 109608 183118 109620
rect 188206 109608 188212 109620
rect 188264 109608 188270 109660
rect 201454 109608 201460 109660
rect 201512 109648 201518 109660
rect 203018 109648 203024 109660
rect 201512 109620 203024 109648
rect 201512 109608 201518 109620
rect 203018 109608 203024 109620
rect 203076 109608 203082 109660
rect 205134 109608 205140 109660
rect 205192 109648 205198 109660
rect 205870 109648 205876 109660
rect 205192 109620 205876 109648
rect 205192 109608 205198 109620
rect 205870 109608 205876 109620
rect 205928 109608 205934 109660
rect 208538 109608 208544 109660
rect 208596 109648 208602 109660
rect 212678 109648 212684 109660
rect 208596 109620 212684 109648
rect 208596 109608 208602 109620
rect 212678 109608 212684 109620
rect 212736 109608 212742 109660
rect 213506 109608 213512 109660
rect 213564 109648 213570 109660
rect 214978 109648 214984 109660
rect 213564 109620 214984 109648
rect 213564 109608 213570 109620
rect 214978 109608 214984 109620
rect 215036 109608 215042 109660
rect 20858 109540 20864 109592
rect 20916 109580 20922 109592
rect 22974 109580 22980 109592
rect 20916 109552 22980 109580
rect 20916 109540 20922 109552
rect 22974 109540 22980 109552
rect 23032 109540 23038 109592
rect 24262 109540 24268 109592
rect 24320 109580 24326 109592
rect 28126 109580 28132 109592
rect 24320 109552 28132 109580
rect 24320 109540 24326 109552
rect 28126 109540 28132 109552
rect 28184 109540 28190 109592
rect 28310 109540 28316 109592
rect 28368 109580 28374 109592
rect 29138 109580 29144 109592
rect 28368 109552 29144 109580
rect 28368 109540 28374 109552
rect 29138 109540 29144 109552
rect 29196 109540 29202 109592
rect 31070 109540 31076 109592
rect 31128 109580 31134 109592
rect 31806 109580 31812 109592
rect 31128 109552 31812 109580
rect 31128 109540 31134 109552
rect 31806 109540 31812 109552
rect 31864 109540 31870 109592
rect 38154 109540 38160 109592
rect 38212 109580 38218 109592
rect 39258 109580 39264 109592
rect 38212 109552 39264 109580
rect 38212 109540 38218 109552
rect 39258 109540 39264 109552
rect 39316 109540 39322 109592
rect 45146 109540 45152 109592
rect 45204 109580 45210 109592
rect 46066 109580 46072 109592
rect 45204 109552 46072 109580
rect 45204 109540 45210 109552
rect 46066 109540 46072 109552
rect 46124 109540 46130 109592
rect 99334 109540 99340 109592
rect 99392 109580 99398 109592
rect 105130 109580 105136 109592
rect 99392 109552 105136 109580
rect 99392 109540 99398 109552
rect 105130 109540 105136 109552
rect 105188 109540 105194 109592
rect 119850 109540 119856 109592
rect 119908 109580 119914 109592
rect 120494 109580 120500 109592
rect 119908 109552 120500 109580
rect 119908 109540 119914 109552
rect 120494 109540 120500 109552
rect 120552 109540 120558 109592
rect 120954 109540 120960 109592
rect 121012 109580 121018 109592
rect 122702 109580 122708 109592
rect 121012 109552 122708 109580
rect 121012 109540 121018 109552
rect 122702 109540 122708 109552
rect 122760 109540 122766 109592
rect 126474 109540 126480 109592
rect 126532 109580 126538 109592
rect 128222 109580 128228 109592
rect 126532 109552 128228 109580
rect 126532 109540 126538 109552
rect 128222 109540 128228 109552
rect 128280 109540 128286 109592
rect 129234 109540 129240 109592
rect 129292 109580 129298 109592
rect 130430 109580 130436 109592
rect 129292 109552 130436 109580
rect 129292 109540 129298 109552
rect 130430 109540 130436 109552
rect 130488 109540 130494 109592
rect 183422 109540 183428 109592
rect 183480 109580 183486 109592
rect 189310 109580 189316 109592
rect 183480 109552 189316 109580
rect 183480 109540 183486 109552
rect 189310 109540 189316 109552
rect 189368 109540 189374 109592
rect 193910 109540 193916 109592
rect 193968 109580 193974 109592
rect 194738 109580 194744 109592
rect 193968 109552 194744 109580
rect 193968 109540 193974 109552
rect 194738 109540 194744 109552
rect 194796 109540 194802 109592
rect 201638 109540 201644 109592
rect 201696 109580 201702 109592
rect 202466 109580 202472 109592
rect 201696 109552 202472 109580
rect 201696 109540 201702 109552
rect 202466 109540 202472 109552
rect 202524 109540 202530 109592
rect 203846 109540 203852 109592
rect 203904 109580 203910 109592
rect 204674 109580 204680 109592
rect 203904 109552 204680 109580
rect 203904 109540 203910 109552
rect 204674 109540 204680 109552
rect 204732 109540 204738 109592
rect 205410 109540 205416 109592
rect 205468 109580 205474 109592
rect 206974 109580 206980 109592
rect 205468 109552 206980 109580
rect 205468 109540 205474 109552
rect 206974 109540 206980 109552
rect 207032 109540 207038 109592
rect 208354 109540 208360 109592
rect 208412 109580 208418 109592
rect 211574 109580 211580 109592
rect 208412 109552 211580 109580
rect 208412 109540 208418 109552
rect 211574 109540 211580 109552
rect 211632 109540 211638 109592
rect 213414 109540 213420 109592
rect 213472 109580 213478 109592
rect 214426 109580 214432 109592
rect 213472 109552 214432 109580
rect 213472 109540 213478 109552
rect 214426 109540 214432 109552
rect 214484 109540 214490 109592
rect 59314 108180 59320 108232
rect 59372 108180 59378 108232
rect 59332 108152 59360 108180
rect 59406 108152 59412 108164
rect 59332 108124 59412 108152
rect 59406 108112 59412 108124
rect 59464 108112 59470 108164
rect 208630 107500 208636 107552
rect 208688 107540 208694 107552
rect 209550 107540 209556 107552
rect 208688 107512 209556 107540
rect 208688 107500 208694 107512
rect 209550 107500 209556 107512
rect 209608 107500 209614 107552
rect 210010 107500 210016 107552
rect 210068 107540 210074 107552
rect 210654 107540 210660 107552
rect 210068 107512 210660 107540
rect 210068 107500 210074 107512
rect 210654 107500 210660 107512
rect 210712 107500 210718 107552
rect 194922 102672 194928 102724
rect 194980 102712 194986 102724
rect 195106 102712 195112 102724
rect 194980 102684 195112 102712
rect 194980 102672 194986 102684
rect 195106 102672 195112 102684
rect 195164 102672 195170 102724
rect 199062 102672 199068 102724
rect 199120 102672 199126 102724
rect 30242 102604 30248 102656
rect 30300 102644 30306 102656
rect 31254 102644 31260 102656
rect 30300 102616 31260 102644
rect 30300 102604 30306 102616
rect 31254 102604 31260 102616
rect 31312 102604 31318 102656
rect 31990 102604 31996 102656
rect 32048 102644 32054 102656
rect 32818 102644 32824 102656
rect 32048 102616 32824 102644
rect 32048 102604 32054 102616
rect 32818 102604 32824 102616
rect 32876 102604 32882 102656
rect 33462 102604 33468 102656
rect 33520 102644 33526 102656
rect 34106 102644 34112 102656
rect 33520 102616 34112 102644
rect 33520 102604 33526 102616
rect 34106 102604 34112 102616
rect 34164 102604 34170 102656
rect 35118 102604 35124 102656
rect 35176 102644 35182 102656
rect 35486 102644 35492 102656
rect 35176 102616 35492 102644
rect 35176 102604 35182 102616
rect 35486 102604 35492 102616
rect 35544 102604 35550 102656
rect 35670 102604 35676 102656
rect 35728 102644 35734 102656
rect 36590 102644 36596 102656
rect 35728 102616 36596 102644
rect 35728 102604 35734 102616
rect 36590 102604 36596 102616
rect 36648 102604 36654 102656
rect 37694 102604 37700 102656
rect 37752 102644 37758 102656
rect 40270 102644 40276 102656
rect 37752 102616 40276 102644
rect 37752 102604 37758 102616
rect 40270 102604 40276 102616
rect 40328 102604 40334 102656
rect 54714 102604 54720 102656
rect 54772 102644 54778 102656
rect 56462 102644 56468 102656
rect 54772 102616 56468 102644
rect 54772 102604 54778 102616
rect 56462 102604 56468 102616
rect 56520 102604 56526 102656
rect 111294 102604 111300 102656
rect 111352 102644 111358 102656
rect 111754 102644 111760 102656
rect 111352 102616 111760 102644
rect 111352 102604 111358 102616
rect 111754 102604 111760 102616
rect 111812 102604 111818 102656
rect 112490 102604 112496 102656
rect 112548 102644 112554 102656
rect 113318 102644 113324 102656
rect 112548 102616 113324 102644
rect 112548 102604 112554 102616
rect 113318 102604 113324 102616
rect 113376 102604 113382 102656
rect 113686 102604 113692 102656
rect 113744 102644 113750 102656
rect 114698 102644 114704 102656
rect 113744 102616 114704 102644
rect 113744 102604 113750 102616
rect 114698 102604 114704 102616
rect 114756 102604 114762 102656
rect 115618 102604 115624 102656
rect 115676 102644 115682 102656
rect 115894 102644 115900 102656
rect 115676 102616 115900 102644
rect 115676 102604 115682 102616
rect 115894 102604 115900 102616
rect 115952 102604 115958 102656
rect 193266 102604 193272 102656
rect 193324 102644 193330 102656
rect 194094 102644 194100 102656
rect 193324 102616 194100 102644
rect 193324 102604 193330 102616
rect 194094 102604 194100 102616
rect 194152 102604 194158 102656
rect 196302 102604 196308 102656
rect 196360 102644 196366 102656
rect 196854 102644 196860 102656
rect 196360 102616 196860 102644
rect 196360 102604 196366 102616
rect 196854 102604 196860 102616
rect 196912 102604 196918 102656
rect 198418 102604 198424 102656
rect 198476 102644 198482 102656
rect 199080 102644 199108 102672
rect 198476 102616 199108 102644
rect 198476 102604 198482 102616
rect 199614 102604 199620 102656
rect 199672 102644 199678 102656
rect 200350 102644 200356 102656
rect 199672 102616 200356 102644
rect 199672 102604 199678 102616
rect 200350 102604 200356 102616
rect 200408 102604 200414 102656
rect 200810 102604 200816 102656
rect 200868 102644 200874 102656
rect 201638 102644 201644 102656
rect 200868 102616 201644 102644
rect 200868 102604 200874 102616
rect 201638 102604 201644 102616
rect 201696 102604 201702 102656
rect 202834 102604 202840 102656
rect 202892 102644 202898 102656
rect 203754 102644 203760 102656
rect 202892 102616 203760 102644
rect 202892 102604 202898 102616
rect 203754 102604 203760 102616
rect 203812 102604 203818 102656
rect 204858 102604 204864 102656
rect 204916 102644 204922 102656
rect 207342 102644 207348 102656
rect 204916 102616 207348 102644
rect 204916 102604 204922 102616
rect 207342 102604 207348 102616
rect 207400 102604 207406 102656
rect 32082 102536 32088 102588
rect 32140 102576 32146 102588
rect 33278 102576 33284 102588
rect 32140 102548 33284 102576
rect 32140 102536 32146 102548
rect 33278 102536 33284 102548
rect 33336 102536 33342 102588
rect 36498 102536 36504 102588
rect 36556 102576 36562 102588
rect 38062 102576 38068 102588
rect 36556 102548 38068 102576
rect 36556 102536 36562 102548
rect 38062 102536 38068 102548
rect 38120 102536 38126 102588
rect 111662 102536 111668 102588
rect 111720 102576 111726 102588
rect 112306 102576 112312 102588
rect 111720 102548 112312 102576
rect 111720 102536 111726 102548
rect 112306 102536 112312 102548
rect 112364 102536 112370 102588
rect 114054 102536 114060 102588
rect 114112 102576 114118 102588
rect 114606 102576 114612 102588
rect 114112 102548 114612 102576
rect 114112 102536 114118 102548
rect 114606 102536 114612 102548
rect 114664 102536 114670 102588
rect 114882 102536 114888 102588
rect 114940 102576 114946 102588
rect 115710 102576 115716 102588
rect 114940 102548 115716 102576
rect 114940 102536 114946 102548
rect 115710 102536 115716 102548
rect 115768 102536 115774 102588
rect 199246 102536 199252 102588
rect 199304 102576 199310 102588
rect 199706 102576 199712 102588
rect 199304 102548 199712 102576
rect 199304 102536 199310 102548
rect 199706 102536 199712 102548
rect 199764 102536 199770 102588
rect 202466 102536 202472 102588
rect 202524 102576 202530 102588
rect 203846 102576 203852 102588
rect 202524 102548 203852 102576
rect 202524 102536 202530 102548
rect 203846 102536 203852 102548
rect 203904 102536 203910 102588
rect 204030 102536 204036 102588
rect 204088 102576 204094 102588
rect 205410 102576 205416 102588
rect 204088 102548 205416 102576
rect 204088 102536 204094 102548
rect 205410 102536 205416 102548
rect 205468 102536 205474 102588
rect 115250 102468 115256 102520
rect 115308 102508 115314 102520
rect 115986 102508 115992 102520
rect 115308 102480 115992 102508
rect 115308 102468 115314 102480
rect 115986 102468 115992 102480
rect 116044 102468 116050 102520
rect 120494 102468 120500 102520
rect 120552 102508 120558 102520
rect 124358 102508 124364 102520
rect 120552 102480 124364 102508
rect 120552 102468 120558 102480
rect 124358 102468 124364 102480
rect 124416 102468 124422 102520
rect 201638 102468 201644 102520
rect 201696 102508 201702 102520
rect 203110 102508 203116 102520
rect 201696 102480 203116 102508
rect 201696 102468 201702 102480
rect 203110 102468 203116 102480
rect 203168 102468 203174 102520
rect 203294 102468 203300 102520
rect 203352 102508 203358 102520
rect 205134 102508 205140 102520
rect 203352 102480 205140 102508
rect 203352 102468 203358 102480
rect 205134 102468 205140 102480
rect 205192 102468 205198 102520
rect 22974 102400 22980 102452
rect 23032 102440 23038 102452
rect 26102 102440 26108 102452
rect 23032 102412 26108 102440
rect 23032 102400 23038 102412
rect 26102 102400 26108 102412
rect 26160 102400 26166 102452
rect 36866 102400 36872 102452
rect 36924 102440 36930 102452
rect 38154 102440 38160 102452
rect 36924 102412 38160 102440
rect 36924 102400 36930 102412
rect 38154 102400 38160 102412
rect 38212 102400 38218 102452
rect 50942 102400 50948 102452
rect 51000 102440 51006 102452
rect 57566 102440 57572 102452
rect 51000 102412 57572 102440
rect 51000 102400 51006 102412
rect 57566 102400 57572 102412
rect 57624 102400 57630 102452
rect 93354 102400 93360 102452
rect 93412 102440 93418 102452
rect 94182 102440 94188 102452
rect 93412 102412 94188 102440
rect 93412 102400 93418 102412
rect 94182 102400 94188 102412
rect 94240 102400 94246 102452
rect 120034 102400 120040 102452
rect 120092 102440 120098 102452
rect 123806 102440 123812 102452
rect 120092 102412 123812 102440
rect 120092 102400 120098 102412
rect 123806 102400 123812 102412
rect 123864 102400 123870 102452
rect 205226 102400 205232 102452
rect 205284 102440 205290 102452
rect 208814 102440 208820 102452
rect 205284 102412 208820 102440
rect 205284 102400 205290 102412
rect 208814 102400 208820 102412
rect 208872 102400 208878 102452
rect 38062 102332 38068 102384
rect 38120 102372 38126 102384
rect 40822 102372 40828 102384
rect 38120 102344 40828 102372
rect 38120 102332 38126 102344
rect 40822 102332 40828 102344
rect 40880 102332 40886 102384
rect 51126 102332 51132 102384
rect 51184 102372 51190 102384
rect 59774 102372 59780 102384
rect 51184 102344 59780 102372
rect 51184 102332 51190 102344
rect 59774 102332 59780 102344
rect 59832 102332 59838 102384
rect 119666 102332 119672 102384
rect 119724 102372 119730 102384
rect 123254 102372 123260 102384
rect 119724 102344 123260 102372
rect 119724 102332 119730 102344
rect 123254 102332 123260 102344
rect 123312 102332 123318 102384
rect 135122 102332 135128 102384
rect 135180 102372 135186 102384
rect 143770 102372 143776 102384
rect 135180 102344 143776 102372
rect 135180 102332 135186 102344
rect 143770 102332 143776 102344
rect 143828 102332 143834 102384
rect 206422 102332 206428 102384
rect 206480 102372 206486 102384
rect 210102 102372 210108 102384
rect 206480 102344 210108 102372
rect 206480 102332 206486 102344
rect 210102 102332 210108 102344
rect 210160 102332 210166 102384
rect 143678 102264 143684 102316
rect 143736 102304 143742 102316
rect 167138 102304 167144 102316
rect 143736 102276 167144 102304
rect 143736 102264 143742 102276
rect 167138 102264 167144 102276
rect 167196 102264 167202 102316
rect 50850 102196 50856 102248
rect 50908 102236 50914 102248
rect 60878 102236 60884 102248
rect 50908 102208 60884 102236
rect 50908 102196 50914 102208
rect 60878 102196 60884 102208
rect 60936 102196 60942 102248
rect 114422 102196 114428 102248
rect 114480 102236 114486 102248
rect 116170 102236 116176 102248
rect 114480 102208 116176 102236
rect 114480 102196 114486 102208
rect 116170 102196 116176 102208
rect 116228 102196 116234 102248
rect 122426 102196 122432 102248
rect 122484 102236 122490 102248
rect 127118 102236 127124 102248
rect 122484 102208 127124 102236
rect 122484 102196 122490 102208
rect 127118 102196 127124 102208
rect 127176 102196 127182 102248
rect 135030 102196 135036 102248
rect 135088 102236 135094 102248
rect 144874 102236 144880 102248
rect 135088 102208 144880 102236
rect 135088 102196 135094 102208
rect 144874 102196 144880 102208
rect 144932 102196 144938 102248
rect 208814 102196 208820 102248
rect 208872 102236 208878 102248
rect 212862 102236 212868 102248
rect 208872 102208 212868 102236
rect 208872 102196 208878 102208
rect 212862 102196 212868 102208
rect 212920 102196 212926 102248
rect 50666 102128 50672 102180
rect 50724 102168 50730 102180
rect 61982 102168 61988 102180
rect 50724 102140 61988 102168
rect 50724 102128 50730 102140
rect 61982 102128 61988 102140
rect 62040 102128 62046 102180
rect 121690 102128 121696 102180
rect 121748 102168 121754 102180
rect 126014 102168 126020 102180
rect 121748 102140 126020 102168
rect 121748 102128 121754 102140
rect 126014 102128 126020 102140
rect 126072 102128 126078 102180
rect 134846 102128 134852 102180
rect 134904 102168 134910 102180
rect 145978 102168 145984 102180
rect 134904 102140 145984 102168
rect 134904 102128 134910 102140
rect 145978 102128 145984 102140
rect 146036 102128 146042 102180
rect 203662 102128 203668 102180
rect 203720 102168 203726 102180
rect 205318 102168 205324 102180
rect 203720 102140 205324 102168
rect 203720 102128 203726 102140
rect 205318 102128 205324 102140
rect 205376 102128 205382 102180
rect 50758 102060 50764 102112
rect 50816 102100 50822 102112
rect 63086 102100 63092 102112
rect 50816 102072 63092 102100
rect 50816 102060 50822 102072
rect 63086 102060 63092 102072
rect 63144 102060 63150 102112
rect 88662 102060 88668 102112
rect 88720 102100 88726 102112
rect 102002 102100 102008 102112
rect 88720 102072 102008 102100
rect 88720 102060 88726 102072
rect 102002 102060 102008 102072
rect 102060 102060 102066 102112
rect 122886 102060 122892 102112
rect 122944 102100 122950 102112
rect 127670 102100 127676 102112
rect 122944 102072 127676 102100
rect 122944 102060 122950 102072
rect 127670 102060 127676 102072
rect 127728 102060 127734 102112
rect 134754 102060 134760 102112
rect 134812 102100 134818 102112
rect 147082 102100 147088 102112
rect 134812 102072 147088 102100
rect 134812 102060 134818 102072
rect 147082 102060 147088 102072
rect 147140 102060 147146 102112
rect 172658 102060 172664 102112
rect 172716 102100 172722 102112
rect 185998 102100 186004 102112
rect 172716 102072 186004 102100
rect 172716 102060 172722 102072
rect 185998 102060 186004 102072
rect 186056 102060 186062 102112
rect 209274 102060 209280 102112
rect 209332 102100 209338 102112
rect 213414 102100 213420 102112
rect 209332 102072 213420 102100
rect 209332 102060 209338 102072
rect 213414 102060 213420 102072
rect 213472 102060 213478 102112
rect 26286 101992 26292 102044
rect 26344 102032 26350 102044
rect 28862 102032 28868 102044
rect 26344 102004 28868 102032
rect 26344 101992 26350 102004
rect 28862 101992 28868 102004
rect 28920 101992 28926 102044
rect 29138 101992 29144 102044
rect 29196 102032 29202 102044
rect 30426 102032 30432 102044
rect 29196 102004 30432 102032
rect 29196 101992 29202 102004
rect 30426 101992 30432 102004
rect 30484 101992 30490 102044
rect 37234 101992 37240 102044
rect 37292 102032 37298 102044
rect 38246 102032 38252 102044
rect 37292 102004 38252 102032
rect 37292 101992 37298 102004
rect 38246 101992 38252 102004
rect 38304 101992 38310 102044
rect 41650 101992 41656 102044
rect 41708 102032 41714 102044
rect 42938 102032 42944 102044
rect 41708 102004 42944 102032
rect 41708 101992 41714 102004
rect 42938 101992 42944 102004
rect 42996 101992 43002 102044
rect 50574 101992 50580 102044
rect 50632 102032 50638 102044
rect 64190 102032 64196 102044
rect 50632 102004 64196 102032
rect 50632 101992 50638 102004
rect 64190 101992 64196 102004
rect 64248 101992 64254 102044
rect 87558 101992 87564 102044
rect 87616 102032 87622 102044
rect 101634 102032 101640 102044
rect 87616 102004 101640 102032
rect 87616 101992 87622 102004
rect 101634 101992 101640 102004
rect 101692 101992 101698 102044
rect 122058 101992 122064 102044
rect 122116 102032 122122 102044
rect 126106 102032 126112 102044
rect 122116 102004 126112 102032
rect 122116 101992 122122 102004
rect 126106 101992 126112 102004
rect 126164 101992 126170 102044
rect 134938 101992 134944 102044
rect 134996 102032 135002 102044
rect 148186 102032 148192 102044
rect 134996 102004 148192 102032
rect 134996 101992 135002 102004
rect 148186 101992 148192 102004
rect 148244 101992 148250 102044
rect 161526 101992 161532 102044
rect 161584 102032 161590 102044
rect 164470 102032 164476 102044
rect 161584 102004 164476 102032
rect 161584 101992 161590 102004
rect 164470 101992 164476 102004
rect 164528 101992 164534 102044
rect 171554 101992 171560 102044
rect 171612 102032 171618 102044
rect 185814 102032 185820 102044
rect 171612 102004 185820 102032
rect 171612 101992 171618 102004
rect 185814 101992 185820 102004
rect 185872 101992 185878 102044
rect 202098 101992 202104 102044
rect 202156 102032 202162 102044
rect 203202 102032 203208 102044
rect 202156 102004 203208 102032
rect 202156 101992 202162 102004
rect 203202 101992 203208 102004
rect 203260 101992 203266 102044
rect 50482 101924 50488 101976
rect 50540 101964 50546 101976
rect 58670 101964 58676 101976
rect 50540 101936 58676 101964
rect 50540 101924 50546 101936
rect 58670 101924 58676 101936
rect 58728 101924 58734 101976
rect 59406 101924 59412 101976
rect 59464 101964 59470 101976
rect 83142 101964 83148 101976
rect 59464 101936 83148 101964
rect 59464 101924 59470 101936
rect 83142 101924 83148 101936
rect 83200 101924 83206 101976
rect 86454 101924 86460 101976
rect 86512 101964 86518 101976
rect 101818 101964 101824 101976
rect 86512 101936 101824 101964
rect 86512 101924 86518 101936
rect 101818 101924 101824 101936
rect 101876 101924 101882 101976
rect 112030 101924 112036 101976
rect 112088 101964 112094 101976
rect 112858 101964 112864 101976
rect 112088 101936 112864 101964
rect 112088 101924 112094 101936
rect 112858 101924 112864 101936
rect 112916 101924 112922 101976
rect 121230 101924 121236 101976
rect 121288 101964 121294 101976
rect 125462 101964 125468 101976
rect 121288 101936 125468 101964
rect 121288 101924 121294 101936
rect 125462 101924 125468 101936
rect 125520 101924 125526 101976
rect 135306 101924 135312 101976
rect 135364 101964 135370 101976
rect 142666 101964 142672 101976
rect 135364 101936 142672 101964
rect 135364 101924 135370 101936
rect 142666 101924 142672 101936
rect 142724 101924 142730 101976
rect 170450 101924 170456 101976
rect 170508 101964 170514 101976
rect 186182 101964 186188 101976
rect 170508 101936 186188 101964
rect 170508 101924 170514 101936
rect 186182 101924 186188 101936
rect 186240 101924 186246 101976
rect 209642 101924 209648 101976
rect 209700 101964 209706 101976
rect 213506 101964 213512 101976
rect 209700 101936 213512 101964
rect 209700 101924 209706 101936
rect 213506 101924 213512 101936
rect 213564 101924 213570 101976
rect 40086 101856 40092 101908
rect 40144 101896 40150 101908
rect 44410 101896 44416 101908
rect 40144 101868 44416 101896
rect 40144 101856 40150 101868
rect 44410 101856 44416 101868
rect 44468 101856 44474 101908
rect 200442 101856 200448 101908
rect 200500 101896 200506 101908
rect 201546 101896 201552 101908
rect 200500 101868 201552 101896
rect 200500 101856 200506 101868
rect 201546 101856 201552 101868
rect 201604 101856 201610 101908
rect 30518 101788 30524 101840
rect 30576 101828 30582 101840
rect 31622 101828 31628 101840
rect 30576 101800 31628 101828
rect 30576 101788 30582 101800
rect 31622 101788 31628 101800
rect 31680 101788 31686 101840
rect 40822 101788 40828 101840
rect 40880 101828 40886 101840
rect 45146 101828 45152 101840
rect 40880 101800 45152 101828
rect 40880 101788 40886 101800
rect 45146 101788 45152 101800
rect 45204 101788 45210 101840
rect 116446 101788 116452 101840
rect 116504 101828 116510 101840
rect 117458 101828 117464 101840
rect 116504 101800 117464 101828
rect 116504 101788 116510 101800
rect 117458 101788 117464 101800
rect 117516 101788 117522 101840
rect 124450 101788 124456 101840
rect 124508 101828 124514 101840
rect 129878 101828 129884 101840
rect 124508 101800 129884 101828
rect 124508 101788 124514 101800
rect 129878 101788 129884 101800
rect 129936 101788 129942 101840
rect 206882 101788 206888 101840
rect 206940 101828 206946 101840
rect 210010 101828 210016 101840
rect 206940 101800 210016 101828
rect 206940 101788 206946 101800
rect 210010 101788 210016 101800
rect 210068 101788 210074 101840
rect 26378 101720 26384 101772
rect 26436 101760 26442 101772
rect 29230 101760 29236 101772
rect 26436 101732 29236 101760
rect 26436 101720 26442 101732
rect 29230 101720 29236 101732
rect 29288 101720 29294 101772
rect 39626 101720 39632 101772
rect 39684 101760 39690 101772
rect 43582 101760 43588 101772
rect 39684 101732 43588 101760
rect 39684 101720 39690 101732
rect 43582 101720 43588 101732
rect 43640 101720 43646 101772
rect 120862 101720 120868 101772
rect 120920 101760 120926 101772
rect 124910 101760 124916 101772
rect 120920 101732 124916 101760
rect 120920 101720 120926 101732
rect 124910 101720 124916 101732
rect 124968 101720 124974 101772
rect 35302 101652 35308 101704
rect 35360 101692 35366 101704
rect 36130 101692 36136 101704
rect 35360 101664 36136 101692
rect 35360 101652 35366 101664
rect 36130 101652 36136 101664
rect 36188 101652 36194 101704
rect 39258 101652 39264 101704
rect 39316 101692 39322 101704
rect 43030 101692 43036 101704
rect 39316 101664 43036 101692
rect 39316 101652 39322 101664
rect 43030 101652 43036 101664
rect 43088 101652 43094 101704
rect 117642 101652 117648 101704
rect 117700 101692 117706 101704
rect 119850 101692 119856 101704
rect 117700 101664 119856 101692
rect 117700 101652 117706 101664
rect 119850 101652 119856 101664
rect 119908 101652 119914 101704
rect 123254 101652 123260 101704
rect 123312 101692 123318 101704
rect 126474 101692 126480 101704
rect 123312 101664 126480 101692
rect 123312 101652 123318 101664
rect 126474 101652 126480 101664
rect 126532 101652 126538 101704
rect 204490 101652 204496 101704
rect 204548 101692 204554 101704
rect 207250 101692 207256 101704
rect 204548 101664 207256 101692
rect 204548 101652 204554 101664
rect 207250 101652 207256 101664
rect 207308 101652 207314 101704
rect 36038 101584 36044 101636
rect 36096 101624 36102 101636
rect 37510 101624 37516 101636
rect 36096 101596 37516 101624
rect 36096 101584 36102 101596
rect 37510 101584 37516 101596
rect 37568 101584 37574 101636
rect 38430 101584 38436 101636
rect 38488 101624 38494 101636
rect 41834 101624 41840 101636
rect 38488 101596 41840 101624
rect 38488 101584 38494 101596
rect 41834 101584 41840 101596
rect 41892 101584 41898 101636
rect 116814 101584 116820 101636
rect 116872 101624 116878 101636
rect 119390 101624 119396 101636
rect 116872 101596 119396 101624
rect 116872 101584 116878 101596
rect 119390 101584 119396 101596
rect 119448 101584 119454 101636
rect 123622 101584 123628 101636
rect 123680 101624 123686 101636
rect 126566 101624 126572 101636
rect 123680 101596 126572 101624
rect 123680 101584 123686 101596
rect 126566 101584 126572 101596
rect 126624 101584 126630 101636
rect 159318 101584 159324 101636
rect 159376 101624 159382 101636
rect 161710 101624 161716 101636
rect 159376 101596 161716 101624
rect 159376 101584 159382 101596
rect 161710 101584 161716 101596
rect 161768 101584 161774 101636
rect 205686 101584 205692 101636
rect 205744 101624 205750 101636
rect 208906 101624 208912 101636
rect 205744 101596 208912 101624
rect 205744 101584 205750 101596
rect 208906 101584 208912 101596
rect 208964 101584 208970 101636
rect 40454 101516 40460 101568
rect 40512 101556 40518 101568
rect 44870 101556 44876 101568
rect 40512 101528 44876 101556
rect 40512 101516 40518 101528
rect 44870 101516 44876 101528
rect 44928 101516 44934 101568
rect 75322 101516 75328 101568
rect 75380 101556 75386 101568
rect 77530 101556 77536 101568
rect 75380 101528 77536 101556
rect 75380 101516 75386 101528
rect 77530 101516 77536 101528
rect 77588 101516 77594 101568
rect 118838 101516 118844 101568
rect 118896 101556 118902 101568
rect 119942 101556 119948 101568
rect 118896 101528 119948 101556
rect 118896 101516 118902 101528
rect 119942 101516 119948 101528
rect 120000 101516 120006 101568
rect 124818 101516 124824 101568
rect 124876 101556 124882 101568
rect 129234 101556 129240 101568
rect 124876 101528 129240 101556
rect 124876 101516 124882 101528
rect 129234 101516 129240 101528
rect 129292 101516 129298 101568
rect 207618 101516 207624 101568
rect 207676 101556 207682 101568
rect 208170 101556 208176 101568
rect 207676 101528 208176 101556
rect 207676 101516 207682 101528
rect 208170 101516 208176 101528
rect 208228 101516 208234 101568
rect 38890 101448 38896 101500
rect 38948 101488 38954 101500
rect 42294 101488 42300 101500
rect 38948 101460 42300 101488
rect 38948 101448 38954 101460
rect 42294 101448 42300 101460
rect 42352 101448 42358 101500
rect 118470 101448 118476 101500
rect 118528 101488 118534 101500
rect 119758 101488 119764 101500
rect 118528 101460 119764 101488
rect 118528 101448 118534 101460
rect 119758 101448 119764 101460
rect 119816 101448 119822 101500
rect 124082 101448 124088 101500
rect 124140 101488 124146 101500
rect 126658 101488 126664 101500
rect 124140 101460 126664 101488
rect 124140 101448 124146 101460
rect 126658 101448 126664 101460
rect 126716 101448 126722 101500
rect 206054 101448 206060 101500
rect 206112 101488 206118 101500
rect 208630 101488 208636 101500
rect 206112 101460 208636 101488
rect 206112 101448 206118 101460
rect 208630 101448 208636 101460
rect 208688 101448 208694 101500
rect 41282 101380 41288 101432
rect 41340 101420 41346 101432
rect 45054 101420 45060 101432
rect 41340 101392 45060 101420
rect 41340 101380 41346 101392
rect 45054 101380 45060 101392
rect 45112 101380 45118 101432
rect 72378 101380 72384 101432
rect 72436 101420 72442 101432
rect 73482 101420 73488 101432
rect 72436 101392 73488 101420
rect 72436 101380 72442 101392
rect 73482 101380 73488 101392
rect 73540 101380 73546 101432
rect 77530 101380 77536 101432
rect 77588 101420 77594 101432
rect 79646 101420 79652 101432
rect 77588 101392 79652 101420
rect 77588 101380 77594 101392
rect 79646 101380 79652 101392
rect 79704 101380 79710 101432
rect 80842 101380 80848 101432
rect 80900 101420 80906 101432
rect 82314 101420 82320 101432
rect 80900 101392 82320 101420
rect 80900 101380 80906 101392
rect 82314 101380 82320 101392
rect 82372 101380 82378 101432
rect 117274 101380 117280 101432
rect 117332 101420 117338 101432
rect 118930 101420 118936 101432
rect 117332 101392 118936 101420
rect 117332 101380 117338 101392
rect 118930 101380 118936 101392
rect 118988 101380 118994 101432
rect 119298 101380 119304 101432
rect 119356 101420 119362 101432
rect 120954 101420 120960 101432
rect 119356 101392 120960 101420
rect 119356 101380 119362 101392
rect 120954 101380 120960 101392
rect 121012 101380 121018 101432
rect 125646 101380 125652 101432
rect 125704 101420 125710 101432
rect 131534 101420 131540 101432
rect 125704 101392 131540 101420
rect 125704 101380 125710 101392
rect 131534 101380 131540 101392
rect 131592 101380 131598 101432
rect 154902 101380 154908 101432
rect 154960 101420 154966 101432
rect 156190 101420 156196 101432
rect 154960 101392 156196 101420
rect 154960 101380 154966 101392
rect 156190 101380 156196 101392
rect 156248 101380 156254 101432
rect 158214 101380 158220 101432
rect 158272 101420 158278 101432
rect 158858 101420 158864 101432
rect 158272 101392 158864 101420
rect 158272 101380 158278 101392
rect 158858 101380 158864 101392
rect 158916 101380 158922 101432
rect 163734 101380 163740 101432
rect 163792 101420 163798 101432
rect 165114 101420 165120 101432
rect 163792 101392 165120 101420
rect 163792 101380 163798 101392
rect 165114 101380 165120 101392
rect 165172 101380 165178 101432
rect 165942 101380 165948 101432
rect 166000 101420 166006 101432
rect 167874 101420 167880 101432
rect 166000 101392 167880 101420
rect 166000 101380 166006 101392
rect 167874 101380 167880 101392
rect 167932 101380 167938 101432
rect 176154 101380 176160 101432
rect 176212 101420 176218 101432
rect 179282 101420 179288 101432
rect 176212 101392 179288 101420
rect 176212 101380 176218 101392
rect 179282 101380 179288 101392
rect 179340 101380 179346 101432
rect 193358 101380 193364 101432
rect 193416 101420 193422 101432
rect 194462 101420 194468 101432
rect 193416 101392 194468 101420
rect 193416 101380 193422 101392
rect 194462 101380 194468 101392
rect 194520 101380 194526 101432
rect 207250 101380 207256 101432
rect 207308 101420 207314 101432
rect 208354 101420 208360 101432
rect 207308 101392 208360 101420
rect 207308 101380 207314 101392
rect 208354 101380 208360 101392
rect 208412 101380 208418 101432
rect 68606 101312 68612 101364
rect 68664 101352 68670 101364
rect 69250 101352 69256 101364
rect 68664 101324 69256 101352
rect 68664 101312 68670 101324
rect 69250 101312 69256 101324
rect 69308 101312 69314 101364
rect 69802 101312 69808 101364
rect 69860 101352 69866 101364
rect 70630 101352 70636 101364
rect 69860 101324 70636 101352
rect 69860 101312 69866 101324
rect 70630 101312 70636 101324
rect 70688 101312 70694 101364
rect 70906 101312 70912 101364
rect 70964 101352 70970 101364
rect 72010 101352 72016 101364
rect 70964 101324 72016 101352
rect 70964 101312 70970 101324
rect 72010 101312 72016 101324
rect 72068 101312 72074 101364
rect 73114 101312 73120 101364
rect 73172 101352 73178 101364
rect 74034 101352 74040 101364
rect 73172 101324 74040 101352
rect 73172 101312 73178 101324
rect 74034 101312 74040 101324
rect 74092 101312 74098 101364
rect 76426 101312 76432 101364
rect 76484 101352 76490 101364
rect 77438 101352 77444 101364
rect 76484 101324 77444 101352
rect 76484 101312 76490 101324
rect 77438 101312 77444 101324
rect 77496 101312 77502 101364
rect 78634 101312 78640 101364
rect 78692 101352 78698 101364
rect 79554 101352 79560 101364
rect 78692 101324 79560 101352
rect 78692 101312 78698 101324
rect 79554 101312 79560 101324
rect 79612 101312 79618 101364
rect 79738 101312 79744 101364
rect 79796 101352 79802 101364
rect 80934 101352 80940 101364
rect 79796 101324 80940 101352
rect 79796 101312 79802 101324
rect 80934 101312 80940 101324
rect 80992 101312 80998 101364
rect 81946 101312 81952 101364
rect 82004 101352 82010 101364
rect 83694 101352 83700 101364
rect 82004 101324 83700 101352
rect 82004 101312 82010 101324
rect 83694 101312 83700 101324
rect 83752 101312 83758 101364
rect 89766 101312 89772 101364
rect 89824 101352 89830 101364
rect 90594 101352 90600 101364
rect 89824 101324 90600 101352
rect 89824 101312 89830 101324
rect 90594 101312 90600 101324
rect 90652 101312 90658 101364
rect 91974 101312 91980 101364
rect 92032 101352 92038 101364
rect 92618 101352 92624 101364
rect 92032 101324 92624 101352
rect 92032 101312 92038 101324
rect 92618 101312 92624 101324
rect 92676 101312 92682 101364
rect 93078 101312 93084 101364
rect 93136 101352 93142 101364
rect 93998 101352 94004 101364
rect 93136 101324 94004 101352
rect 93136 101312 93142 101324
rect 93998 101312 94004 101324
rect 94056 101312 94062 101364
rect 118102 101312 118108 101364
rect 118160 101352 118166 101364
rect 119574 101352 119580 101364
rect 118160 101324 119580 101352
rect 118160 101312 118166 101324
rect 119574 101312 119580 101324
rect 119632 101312 119638 101364
rect 125278 101312 125284 101364
rect 125336 101352 125342 101364
rect 129326 101352 129332 101364
rect 125336 101324 129332 101352
rect 125336 101312 125342 101324
rect 129326 101312 129332 101324
rect 129384 101312 129390 101364
rect 135214 101312 135220 101364
rect 135272 101352 135278 101364
rect 140458 101352 140464 101364
rect 135272 101324 140464 101352
rect 135272 101312 135278 101324
rect 140458 101312 140464 101324
rect 140516 101312 140522 101364
rect 152602 101312 152608 101364
rect 152660 101352 152666 101364
rect 153430 101352 153436 101364
rect 152660 101324 153436 101352
rect 152660 101312 152666 101324
rect 153430 101312 153436 101324
rect 153488 101312 153494 101364
rect 153798 101312 153804 101364
rect 153856 101352 153862 101364
rect 154810 101352 154816 101364
rect 153856 101324 154816 101352
rect 153856 101312 153862 101324
rect 154810 101312 154816 101324
rect 154868 101312 154874 101364
rect 156006 101312 156012 101364
rect 156064 101352 156070 101364
rect 156834 101352 156840 101364
rect 156064 101324 156840 101352
rect 156064 101312 156070 101324
rect 156834 101312 156840 101324
rect 156892 101312 156898 101364
rect 157110 101312 157116 101364
rect 157168 101352 157174 101364
rect 158306 101352 158312 101364
rect 157168 101324 158312 101352
rect 157168 101312 157174 101324
rect 158306 101312 158312 101324
rect 158364 101312 158370 101364
rect 160422 101312 160428 101364
rect 160480 101352 160486 101364
rect 161618 101352 161624 101364
rect 160480 101324 161624 101352
rect 160480 101312 160486 101324
rect 161618 101312 161624 101324
rect 161676 101312 161682 101364
rect 162630 101312 162636 101364
rect 162688 101352 162694 101364
rect 163826 101352 163832 101364
rect 162688 101324 163832 101352
rect 162688 101312 162694 101324
rect 163826 101312 163832 101324
rect 163884 101312 163890 101364
rect 164838 101312 164844 101364
rect 164896 101352 164902 101364
rect 166494 101352 166500 101364
rect 164896 101324 166500 101352
rect 164896 101312 164902 101324
rect 166494 101312 166500 101324
rect 166552 101312 166558 101364
rect 173762 101312 173768 101364
rect 173820 101352 173826 101364
rect 174774 101352 174780 101364
rect 173820 101324 174780 101352
rect 173820 101312 173826 101324
rect 174774 101312 174780 101324
rect 174832 101312 174838 101364
rect 175970 101312 175976 101364
rect 176028 101352 176034 101364
rect 176798 101352 176804 101364
rect 176028 101324 176804 101352
rect 176028 101312 176034 101324
rect 176798 101312 176804 101324
rect 176856 101312 176862 101364
rect 177074 101312 177080 101364
rect 177132 101352 177138 101364
rect 178178 101352 178184 101364
rect 177132 101324 178184 101352
rect 177132 101312 177138 101324
rect 178178 101312 178184 101324
rect 178236 101312 178242 101364
rect 194646 101312 194652 101364
rect 194704 101352 194710 101364
rect 194704 101324 194876 101352
rect 194704 101312 194710 101324
rect 194848 101216 194876 101324
rect 194922 101312 194928 101364
rect 194980 101352 194986 101364
rect 196026 101352 196032 101364
rect 194980 101324 196032 101352
rect 194980 101312 194986 101324
rect 196026 101312 196032 101324
rect 196084 101312 196090 101364
rect 208078 101312 208084 101364
rect 208136 101352 208142 101364
rect 208538 101352 208544 101364
rect 208136 101324 208544 101352
rect 208136 101312 208142 101324
rect 208538 101312 208544 101324
rect 208596 101312 208602 101364
rect 194922 101216 194928 101228
rect 194848 101188 194928 101216
rect 194922 101176 194928 101188
rect 194980 101176 194986 101228
rect 98782 97164 98788 97216
rect 98840 97204 98846 97216
rect 106786 97204 106792 97216
rect 98840 97176 106792 97204
rect 98840 97164 98846 97176
rect 106786 97164 106792 97176
rect 106844 97164 106850 97216
rect 18098 97096 18104 97148
rect 18156 97136 18162 97148
rect 22330 97136 22336 97148
rect 18156 97108 22336 97136
rect 18156 97096 18162 97108
rect 22330 97096 22336 97108
rect 22388 97096 22394 97148
rect 212310 97096 212316 97148
rect 212368 97136 212374 97148
rect 220958 97136 220964 97148
rect 212368 97108 220964 97136
rect 212368 97096 212374 97108
rect 220958 97096 220964 97108
rect 221016 97096 221022 97148
rect 99518 95804 99524 95856
rect 99576 95844 99582 95856
rect 106786 95844 106792 95856
rect 99576 95816 106792 95844
rect 99576 95804 99582 95816
rect 106786 95804 106792 95816
rect 106844 95804 106850 95856
rect 188574 94376 188580 94428
rect 188632 94416 188638 94428
rect 191978 94416 191984 94428
rect 188632 94388 191984 94416
rect 188632 94376 188638 94388
rect 191978 94376 191984 94388
rect 192036 94376 192042 94428
rect 98690 93016 98696 93068
rect 98748 93056 98754 93068
rect 106510 93056 106516 93068
rect 98748 93028 106516 93056
rect 98748 93016 98754 93028
rect 106510 93016 106516 93028
rect 106568 93016 106574 93068
rect 105038 90228 105044 90280
rect 105096 90268 105102 90280
rect 106786 90268 106792 90280
rect 105096 90240 106792 90268
rect 105096 90228 105102 90240
rect 106786 90228 106792 90240
rect 106844 90228 106850 90280
rect 13314 90160 13320 90212
rect 13372 90200 13378 90212
rect 22330 90200 22336 90212
rect 13372 90172 22336 90200
rect 13372 90160 13378 90172
rect 22330 90160 22336 90172
rect 22388 90160 22394 90212
rect 182870 90160 182876 90212
rect 182928 90200 182934 90212
rect 188574 90200 188580 90212
rect 182928 90172 188580 90200
rect 182928 90160 182934 90172
rect 188574 90160 188580 90172
rect 188632 90160 188638 90212
rect 104946 88868 104952 88920
rect 105004 88908 105010 88920
rect 106786 88908 106792 88920
rect 105004 88880 106792 88908
rect 105004 88868 105010 88880
rect 106786 88868 106792 88880
rect 106844 88868 106850 88920
rect 128498 88868 128504 88920
rect 128556 88908 128562 88920
rect 131994 88908 132000 88920
rect 128556 88880 132000 88908
rect 128556 88868 128562 88880
rect 131994 88868 132000 88880
rect 132052 88868 132058 88920
rect 183514 88800 183520 88852
rect 183572 88840 183578 88852
rect 191150 88840 191156 88852
rect 183572 88812 191156 88840
rect 183572 88800 183578 88812
rect 191150 88800 191156 88812
rect 191208 88800 191214 88852
rect 183698 87440 183704 87492
rect 183756 87480 183762 87492
rect 190782 87480 190788 87492
rect 183756 87452 190788 87480
rect 183756 87440 183762 87452
rect 190782 87440 190788 87452
rect 190840 87440 190846 87492
rect 183698 86012 183704 86064
rect 183756 86052 183762 86064
rect 191702 86052 191708 86064
rect 183756 86024 191708 86052
rect 183756 86012 183762 86024
rect 191702 86012 191708 86024
rect 191760 86012 191766 86064
rect 99518 85196 99524 85248
rect 99576 85236 99582 85248
rect 105038 85236 105044 85248
rect 99576 85208 105044 85236
rect 99576 85196 99582 85208
rect 105038 85196 105044 85208
rect 105096 85196 105102 85248
rect 44410 84720 44416 84772
rect 44468 84760 44474 84772
rect 52690 84760 52696 84772
rect 44468 84732 52696 84760
rect 44468 84720 44474 84732
rect 52690 84720 52696 84732
rect 52748 84720 52754 84772
rect 99426 84652 99432 84704
rect 99484 84692 99490 84704
rect 106786 84692 106792 84704
rect 99484 84664 106792 84692
rect 99484 84652 99490 84664
rect 106786 84652 106792 84664
rect 106844 84652 106850 84704
rect 182502 84652 182508 84704
rect 182560 84692 182566 84704
rect 191978 84692 191984 84704
rect 182560 84664 191984 84692
rect 182560 84652 182566 84664
rect 191978 84652 191984 84664
rect 192036 84652 192042 84704
rect 99518 84584 99524 84636
rect 99576 84624 99582 84636
rect 104946 84624 104952 84636
rect 99576 84596 104952 84624
rect 99576 84584 99582 84596
rect 104946 84584 104952 84596
rect 105004 84584 105010 84636
rect 183698 84584 183704 84636
rect 183756 84624 183762 84636
rect 191610 84624 191616 84636
rect 183756 84596 191616 84624
rect 183756 84584 183762 84596
rect 191610 84584 191616 84596
rect 191668 84584 191674 84636
rect 13406 83292 13412 83344
rect 13464 83332 13470 83344
rect 22330 83332 22336 83344
rect 13464 83304 22336 83332
rect 13464 83292 13470 83304
rect 22330 83292 22336 83304
rect 22388 83292 22394 83344
rect 99518 83292 99524 83344
rect 99576 83332 99582 83344
rect 107798 83332 107804 83344
rect 99576 83304 107804 83332
rect 99576 83292 99582 83304
rect 107798 83292 107804 83304
rect 107856 83292 107862 83344
rect 183698 82612 183704 82664
rect 183756 82652 183762 82664
rect 191978 82652 191984 82664
rect 183756 82624 191984 82652
rect 183756 82612 183762 82624
rect 191978 82612 191984 82624
rect 192036 82612 192042 82664
rect 106786 82108 106792 82120
rect 103768 82080 106792 82108
rect 99518 81932 99524 81984
rect 99576 81972 99582 81984
rect 103768 81972 103796 82080
rect 106786 82068 106792 82080
rect 106844 82068 106850 82120
rect 99576 81944 103796 81972
rect 99576 81932 99582 81944
rect 183238 81252 183244 81304
rect 183296 81292 183302 81304
rect 191886 81292 191892 81304
rect 183296 81264 191892 81292
rect 183296 81252 183302 81264
rect 191886 81252 191892 81264
rect 191944 81252 191950 81304
rect 131994 80504 132000 80556
rect 132052 80544 132058 80556
rect 136870 80544 136876 80556
rect 132052 80516 136876 80544
rect 132052 80504 132058 80516
rect 136870 80504 136876 80516
rect 136928 80504 136934 80556
rect 99518 79824 99524 79876
rect 99576 79864 99582 79876
rect 106786 79864 106792 79876
rect 99576 79836 106792 79864
rect 99576 79824 99582 79836
rect 106786 79824 106792 79836
rect 106844 79824 106850 79876
rect 183698 79212 183704 79264
rect 183756 79252 183762 79264
rect 183756 79224 187976 79252
rect 183756 79212 183762 79224
rect 187948 79184 187976 79224
rect 191978 79184 191984 79196
rect 187948 79156 191984 79184
rect 191978 79144 191984 79156
rect 192036 79144 192042 79196
rect 99518 77852 99524 77904
rect 99576 77892 99582 77904
rect 106510 77892 106516 77904
rect 99576 77864 106516 77892
rect 99576 77852 99582 77864
rect 106510 77852 106516 77864
rect 106568 77852 106574 77904
rect 183514 77852 183520 77904
rect 183572 77892 183578 77904
rect 191978 77892 191984 77904
rect 183572 77864 191984 77892
rect 183572 77852 183578 77864
rect 191978 77852 191984 77864
rect 192036 77852 192042 77904
rect 13498 77784 13504 77836
rect 13556 77824 13562 77836
rect 22330 77824 22336 77836
rect 13556 77796 22336 77824
rect 13556 77784 13562 77796
rect 22330 77784 22336 77796
rect 22388 77784 22394 77836
rect 99518 76424 99524 76476
rect 99576 76464 99582 76476
rect 100990 76464 100996 76476
rect 99576 76436 100996 76464
rect 99576 76424 99582 76436
rect 100990 76424 100996 76436
rect 101048 76424 101054 76476
rect 183054 76424 183060 76476
rect 183112 76464 183118 76476
rect 185170 76464 185176 76476
rect 183112 76436 185176 76464
rect 183112 76424 183118 76436
rect 185170 76424 185176 76436
rect 185228 76424 185234 76476
rect 98230 75064 98236 75116
rect 98288 75104 98294 75116
rect 98288 75076 100944 75104
rect 98288 75064 98294 75076
rect 100916 74900 100944 75076
rect 183238 75064 183244 75116
rect 183296 75104 183302 75116
rect 186182 75104 186188 75116
rect 183296 75076 186188 75104
rect 183296 75064 183302 75076
rect 186182 75064 186188 75076
rect 186240 75064 186246 75116
rect 100990 74996 100996 75048
rect 101048 75036 101054 75048
rect 106786 75036 106792 75048
rect 101048 75008 106792 75036
rect 101048 74996 101054 75008
rect 106786 74996 106792 75008
rect 106844 74996 106850 75048
rect 185170 74996 185176 75048
rect 185228 75036 185234 75048
rect 191518 75036 191524 75048
rect 185228 75008 191524 75036
rect 185228 74996 185234 75008
rect 191518 74996 191524 75008
rect 191576 74996 191582 75048
rect 212126 74996 212132 75048
rect 212184 75036 212190 75048
rect 222338 75036 222344 75048
rect 212184 75008 222344 75036
rect 212184 74996 212190 75008
rect 222338 74996 222344 75008
rect 222396 74996 222402 75048
rect 100990 74900 100996 74912
rect 100916 74872 100996 74900
rect 100990 74860 100996 74872
rect 101048 74860 101054 74912
rect 44410 74316 44416 74368
rect 44468 74356 44474 74368
rect 53334 74356 53340 74368
rect 44468 74328 53340 74356
rect 44468 74316 44474 74328
rect 53334 74316 53340 74328
rect 53392 74316 53398 74368
rect 99518 73840 99524 73892
rect 99576 73880 99582 73892
rect 105130 73880 105136 73892
rect 99576 73852 105136 73880
rect 99576 73840 99582 73852
rect 105130 73840 105136 73852
rect 105188 73840 105194 73892
rect 183698 73840 183704 73892
rect 183756 73880 183762 73892
rect 183756 73852 188620 73880
rect 183756 73840 183762 73852
rect 99426 73704 99432 73756
rect 99484 73744 99490 73756
rect 106694 73744 106700 73756
rect 99484 73716 106700 73744
rect 99484 73704 99490 73716
rect 106694 73704 106700 73716
rect 106752 73704 106758 73756
rect 183698 73704 183704 73756
rect 183756 73744 183762 73756
rect 188482 73744 188488 73756
rect 183756 73716 188488 73744
rect 183756 73704 183762 73716
rect 188482 73704 188488 73716
rect 188540 73704 188546 73756
rect 188592 73744 188620 73852
rect 190782 73744 190788 73756
rect 188592 73716 190788 73744
rect 190782 73704 190788 73716
rect 190840 73704 190846 73756
rect 100990 73636 100996 73688
rect 101048 73676 101054 73688
rect 106786 73676 106792 73688
rect 101048 73648 106792 73676
rect 101048 73636 101054 73648
rect 106786 73636 106792 73648
rect 106844 73636 106850 73688
rect 186182 73636 186188 73688
rect 186240 73676 186246 73688
rect 191978 73676 191984 73688
rect 186240 73648 191984 73676
rect 186240 73636 186246 73648
rect 191978 73636 191984 73648
rect 192036 73636 192042 73688
rect 99518 72344 99524 72396
rect 99576 72384 99582 72396
rect 106510 72384 106516 72396
rect 99576 72356 106516 72384
rect 99576 72344 99582 72356
rect 106510 72344 106516 72356
rect 106568 72344 106574 72396
rect 99518 70984 99524 71036
rect 99576 71024 99582 71036
rect 104486 71024 104492 71036
rect 99576 70996 104492 71024
rect 99576 70984 99582 70996
rect 104486 70984 104492 70996
rect 104544 70984 104550 71036
rect 183698 70916 183704 70968
rect 183756 70956 183762 70968
rect 191518 70956 191524 70968
rect 183756 70928 191524 70956
rect 183756 70916 183762 70928
rect 191518 70916 191524 70928
rect 191576 70916 191582 70968
rect 128498 70168 128504 70220
rect 128556 70208 128562 70220
rect 133374 70208 133380 70220
rect 128556 70180 133380 70208
rect 128556 70168 128562 70180
rect 133374 70168 133380 70180
rect 133432 70208 133438 70220
rect 136870 70208 136876 70220
rect 133432 70180 136876 70208
rect 133432 70168 133438 70180
rect 136870 70168 136876 70180
rect 136928 70168 136934 70220
rect 182870 69896 182876 69948
rect 182928 69936 182934 69948
rect 189954 69936 189960 69948
rect 182928 69908 189960 69936
rect 182928 69896 182934 69908
rect 189954 69896 189960 69908
rect 190012 69896 190018 69948
rect 212678 69760 212684 69812
rect 212736 69800 212742 69812
rect 215622 69800 215628 69812
rect 212736 69772 215628 69800
rect 212736 69760 212742 69772
rect 215622 69760 215628 69772
rect 215680 69760 215686 69812
rect 99518 69556 99524 69608
rect 99576 69596 99582 69608
rect 104394 69596 104400 69608
rect 99576 69568 104400 69596
rect 99576 69556 99582 69568
rect 104394 69556 104400 69568
rect 104452 69556 104458 69608
rect 188482 69488 188488 69540
rect 188540 69528 188546 69540
rect 190966 69528 190972 69540
rect 188540 69500 190972 69528
rect 188540 69488 188546 69500
rect 190966 69488 190972 69500
rect 191024 69488 191030 69540
rect 105130 68128 105136 68180
rect 105188 68168 105194 68180
rect 106602 68168 106608 68180
rect 105188 68140 106608 68168
rect 105188 68128 105194 68140
rect 106602 68128 106608 68140
rect 106660 68128 106666 68180
rect 183790 68128 183796 68180
rect 183848 68168 183854 68180
rect 191334 68168 191340 68180
rect 183848 68140 191340 68168
rect 183848 68128 183854 68140
rect 191334 68128 191340 68140
rect 191392 68128 191398 68180
rect 104486 63640 104492 63692
rect 104544 63680 104550 63692
rect 106602 63680 106608 63692
rect 104544 63652 106608 63680
rect 104544 63640 104550 63652
rect 106602 63640 106608 63652
rect 106660 63640 106666 63692
rect 183698 61464 183704 61516
rect 183756 61504 183762 61516
rect 188022 61504 188028 61516
rect 183756 61476 188028 61504
rect 183756 61464 183762 61476
rect 188022 61464 188028 61476
rect 188080 61464 188086 61516
rect 99518 61328 99524 61380
rect 99576 61368 99582 61380
rect 105314 61368 105320 61380
rect 99576 61340 105320 61368
rect 99576 61328 99582 61340
rect 105314 61328 105320 61340
rect 105372 61328 105378 61380
rect 104394 61192 104400 61244
rect 104452 61232 104458 61244
rect 107154 61232 107160 61244
rect 104452 61204 107160 61232
rect 104452 61192 104458 61204
rect 107154 61192 107160 61204
rect 107212 61192 107218 61244
rect 182686 60376 182692 60428
rect 182744 60416 182750 60428
rect 184434 60416 184440 60428
rect 182744 60388 184440 60416
rect 182744 60376 182750 60388
rect 184434 60376 184440 60388
rect 184492 60376 184498 60428
rect 26746 59968 26752 60020
rect 26804 60008 26810 60020
rect 26930 60008 26936 60020
rect 26804 59980 26936 60008
rect 26804 59968 26810 59980
rect 26930 59968 26936 59980
rect 26988 59968 26994 60020
rect 137974 59832 137980 59884
rect 138032 59872 138038 59884
rect 138158 59872 138164 59884
rect 138032 59844 138164 59872
rect 138032 59832 138038 59844
rect 138158 59832 138164 59844
rect 138216 59832 138222 59884
rect 112398 58540 112404 58592
rect 112456 58580 112462 58592
rect 112858 58580 112864 58592
rect 112456 58552 112864 58580
rect 112456 58540 112462 58552
rect 112858 58540 112864 58552
rect 112916 58540 112922 58592
rect 36130 58472 36136 58524
rect 36188 58512 36194 58524
rect 37602 58512 37608 58524
rect 36188 58484 37608 58512
rect 36188 58472 36194 58484
rect 37602 58472 37608 58484
rect 37660 58472 37666 58524
rect 79186 58472 79192 58524
rect 79244 58512 79250 58524
rect 96114 58512 96120 58524
rect 79244 58484 96120 58512
rect 79244 58472 79250 58484
rect 96114 58472 96120 58484
rect 96172 58512 96178 58524
rect 163182 58512 163188 58524
rect 96172 58484 163188 58512
rect 96172 58472 96178 58484
rect 163182 58472 163188 58484
rect 163240 58472 163246 58524
rect 199614 58472 199620 58524
rect 199672 58512 199678 58524
rect 200350 58512 200356 58524
rect 199672 58484 200356 58512
rect 199672 58472 199678 58484
rect 200350 58472 200356 58484
rect 200408 58472 200414 58524
rect 208078 58472 208084 58524
rect 208136 58512 208142 58524
rect 210654 58512 210660 58524
rect 208136 58484 210660 58512
rect 208136 58472 208142 58484
rect 210654 58472 210660 58484
rect 210712 58472 210718 58524
rect 41282 58404 41288 58456
rect 41340 58444 41346 58456
rect 45882 58444 45888 58456
rect 41340 58416 45888 58444
rect 41340 58404 41346 58416
rect 45882 58404 45888 58416
rect 45940 58404 45946 58456
rect 72562 58404 72568 58456
rect 72620 58444 72626 58456
rect 98874 58444 98880 58456
rect 72620 58416 98880 58444
rect 72620 58404 72626 58416
rect 98874 58404 98880 58416
rect 98932 58444 98938 58456
rect 156558 58444 156564 58456
rect 98932 58416 156564 58444
rect 98932 58404 98938 58416
rect 156558 58404 156564 58416
rect 156616 58404 156622 58456
rect 209642 58404 209648 58456
rect 209700 58444 209706 58456
rect 212310 58444 212316 58456
rect 209700 58416 212316 58444
rect 209700 58404 209706 58416
rect 212310 58404 212316 58416
rect 212368 58404 212374 58456
rect 41650 58336 41656 58388
rect 41708 58376 41714 58388
rect 46434 58376 46440 58388
rect 41708 58348 46440 58376
rect 41708 58336 41714 58348
rect 46434 58336 46440 58348
rect 46492 58336 46498 58388
rect 121230 58336 121236 58388
rect 121288 58376 121294 58388
rect 123714 58376 123720 58388
rect 121288 58348 123720 58376
rect 121288 58336 121294 58348
rect 123714 58336 123720 58348
rect 123772 58336 123778 58388
rect 207618 58336 207624 58388
rect 207676 58376 207682 58388
rect 210746 58376 210752 58388
rect 207676 58348 210752 58376
rect 207676 58336 207682 58348
rect 210746 58336 210752 58348
rect 210804 58336 210810 58388
rect 122426 58268 122432 58320
rect 122484 58308 122490 58320
rect 125094 58308 125100 58320
rect 122484 58280 125100 58308
rect 122484 58268 122490 58280
rect 125094 58268 125100 58280
rect 125152 58268 125158 58320
rect 208814 58268 208820 58320
rect 208872 58308 208878 58320
rect 212218 58308 212224 58320
rect 208872 58280 212224 58308
rect 208872 58268 208878 58280
rect 212218 58268 212224 58280
rect 212276 58268 212282 58320
rect 123254 58200 123260 58252
rect 123312 58240 123318 58252
rect 127302 58240 127308 58252
rect 123312 58212 127308 58240
rect 123312 58200 123318 58212
rect 127302 58200 127308 58212
rect 127360 58200 127366 58252
rect 207250 58200 207256 58252
rect 207308 58240 207314 58252
rect 210838 58240 210844 58252
rect 207308 58212 210844 58240
rect 207308 58200 207314 58212
rect 210838 58200 210844 58212
rect 210896 58200 210902 58252
rect 120494 58064 120500 58116
rect 120552 58104 120558 58116
rect 123254 58104 123260 58116
rect 120552 58076 123260 58104
rect 120552 58064 120558 58076
rect 123254 58064 123260 58076
rect 123312 58064 123318 58116
rect 209274 58064 209280 58116
rect 209332 58104 209338 58116
rect 212126 58104 212132 58116
rect 209332 58076 212132 58104
rect 209332 58064 209338 58076
rect 212126 58064 212132 58076
rect 212184 58064 212190 58116
rect 120862 57928 120868 57980
rect 120920 57968 120926 57980
rect 123438 57968 123444 57980
rect 120920 57940 123444 57968
rect 120920 57928 120926 57940
rect 123438 57928 123444 57940
rect 123496 57928 123502 57980
rect 70538 57860 70544 57912
rect 70596 57900 70602 57912
rect 92526 57900 92532 57912
rect 70596 57872 92532 57900
rect 70596 57860 70602 57872
rect 92526 57860 92532 57872
rect 92584 57860 92590 57912
rect 13314 57792 13320 57844
rect 13372 57832 13378 57844
rect 72562 57832 72568 57844
rect 13372 57804 72568 57832
rect 13372 57792 13378 57804
rect 72562 57792 72568 57804
rect 72620 57792 72626 57844
rect 122058 57792 122064 57844
rect 122116 57832 122122 57844
rect 125186 57832 125192 57844
rect 122116 57804 125192 57832
rect 122116 57792 122122 57804
rect 125186 57792 125192 57804
rect 125244 57792 125250 57844
rect 156098 57792 156104 57844
rect 156156 57832 156162 57844
rect 169898 57832 169904 57844
rect 156156 57804 169904 57832
rect 156156 57792 156162 57804
rect 169898 57792 169904 57804
rect 169956 57792 169962 57844
rect 208446 57792 208452 57844
rect 208504 57832 208510 57844
rect 212862 57832 212868 57844
rect 208504 57804 212868 57832
rect 208504 57792 208510 57804
rect 212862 57792 212868 57804
rect 212920 57792 212926 57844
rect 40822 57724 40828 57776
rect 40880 57764 40886 57776
rect 45790 57764 45796 57776
rect 40880 57736 45796 57764
rect 40880 57724 40886 57736
rect 45790 57724 45796 57736
rect 45848 57724 45854 57776
rect 114054 57724 114060 57776
rect 114112 57764 114118 57776
rect 114974 57764 114980 57776
rect 114112 57736 114980 57764
rect 114112 57724 114118 57736
rect 114974 57724 114980 57736
rect 115032 57724 115038 57776
rect 116814 57656 116820 57708
rect 116872 57696 116878 57708
rect 118378 57696 118384 57708
rect 116872 57668 118384 57696
rect 116872 57656 116878 57668
rect 118378 57656 118384 57668
rect 118436 57656 118442 57708
rect 125278 57656 125284 57708
rect 125336 57696 125342 57708
rect 129970 57696 129976 57708
rect 125336 57668 129976 57696
rect 125336 57656 125342 57668
rect 129970 57656 129976 57668
rect 130028 57656 130034 57708
rect 116078 57588 116084 57640
rect 116136 57628 116142 57640
rect 117734 57628 117740 57640
rect 116136 57600 117740 57628
rect 116136 57588 116142 57600
rect 117734 57588 117740 57600
rect 117792 57588 117798 57640
rect 206422 57588 206428 57640
rect 206480 57628 206486 57640
rect 210102 57628 210108 57640
rect 206480 57600 210108 57628
rect 206480 57588 206486 57600
rect 210102 57588 210108 57600
rect 210160 57588 210166 57640
rect 40086 57520 40092 57572
rect 40144 57560 40150 57572
rect 43766 57560 43772 57572
rect 40144 57532 43772 57560
rect 40144 57520 40150 57532
rect 43766 57520 43772 57532
rect 43824 57520 43830 57572
rect 118838 57520 118844 57572
rect 118896 57560 118902 57572
rect 121230 57560 121236 57572
rect 118896 57532 121236 57560
rect 118896 57520 118902 57532
rect 121230 57520 121236 57532
rect 121288 57520 121294 57572
rect 122886 57520 122892 57572
rect 122944 57560 122950 57572
rect 125278 57560 125284 57572
rect 122944 57532 125284 57560
rect 122944 57520 122950 57532
rect 125278 57520 125284 57532
rect 125336 57520 125342 57572
rect 204490 57520 204496 57572
rect 204548 57560 204554 57572
rect 207250 57560 207256 57572
rect 204548 57532 207256 57560
rect 204548 57520 204554 57532
rect 207250 57520 207256 57532
rect 207308 57520 207314 57572
rect 39258 57452 39264 57504
rect 39316 57492 39322 57504
rect 43030 57492 43036 57504
rect 39316 57464 43036 57492
rect 39316 57452 39322 57464
rect 43030 57452 43036 57464
rect 43088 57452 43094 57504
rect 118102 57452 118108 57504
rect 118160 57492 118166 57504
rect 120494 57492 120500 57504
rect 118160 57464 120500 57492
rect 118160 57452 118166 57464
rect 120494 57452 120500 57464
rect 120552 57452 120558 57504
rect 124082 57452 124088 57504
rect 124140 57492 124146 57504
rect 128774 57492 128780 57504
rect 124140 57464 128780 57492
rect 124140 57452 124146 57464
rect 128774 57452 128780 57464
rect 128832 57452 128838 57504
rect 205226 57452 205232 57504
rect 205284 57492 205290 57504
rect 207986 57492 207992 57504
rect 205284 57464 207992 57492
rect 205284 57452 205290 57464
rect 207986 57452 207992 57464
rect 208044 57452 208050 57504
rect 39626 57384 39632 57436
rect 39684 57424 39690 57436
rect 43122 57424 43128 57436
rect 39684 57396 43128 57424
rect 39684 57384 39690 57396
rect 43122 57384 43128 57396
rect 43180 57384 43186 57436
rect 118470 57384 118476 57436
rect 118528 57424 118534 57436
rect 120770 57424 120776 57436
rect 118528 57396 120776 57424
rect 118528 57384 118534 57396
rect 120770 57384 120776 57396
rect 120828 57384 120834 57436
rect 121690 57384 121696 57436
rect 121748 57424 121754 57436
rect 124910 57424 124916 57436
rect 121748 57396 124916 57424
rect 121748 57384 121754 57396
rect 124910 57384 124916 57396
rect 124968 57384 124974 57436
rect 203294 57384 203300 57436
rect 203352 57424 203358 57436
rect 205318 57424 205324 57436
rect 203352 57396 205324 57424
rect 203352 57384 203358 57396
rect 205318 57384 205324 57396
rect 205376 57384 205382 57436
rect 206882 57384 206888 57436
rect 206940 57424 206946 57436
rect 210010 57424 210016 57436
rect 206940 57396 210016 57424
rect 206940 57384 206946 57396
rect 210010 57384 210016 57396
rect 210068 57384 210074 57436
rect 29138 57316 29144 57368
rect 29196 57356 29202 57368
rect 30426 57356 30432 57368
rect 29196 57328 30432 57356
rect 29196 57316 29202 57328
rect 30426 57316 30432 57328
rect 30484 57316 30490 57368
rect 37694 57316 37700 57368
rect 37752 57356 37758 57368
rect 40270 57356 40276 57368
rect 37752 57328 40276 57356
rect 37752 57316 37758 57328
rect 40270 57316 40276 57328
rect 40328 57316 40334 57368
rect 124450 57316 124456 57368
rect 124508 57356 124514 57368
rect 128866 57356 128872 57368
rect 124508 57328 128872 57356
rect 124508 57316 124514 57328
rect 128866 57316 128872 57328
rect 128924 57316 128930 57368
rect 200718 57316 200724 57368
rect 200776 57356 200782 57368
rect 201822 57356 201828 57368
rect 200776 57328 201828 57356
rect 200776 57316 200782 57328
rect 201822 57316 201828 57328
rect 201880 57316 201886 57368
rect 202466 57316 202472 57368
rect 202524 57356 202530 57368
rect 204582 57356 204588 57368
rect 202524 57328 204588 57356
rect 202524 57316 202530 57328
rect 204582 57316 204588 57328
rect 204640 57316 204646 57368
rect 204858 57316 204864 57368
rect 204916 57356 204922 57368
rect 207342 57356 207348 57368
rect 204916 57328 207348 57356
rect 204916 57316 204922 57328
rect 207342 57316 207348 57328
rect 207400 57316 207406 57368
rect 36866 57248 36872 57300
rect 36924 57288 36930 57300
rect 38246 57288 38252 57300
rect 36924 57260 38252 57288
rect 36924 57248 36930 57260
rect 38246 57248 38252 57260
rect 38304 57248 38310 57300
rect 38890 57248 38896 57300
rect 38948 57288 38954 57300
rect 41834 57288 41840 57300
rect 38948 57260 41840 57288
rect 38948 57248 38954 57260
rect 41834 57248 41840 57260
rect 41892 57248 41898 57300
rect 115250 57248 115256 57300
rect 115308 57288 115314 57300
rect 116262 57288 116268 57300
rect 115308 57260 116268 57288
rect 115308 57248 115314 57260
rect 116262 57248 116268 57260
rect 116320 57248 116326 57300
rect 117642 57248 117648 57300
rect 117700 57288 117706 57300
rect 118838 57288 118844 57300
rect 117700 57260 118844 57288
rect 117700 57248 117706 57260
rect 118838 57248 118844 57260
rect 118896 57248 118902 57300
rect 119298 57248 119304 57300
rect 119356 57288 119362 57300
rect 121046 57288 121052 57300
rect 119356 57260 121052 57288
rect 119356 57248 119362 57260
rect 121046 57248 121052 57260
rect 121104 57248 121110 57300
rect 123622 57248 123628 57300
rect 123680 57288 123686 57300
rect 127210 57288 127216 57300
rect 123680 57260 127216 57288
rect 123680 57248 123686 57260
rect 127210 57248 127216 57260
rect 127268 57248 127274 57300
rect 194646 57248 194652 57300
rect 194704 57288 194710 57300
rect 195290 57288 195296 57300
rect 194704 57260 195296 57288
rect 194704 57248 194710 57260
rect 195290 57248 195296 57260
rect 195348 57248 195354 57300
rect 198878 57248 198884 57300
rect 198936 57288 198942 57300
rect 199154 57288 199160 57300
rect 198936 57260 199160 57288
rect 198936 57248 198942 57260
rect 199154 57248 199160 57260
rect 199212 57248 199218 57300
rect 201270 57248 201276 57300
rect 201328 57288 201334 57300
rect 202190 57288 202196 57300
rect 201328 57260 202196 57288
rect 201328 57248 201334 57260
rect 202190 57248 202196 57260
rect 202248 57248 202254 57300
rect 203662 57248 203668 57300
rect 203720 57288 203726 57300
rect 205226 57288 205232 57300
rect 203720 57260 205232 57288
rect 203720 57248 203726 57260
rect 205226 57248 205232 57260
rect 205284 57248 205290 57300
rect 30426 57180 30432 57232
rect 30484 57220 30490 57232
rect 31254 57220 31260 57232
rect 30484 57192 31260 57220
rect 30484 57180 30490 57192
rect 31254 57180 31260 57192
rect 31312 57180 31318 57232
rect 37234 57180 37240 57232
rect 37292 57220 37298 57232
rect 38154 57220 38160 57232
rect 37292 57192 38160 57220
rect 37292 57180 37298 57192
rect 38154 57180 38160 57192
rect 38212 57180 38218 57232
rect 38430 57180 38436 57232
rect 38488 57220 38494 57232
rect 40914 57220 40920 57232
rect 38488 57192 40920 57220
rect 38488 57180 38494 57192
rect 40914 57180 40920 57192
rect 40972 57180 40978 57232
rect 109270 57180 109276 57232
rect 109328 57220 109334 57232
rect 110466 57220 110472 57232
rect 109328 57192 110472 57220
rect 109328 57180 109334 57192
rect 110466 57180 110472 57192
rect 110524 57180 110530 57232
rect 114422 57180 114428 57232
rect 114480 57220 114486 57232
rect 115342 57220 115348 57232
rect 114480 57192 115348 57220
rect 114480 57180 114486 57192
rect 115342 57180 115348 57192
rect 115400 57180 115406 57232
rect 116446 57180 116452 57232
rect 116504 57220 116510 57232
rect 118102 57220 118108 57232
rect 116504 57192 118108 57220
rect 116504 57180 116510 57192
rect 118102 57180 118108 57192
rect 118160 57180 118166 57232
rect 120034 57180 120040 57232
rect 120092 57220 120098 57232
rect 121138 57220 121144 57232
rect 120092 57192 121144 57220
rect 120092 57180 120098 57192
rect 121138 57180 121144 57192
rect 121196 57180 121202 57232
rect 124818 57180 124824 57232
rect 124876 57220 124882 57232
rect 129510 57220 129516 57232
rect 124876 57192 129516 57220
rect 124876 57180 124882 57192
rect 129510 57180 129516 57192
rect 129568 57180 129574 57232
rect 193358 57180 193364 57232
rect 193416 57220 193422 57232
rect 194462 57220 194468 57232
rect 193416 57192 194468 57220
rect 193416 57180 193422 57192
rect 194462 57180 194468 57192
rect 194520 57180 194526 57232
rect 195106 57180 195112 57232
rect 195164 57220 195170 57232
rect 196026 57220 196032 57232
rect 195164 57192 196032 57220
rect 195164 57180 195170 57192
rect 196026 57180 196032 57192
rect 196084 57180 196090 57232
rect 196394 57180 196400 57232
rect 196452 57220 196458 57232
rect 196854 57220 196860 57232
rect 196452 57192 196860 57220
rect 196452 57180 196458 57192
rect 196854 57180 196860 57192
rect 196912 57180 196918 57232
rect 201638 57180 201644 57232
rect 201696 57220 201702 57232
rect 202374 57220 202380 57232
rect 201696 57192 202380 57220
rect 201696 57180 201702 57192
rect 202374 57180 202380 57192
rect 202432 57180 202438 57232
rect 202834 57180 202840 57232
rect 202892 57220 202898 57232
rect 204490 57220 204496 57232
rect 202892 57192 204496 57220
rect 202892 57180 202898 57192
rect 204490 57180 204496 57192
rect 204548 57180 204554 57232
rect 205686 57180 205692 57232
rect 205744 57220 205750 57232
rect 207894 57220 207900 57232
rect 205744 57192 207900 57220
rect 205744 57180 205750 57192
rect 207894 57180 207900 57192
rect 207952 57180 207958 57232
rect 26562 57112 26568 57164
rect 26620 57152 26626 57164
rect 27022 57152 27028 57164
rect 26620 57124 27028 57152
rect 26620 57112 26626 57124
rect 27022 57112 27028 57124
rect 27080 57112 27086 57164
rect 27850 57112 27856 57164
rect 27908 57152 27914 57164
rect 28586 57152 28592 57164
rect 27908 57124 28592 57152
rect 27908 57112 27914 57124
rect 28586 57112 28592 57124
rect 28644 57112 28650 57164
rect 29322 57112 29328 57164
rect 29380 57152 29386 57164
rect 29598 57152 29604 57164
rect 29380 57124 29604 57152
rect 29380 57112 29386 57124
rect 29598 57112 29604 57124
rect 29656 57112 29662 57164
rect 30518 57112 30524 57164
rect 30576 57152 30582 57164
rect 31622 57152 31628 57164
rect 30576 57124 31628 57152
rect 30576 57112 30582 57124
rect 31622 57112 31628 57124
rect 31680 57112 31686 57164
rect 33278 57152 33284 57164
rect 32100 57124 33284 57152
rect 26470 57044 26476 57096
rect 26528 57084 26534 57096
rect 27390 57084 27396 57096
rect 26528 57056 27396 57084
rect 26528 57044 26534 57056
rect 27390 57044 27396 57056
rect 27448 57044 27454 57096
rect 29414 57044 29420 57096
rect 29472 57084 29478 57096
rect 29782 57084 29788 57096
rect 29472 57056 29788 57084
rect 29472 57044 29478 57056
rect 29782 57044 29788 57056
rect 29840 57044 29846 57096
rect 32100 56824 32128 57124
rect 33278 57112 33284 57124
rect 33336 57112 33342 57164
rect 33462 57112 33468 57164
rect 33520 57152 33526 57164
rect 34106 57152 34112 57164
rect 33520 57124 34112 57152
rect 33520 57112 33526 57124
rect 34106 57112 34112 57124
rect 34164 57112 34170 57164
rect 35302 57112 35308 57164
rect 35360 57152 35366 57164
rect 36038 57152 36044 57164
rect 35360 57124 36044 57152
rect 35360 57112 35366 57124
rect 36038 57112 36044 57124
rect 36096 57112 36102 57164
rect 36498 57112 36504 57164
rect 36556 57152 36562 57164
rect 37510 57152 37516 57164
rect 36556 57124 37516 57152
rect 36556 57112 36562 57124
rect 37510 57112 37516 57124
rect 37568 57112 37574 57164
rect 38062 57112 38068 57164
rect 38120 57152 38126 57164
rect 40362 57152 40368 57164
rect 38120 57124 40368 57152
rect 38120 57112 38126 57124
rect 40362 57112 40368 57124
rect 40420 57112 40426 57164
rect 40454 57112 40460 57164
rect 40512 57152 40518 57164
rect 43674 57152 43680 57164
rect 40512 57124 43680 57152
rect 40512 57112 40518 57124
rect 43674 57112 43680 57124
rect 43732 57112 43738 57164
rect 109178 57112 109184 57164
rect 109236 57152 109242 57164
rect 110098 57152 110104 57164
rect 109236 57124 110104 57152
rect 109236 57112 109242 57124
rect 110098 57112 110104 57124
rect 110156 57112 110162 57164
rect 111110 57112 111116 57164
rect 111168 57152 111174 57164
rect 111662 57152 111668 57164
rect 111168 57124 111668 57152
rect 111168 57112 111174 57124
rect 111662 57112 111668 57124
rect 111720 57112 111726 57164
rect 114882 57112 114888 57164
rect 114940 57152 114946 57164
rect 115526 57152 115532 57164
rect 114940 57124 115532 57152
rect 114940 57112 114946 57124
rect 115526 57112 115532 57124
rect 115584 57112 115590 57164
rect 115986 57112 115992 57164
rect 116044 57152 116050 57164
rect 116630 57152 116636 57164
rect 116044 57124 116636 57152
rect 116044 57112 116050 57124
rect 116630 57112 116636 57124
rect 116688 57112 116694 57164
rect 117274 57112 117280 57164
rect 117332 57152 117338 57164
rect 118194 57152 118200 57164
rect 117332 57124 118200 57152
rect 117332 57112 117338 57124
rect 118194 57112 118200 57124
rect 118252 57112 118258 57164
rect 119666 57112 119672 57164
rect 119724 57152 119730 57164
rect 120954 57152 120960 57164
rect 119724 57124 120960 57152
rect 119724 57112 119730 57124
rect 120954 57112 120960 57124
rect 121012 57112 121018 57164
rect 125646 57112 125652 57164
rect 125704 57152 125710 57164
rect 130062 57152 130068 57164
rect 125704 57124 130068 57152
rect 125704 57112 125710 57124
rect 130062 57112 130068 57124
rect 130120 57112 130126 57164
rect 193266 57112 193272 57164
rect 193324 57152 193330 57164
rect 194094 57152 194100 57164
rect 193324 57124 194100 57152
rect 193324 57112 193330 57124
rect 194094 57112 194100 57124
rect 194152 57112 194158 57164
rect 194922 57112 194928 57164
rect 194980 57152 194986 57164
rect 195658 57152 195664 57164
rect 194980 57124 195664 57152
rect 194980 57112 194986 57124
rect 195658 57112 195664 57124
rect 195716 57112 195722 57164
rect 196302 57112 196308 57164
rect 196360 57152 196366 57164
rect 197222 57152 197228 57164
rect 196360 57124 197228 57152
rect 196360 57112 196366 57124
rect 197222 57112 197228 57124
rect 197280 57112 197286 57164
rect 200810 57112 200816 57164
rect 200868 57152 200874 57164
rect 201914 57152 201920 57164
rect 200868 57124 201920 57152
rect 200868 57112 200874 57124
rect 201914 57112 201920 57124
rect 201972 57112 201978 57164
rect 202098 57112 202104 57164
rect 202156 57152 202162 57164
rect 203018 57152 203024 57164
rect 202156 57124 203024 57152
rect 202156 57112 202162 57124
rect 203018 57112 203024 57124
rect 203076 57112 203082 57164
rect 204030 57112 204036 57164
rect 204088 57152 204094 57164
rect 205134 57152 205140 57164
rect 204088 57124 205140 57152
rect 204088 57112 204094 57124
rect 205134 57112 205140 57124
rect 205192 57112 205198 57164
rect 206054 57112 206060 57164
rect 206112 57152 206118 57164
rect 207158 57152 207164 57164
rect 206112 57124 207164 57152
rect 206112 57112 206118 57124
rect 207158 57112 207164 57124
rect 207216 57112 207222 57164
rect 32082 56772 32088 56824
rect 32140 56772 32146 56824
rect 138158 55684 138164 55736
rect 138216 55724 138222 55736
rect 138342 55724 138348 55736
rect 138216 55696 138348 55724
rect 138216 55684 138222 55696
rect 138342 55684 138348 55696
rect 138400 55684 138406 55736
rect 194186 54324 194192 54376
rect 194244 54364 194250 54376
rect 194738 54364 194744 54376
rect 194244 54336 194744 54364
rect 194244 54324 194250 54336
rect 194738 54324 194744 54336
rect 194796 54324 194802 54376
rect 198970 54324 198976 54376
rect 199028 54364 199034 54376
rect 199246 54364 199252 54376
rect 199028 54336 199252 54364
rect 199028 54324 199034 54336
rect 199246 54324 199252 54336
rect 199304 54324 199310 54376
rect 210654 50516 210660 50568
rect 210712 50556 210718 50568
rect 210930 50556 210936 50568
rect 210712 50528 210936 50556
rect 210712 50516 210718 50528
rect 210930 50516 210936 50528
rect 210988 50516 210994 50568
rect 127210 50380 127216 50432
rect 127268 50420 127274 50432
rect 127854 50420 127860 50432
rect 127268 50392 127860 50420
rect 127268 50380 127274 50392
rect 127854 50380 127860 50392
rect 127912 50380 127918 50432
rect 196210 50380 196216 50432
rect 196268 50420 196274 50432
rect 197038 50420 197044 50432
rect 196268 50392 197044 50420
rect 196268 50380 196274 50392
rect 197038 50380 197044 50392
rect 197096 50380 197102 50432
rect 197682 50380 197688 50432
rect 197740 50420 197746 50432
rect 198142 50420 198148 50432
rect 197740 50392 198148 50420
rect 197740 50380 197746 50392
rect 198142 50380 198148 50392
rect 198200 50380 198206 50432
rect 199062 50380 199068 50432
rect 199120 50420 199126 50432
rect 199798 50420 199804 50432
rect 199120 50392 199804 50420
rect 199120 50380 199126 50392
rect 199798 50380 199804 50392
rect 199856 50380 199862 50432
rect 204490 50380 204496 50432
rect 204548 50420 204554 50432
rect 204950 50420 204956 50432
rect 204548 50392 204956 50420
rect 204548 50380 204554 50392
rect 204950 50380 204956 50392
rect 205008 50380 205014 50432
rect 210010 50380 210016 50432
rect 210068 50420 210074 50432
rect 210654 50420 210660 50432
rect 210068 50392 210660 50420
rect 210068 50380 210074 50392
rect 210654 50380 210660 50392
rect 210712 50380 210718 50432
rect 212126 50312 212132 50364
rect 212184 50312 212190 50364
rect 33462 50244 33468 50296
rect 33520 50284 33526 50296
rect 34290 50284 34296 50296
rect 33520 50256 34296 50284
rect 33520 50244 33526 50256
rect 34290 50244 34296 50256
rect 34348 50244 34354 50296
rect 112306 50244 112312 50296
rect 112364 50284 112370 50296
rect 112490 50284 112496 50296
rect 112364 50256 112496 50284
rect 112364 50244 112370 50256
rect 112490 50244 112496 50256
rect 112548 50244 112554 50296
rect 199062 50244 199068 50296
rect 199120 50284 199126 50296
rect 199246 50284 199252 50296
rect 199120 50256 199252 50284
rect 199120 50244 199126 50256
rect 199246 50244 199252 50256
rect 199304 50244 199310 50296
rect 212144 50284 212172 50312
rect 212144 50256 212264 50284
rect 25642 50176 25648 50228
rect 25700 50216 25706 50228
rect 27850 50216 27856 50228
rect 25700 50188 27856 50216
rect 25700 50176 25706 50188
rect 27850 50176 27856 50188
rect 27908 50176 27914 50228
rect 28310 50176 28316 50228
rect 28368 50216 28374 50228
rect 29138 50216 29144 50228
rect 28368 50188 29144 50216
rect 28368 50176 28374 50188
rect 29138 50176 29144 50188
rect 29196 50176 29202 50228
rect 29690 50176 29696 50228
rect 29748 50216 29754 50228
rect 30426 50216 30432 50228
rect 29748 50188 30432 50216
rect 29748 50176 29754 50188
rect 30426 50176 30432 50188
rect 30484 50176 30490 50228
rect 31070 50176 31076 50228
rect 31128 50216 31134 50228
rect 31806 50216 31812 50228
rect 31128 50188 31812 50216
rect 31128 50176 31134 50188
rect 31806 50176 31812 50188
rect 31864 50176 31870 50228
rect 38246 50176 38252 50228
rect 38304 50216 38310 50228
rect 39258 50216 39264 50228
rect 38304 50188 39264 50216
rect 38304 50176 38310 50188
rect 39258 50176 39264 50188
rect 39316 50176 39322 50228
rect 40914 50176 40920 50228
rect 40972 50216 40978 50228
rect 42018 50216 42024 50228
rect 40972 50188 42024 50216
rect 40972 50176 40978 50188
rect 42018 50176 42024 50188
rect 42076 50176 42082 50228
rect 43766 50176 43772 50228
rect 43824 50216 43830 50228
rect 44686 50216 44692 50228
rect 43824 50188 44692 50216
rect 43824 50176 43830 50188
rect 44686 50176 44692 50188
rect 44744 50176 44750 50228
rect 46434 50176 46440 50228
rect 46492 50216 46498 50228
rect 47446 50216 47452 50228
rect 46492 50188 47452 50216
rect 46492 50176 46498 50188
rect 47446 50176 47452 50188
rect 47504 50176 47510 50228
rect 100254 50176 100260 50228
rect 100312 50216 100318 50228
rect 104762 50216 104768 50228
rect 100312 50188 104768 50216
rect 100312 50176 100318 50188
rect 104762 50176 104768 50188
rect 104820 50176 104826 50228
rect 118194 50176 118200 50228
rect 118252 50216 118258 50228
rect 119298 50216 119304 50228
rect 118252 50188 119304 50216
rect 118252 50176 118258 50188
rect 119298 50176 119304 50188
rect 119356 50176 119362 50228
rect 120954 50176 120960 50228
rect 121012 50216 121018 50228
rect 122610 50216 122616 50228
rect 121012 50188 122616 50216
rect 121012 50176 121018 50188
rect 122610 50176 122616 50188
rect 122668 50176 122674 50228
rect 123714 50176 123720 50228
rect 123772 50216 123778 50228
rect 124818 50216 124824 50228
rect 123772 50188 124824 50216
rect 123772 50176 123778 50188
rect 124818 50176 124824 50188
rect 124876 50176 124882 50228
rect 184434 50176 184440 50228
rect 184492 50216 184498 50228
rect 188206 50216 188212 50228
rect 184492 50188 188212 50216
rect 184492 50176 184498 50188
rect 188206 50176 188212 50188
rect 188264 50176 188270 50228
rect 205318 50176 205324 50228
rect 205376 50216 205382 50228
rect 205870 50216 205876 50228
rect 205376 50188 205876 50216
rect 205376 50176 205382 50188
rect 205870 50176 205876 50188
rect 205928 50176 205934 50228
rect 207986 50176 207992 50228
rect 208044 50216 208050 50228
rect 208722 50216 208728 50228
rect 208044 50188 208728 50216
rect 208044 50176 208050 50188
rect 208722 50176 208728 50188
rect 208780 50176 208786 50228
rect 210746 50176 210752 50228
rect 210804 50216 210810 50228
rect 212126 50216 212132 50228
rect 210804 50188 212132 50216
rect 210804 50176 210810 50188
rect 212126 50176 212132 50188
rect 212184 50176 212190 50228
rect 212236 50216 212264 50256
rect 214426 50216 214432 50228
rect 212236 50188 214432 50216
rect 214426 50176 214432 50188
rect 214484 50176 214490 50228
rect 29046 50108 29052 50160
rect 29104 50148 29110 50160
rect 30702 50148 30708 50160
rect 29104 50120 30708 50148
rect 29104 50108 29110 50120
rect 30702 50108 30708 50120
rect 30760 50108 30766 50160
rect 38154 50108 38160 50160
rect 38212 50148 38218 50160
rect 39994 50148 40000 50160
rect 38212 50120 40000 50148
rect 38212 50108 38218 50120
rect 39994 50108 40000 50120
rect 40052 50108 40058 50160
rect 99334 50108 99340 50160
rect 99392 50148 99398 50160
rect 105866 50148 105872 50160
rect 99392 50120 105872 50148
rect 99392 50108 99398 50120
rect 105866 50108 105872 50120
rect 105924 50108 105930 50160
rect 205226 50108 205232 50160
rect 205284 50148 205290 50160
rect 206422 50148 206428 50160
rect 205284 50120 206428 50148
rect 205284 50108 205290 50120
rect 206422 50108 206428 50120
rect 206480 50108 206486 50160
rect 207894 50108 207900 50160
rect 207952 50148 207958 50160
rect 209274 50148 209280 50160
rect 207952 50120 209280 50148
rect 207952 50108 207958 50120
rect 209274 50108 209280 50120
rect 209332 50108 209338 50160
rect 210930 50108 210936 50160
rect 210988 50148 210994 50160
rect 212678 50148 212684 50160
rect 210988 50120 212684 50148
rect 210988 50108 210994 50120
rect 212678 50108 212684 50120
rect 212736 50108 212742 50160
rect 22238 50040 22244 50092
rect 22296 50080 22302 50092
rect 26654 50080 26660 50092
rect 22296 50052 26660 50080
rect 22296 50040 22302 50052
rect 26654 50040 26660 50052
rect 26712 50040 26718 50092
rect 37510 50040 37516 50092
rect 37568 50080 37574 50092
rect 38246 50080 38252 50092
rect 37568 50052 38252 50080
rect 37568 50040 37574 50052
rect 38246 50040 38252 50052
rect 38304 50040 38310 50092
rect 99518 50040 99524 50092
rect 99576 50080 99582 50092
rect 106418 50080 106424 50092
rect 99576 50052 106424 50080
rect 99576 50040 99582 50052
rect 106418 50040 106424 50052
rect 106476 50040 106482 50092
rect 121138 50040 121144 50092
rect 121196 50080 121202 50092
rect 123162 50080 123168 50092
rect 121196 50052 123168 50080
rect 121196 50040 121202 50052
rect 123162 50040 123168 50052
rect 123220 50040 123226 50092
rect 202374 50040 202380 50092
rect 202432 50080 202438 50092
rect 203570 50080 203576 50092
rect 202432 50052 203576 50080
rect 202432 50040 202438 50052
rect 203570 50040 203576 50052
rect 203628 50040 203634 50092
rect 205134 50040 205140 50092
rect 205192 50080 205198 50092
rect 206974 50080 206980 50092
rect 205192 50052 206980 50080
rect 205192 50040 205198 50052
rect 206974 50040 206980 50052
rect 207032 50040 207038 50092
rect 21502 49972 21508 50024
rect 21560 50012 21566 50024
rect 26930 50012 26936 50024
rect 21560 49984 26936 50012
rect 21560 49972 21566 49984
rect 26930 49972 26936 49984
rect 26988 49972 26994 50024
rect 125186 49904 125192 49956
rect 125244 49944 125250 49956
rect 126014 49944 126020 49956
rect 125244 49916 126020 49944
rect 125244 49904 125250 49916
rect 126014 49904 126020 49916
rect 126072 49904 126078 49956
rect 20858 49836 20864 49888
rect 20916 49876 20922 49888
rect 25090 49876 25096 49888
rect 20916 49848 25096 49876
rect 20916 49836 20922 49848
rect 25090 49836 25096 49848
rect 25148 49836 25154 49888
rect 26470 49876 26476 49888
rect 25200 49848 26476 49876
rect 23618 49700 23624 49752
rect 23676 49740 23682 49752
rect 25200 49740 25228 49848
rect 26470 49836 26476 49848
rect 26528 49836 26534 49888
rect 27942 49808 27948 49820
rect 23676 49712 25228 49740
rect 25292 49780 27948 49808
rect 23676 49700 23682 49712
rect 24262 49632 24268 49684
rect 24320 49672 24326 49684
rect 25292 49672 25320 49780
rect 27942 49768 27948 49780
rect 28000 49768 28006 49820
rect 43674 49768 43680 49820
rect 43732 49808 43738 49820
rect 45422 49808 45428 49820
rect 43732 49780 45428 49808
rect 43732 49768 43738 49780
rect 45422 49768 45428 49780
rect 45480 49768 45486 49820
rect 99242 49768 99248 49820
rect 99300 49808 99306 49820
rect 106970 49808 106976 49820
rect 99300 49780 106976 49808
rect 99300 49768 99306 49780
rect 106970 49768 106976 49780
rect 107028 49768 107034 49820
rect 26286 49700 26292 49752
rect 26344 49740 26350 49752
rect 29506 49740 29512 49752
rect 26344 49712 29512 49740
rect 26344 49700 26350 49712
rect 29506 49700 29512 49712
rect 29564 49700 29570 49752
rect 121046 49700 121052 49752
rect 121104 49740 121110 49752
rect 122058 49740 122064 49752
rect 121104 49712 122064 49740
rect 121104 49700 121110 49712
rect 122058 49700 122064 49712
rect 122116 49700 122122 49752
rect 24320 49644 25320 49672
rect 24320 49632 24326 49644
rect 99150 49632 99156 49684
rect 99208 49672 99214 49684
rect 107522 49672 107528 49684
rect 99208 49644 107528 49672
rect 99208 49632 99214 49644
rect 107522 49632 107528 49644
rect 107580 49632 107586 49684
rect 183238 49632 183244 49684
rect 183296 49672 183302 49684
rect 191058 49672 191064 49684
rect 183296 49644 191064 49672
rect 183296 49632 183302 49644
rect 191058 49632 191064 49644
rect 191116 49632 191122 49684
rect 212218 49632 212224 49684
rect 212276 49672 212282 49684
rect 213874 49672 213880 49684
rect 212276 49644 213880 49672
rect 212276 49632 212282 49644
rect 213874 49632 213880 49644
rect 213932 49632 213938 49684
rect 99058 49564 99064 49616
rect 99116 49604 99122 49616
rect 108074 49604 108080 49616
rect 99116 49576 108080 49604
rect 99116 49564 99122 49576
rect 108074 49564 108080 49576
rect 108132 49564 108138 49616
rect 183054 49564 183060 49616
rect 183112 49604 183118 49616
rect 192162 49604 192168 49616
rect 183112 49576 192168 49604
rect 183112 49564 183118 49576
rect 192162 49564 192168 49576
rect 192220 49564 192226 49616
rect 215530 49604 215536 49616
rect 210764 49576 215536 49604
rect 20214 49496 20220 49548
rect 20272 49536 20278 49548
rect 44410 49536 44416 49548
rect 20272 49508 44416 49536
rect 20272 49496 20278 49508
rect 44410 49496 44416 49508
rect 44468 49496 44474 49548
rect 98966 49496 98972 49548
rect 99024 49536 99030 49548
rect 108626 49536 108632 49548
rect 99024 49508 108632 49536
rect 99024 49496 99030 49508
rect 108626 49496 108632 49508
rect 108684 49496 108690 49548
rect 125094 49496 125100 49548
rect 125152 49536 125158 49548
rect 126566 49536 126572 49548
rect 125152 49508 126572 49536
rect 125152 49496 125158 49508
rect 126566 49496 126572 49508
rect 126624 49496 126630 49548
rect 183146 49496 183152 49548
rect 183204 49536 183210 49548
rect 191610 49536 191616 49548
rect 183204 49508 191616 49536
rect 183204 49496 183210 49508
rect 191610 49496 191616 49508
rect 191668 49496 191674 49548
rect 191978 49496 191984 49548
rect 192036 49536 192042 49548
rect 210764 49536 210792 49576
rect 215530 49564 215536 49576
rect 215588 49564 215594 49616
rect 192036 49508 210792 49536
rect 192036 49496 192042 49508
rect 210838 49496 210844 49548
rect 210896 49536 210902 49548
rect 211574 49536 211580 49548
rect 210896 49508 211580 49536
rect 210896 49496 210902 49508
rect 211574 49496 211580 49508
rect 211632 49496 211638 49548
rect 212310 49496 212316 49548
rect 212368 49536 212374 49548
rect 214978 49536 214984 49548
rect 212368 49508 214984 49536
rect 212368 49496 212374 49508
rect 214978 49496 214984 49508
rect 215036 49496 215042 49548
rect 24906 49360 24912 49412
rect 24964 49400 24970 49412
rect 28034 49400 28040 49412
rect 24964 49372 28040 49400
rect 24964 49360 24970 49372
rect 28034 49360 28040 49372
rect 28092 49360 28098 49412
rect 183422 49292 183428 49344
rect 183480 49332 183486 49344
rect 189310 49332 189316 49344
rect 183480 49304 189316 49332
rect 183480 49292 183486 49304
rect 189310 49292 189316 49304
rect 189368 49292 189374 49344
rect 22882 49224 22888 49276
rect 22940 49264 22946 49276
rect 26562 49264 26568 49276
rect 22940 49236 26568 49264
rect 22940 49224 22946 49236
rect 26562 49224 26568 49236
rect 26620 49224 26626 49276
rect 27666 49224 27672 49276
rect 27724 49264 27730 49276
rect 29414 49264 29420 49276
rect 27724 49236 29420 49264
rect 27724 49224 27730 49236
rect 29414 49224 29420 49236
rect 29472 49224 29478 49276
rect 183606 49224 183612 49276
rect 183664 49264 183670 49276
rect 189862 49264 189868 49276
rect 183664 49236 189868 49264
rect 183664 49224 183670 49236
rect 189862 49224 189868 49236
rect 189920 49224 189926 49276
rect 125278 49156 125284 49208
rect 125336 49196 125342 49208
rect 127118 49196 127124 49208
rect 125336 49168 127124 49196
rect 125336 49156 125342 49168
rect 127118 49156 127124 49168
rect 127176 49156 127182 49208
rect 207158 49156 207164 49208
rect 207216 49196 207222 49208
rect 209826 49196 209832 49208
rect 207216 49168 209832 49196
rect 207216 49156 207222 49168
rect 209826 49156 209832 49168
rect 209884 49156 209890 49208
rect 118838 49088 118844 49140
rect 118896 49128 118902 49140
rect 119850 49128 119856 49140
rect 118896 49100 119856 49128
rect 118896 49088 118902 49100
rect 119850 49088 119856 49100
rect 119908 49088 119914 49140
rect 183330 49088 183336 49140
rect 183388 49128 183394 49140
rect 190414 49128 190420 49140
rect 183388 49100 190420 49128
rect 183388 49088 183394 49100
rect 190414 49088 190420 49100
rect 190472 49088 190478 49140
rect 203018 49088 203024 49140
rect 203076 49128 203082 49140
rect 204122 49128 204128 49140
rect 203076 49100 204128 49128
rect 203076 49088 203082 49100
rect 204122 49088 204128 49100
rect 204180 49088 204186 49140
rect 27022 49020 27028 49072
rect 27080 49060 27086 49072
rect 29322 49060 29328 49072
rect 27080 49032 29328 49060
rect 27080 49020 27086 49032
rect 29322 49020 29328 49032
rect 29380 49020 29386 49072
rect 36130 48884 36136 48936
rect 36188 48924 36194 48936
rect 37234 48924 37240 48936
rect 36188 48896 37240 48924
rect 36188 48884 36194 48896
rect 37234 48884 37240 48896
rect 37292 48884 37298 48936
rect 90686 48884 90692 48936
rect 90744 48924 90750 48936
rect 104210 48924 104216 48936
rect 90744 48896 104216 48924
rect 90744 48884 90750 48896
rect 104210 48884 104216 48896
rect 104268 48884 104274 48936
rect 212034 48816 212040 48868
rect 212092 48856 212098 48868
rect 222246 48856 222252 48868
rect 212092 48828 222252 48856
rect 212092 48816 212098 48828
rect 222246 48816 222252 48828
rect 222304 48816 222310 48868
rect 50390 47048 50396 47100
rect 50448 47088 50454 47100
rect 53334 47088 53340 47100
rect 50448 47060 53340 47088
rect 50448 47048 50454 47060
rect 53334 47048 53340 47060
rect 53392 47048 53398 47100
rect 110742 46912 110748 46964
rect 110800 46952 110806 46964
rect 110926 46952 110932 46964
rect 110800 46924 110932 46952
rect 110800 46912 110806 46924
rect 110926 46912 110932 46924
rect 110984 46912 110990 46964
rect 134570 46504 134576 46556
rect 134628 46544 134634 46556
rect 145334 46544 145340 46556
rect 134628 46516 145340 46544
rect 134628 46504 134634 46516
rect 145334 46504 145340 46516
rect 145392 46504 145398 46556
rect 50574 46436 50580 46488
rect 50632 46476 50638 46488
rect 61338 46476 61344 46488
rect 50632 46448 61344 46476
rect 50632 46436 50638 46448
rect 61338 46436 61344 46448
rect 61396 46436 61402 46488
rect 134754 46436 134760 46488
rect 134812 46476 134818 46488
rect 142574 46476 142580 46488
rect 134812 46448 142580 46476
rect 134812 46436 134818 46448
rect 142574 46436 142580 46448
rect 142632 46436 142638 46488
rect 50758 46368 50764 46420
rect 50816 46408 50822 46420
rect 62810 46408 62816 46420
rect 50816 46380 62816 46408
rect 50816 46368 50822 46380
rect 62810 46368 62816 46380
rect 62868 46368 62874 46420
rect 135214 46368 135220 46420
rect 135272 46408 135278 46420
rect 146806 46408 146812 46420
rect 135272 46380 146812 46408
rect 135272 46368 135278 46380
rect 146806 46368 146812 46380
rect 146864 46368 146870 46420
rect 50850 46300 50856 46352
rect 50908 46340 50914 46352
rect 64282 46340 64288 46352
rect 50908 46312 64288 46340
rect 50908 46300 50914 46312
rect 64282 46300 64288 46312
rect 64340 46300 64346 46352
rect 135030 46300 135036 46352
rect 135088 46340 135094 46352
rect 148278 46340 148284 46352
rect 135088 46312 148284 46340
rect 135088 46300 135094 46312
rect 148278 46300 148284 46312
rect 148336 46300 148342 46352
rect 51034 46232 51040 46284
rect 51092 46272 51098 46284
rect 65754 46272 65760 46284
rect 51092 46244 65760 46272
rect 51092 46232 51098 46244
rect 65754 46232 65760 46244
rect 65812 46232 65818 46284
rect 82958 46232 82964 46284
rect 83016 46272 83022 46284
rect 93354 46272 93360 46284
rect 83016 46244 93360 46272
rect 83016 46232 83022 46244
rect 93354 46232 93360 46244
rect 93412 46232 93418 46284
rect 134938 46232 134944 46284
rect 134996 46272 135002 46284
rect 149750 46272 149756 46284
rect 134996 46244 149756 46272
rect 134996 46232 135002 46244
rect 149750 46232 149756 46244
rect 149808 46232 149814 46284
rect 50666 46164 50672 46216
rect 50724 46204 50730 46216
rect 67318 46204 67324 46216
rect 50724 46176 67324 46204
rect 50724 46164 50730 46176
rect 67318 46164 67324 46176
rect 67376 46164 67382 46216
rect 84062 46164 84068 46216
rect 84120 46204 84126 46216
rect 94734 46204 94740 46216
rect 84120 46176 94740 46204
rect 84120 46164 84126 46176
rect 94734 46164 94740 46176
rect 94792 46164 94798 46216
rect 135122 46164 135128 46216
rect 135180 46204 135186 46216
rect 151314 46204 151320 46216
rect 135180 46176 151320 46204
rect 135180 46164 135186 46176
rect 151314 46164 151320 46176
rect 151372 46164 151378 46216
rect 168426 46164 168432 46216
rect 168484 46204 168490 46216
rect 177534 46204 177540 46216
rect 168484 46176 177540 46204
rect 168484 46164 168490 46176
rect 177534 46164 177540 46176
rect 177592 46164 177598 46216
rect 50942 46096 50948 46148
rect 51000 46136 51006 46148
rect 68790 46136 68796 46148
rect 51000 46108 68796 46136
rect 51000 46096 51006 46108
rect 68790 46096 68796 46108
rect 68848 46096 68854 46148
rect 88938 46096 88944 46148
rect 88996 46136 89002 46148
rect 96114 46136 96120 46148
rect 88996 46108 96120 46136
rect 88996 46096 89002 46108
rect 96114 46096 96120 46108
rect 96172 46096 96178 46148
rect 135306 46096 135312 46148
rect 135364 46136 135370 46148
rect 152786 46136 152792 46148
rect 135364 46108 152792 46136
rect 135364 46096 135370 46108
rect 152786 46096 152792 46108
rect 152844 46096 152850 46148
rect 166954 46096 166960 46148
rect 167012 46136 167018 46148
rect 176154 46136 176160 46148
rect 167012 46108 176160 46136
rect 167012 46096 167018 46108
rect 176154 46096 176160 46108
rect 176212 46096 176218 46148
rect 181030 45280 181036 45332
rect 181088 45320 181094 45332
rect 185170 45320 185176 45332
rect 181088 45292 185176 45320
rect 181088 45280 181094 45292
rect 185170 45280 185176 45292
rect 185228 45280 185234 45332
rect 134754 44872 134760 44924
rect 134812 44912 134818 44924
rect 142666 44912 142672 44924
rect 134812 44884 142672 44912
rect 134812 44872 134818 44884
rect 142666 44872 142672 44884
rect 142724 44872 142730 44924
rect 134294 44804 134300 44856
rect 134352 44844 134358 44856
rect 142482 44844 142488 44856
rect 134352 44816 142488 44844
rect 134352 44804 134358 44816
rect 142482 44804 142488 44816
rect 142540 44804 142546 44856
rect 51218 44736 51224 44788
rect 51276 44776 51282 44788
rect 51276 44748 51356 44776
rect 51276 44736 51282 44748
rect 51328 44708 51356 44748
rect 134846 44736 134852 44788
rect 134904 44776 134910 44788
rect 134904 44748 135536 44776
rect 134904 44736 134910 44748
rect 58302 44708 58308 44720
rect 51328 44680 58308 44708
rect 58302 44668 58308 44680
rect 58360 44668 58366 44720
rect 93906 44668 93912 44720
rect 93964 44708 93970 44720
rect 100990 44708 100996 44720
rect 93964 44680 100996 44708
rect 93964 44668 93970 44680
rect 100990 44668 100996 44680
rect 101048 44668 101054 44720
rect 135508 44708 135536 44748
rect 142390 44708 142396 44720
rect 135508 44680 142396 44708
rect 142390 44668 142396 44680
rect 142448 44668 142454 44720
rect 177718 44668 177724 44720
rect 177776 44708 177782 44720
rect 185814 44708 185820 44720
rect 177776 44680 185820 44708
rect 177776 44668 177782 44680
rect 185814 44668 185820 44680
rect 185872 44668 185878 44720
rect 51310 44600 51316 44652
rect 51368 44640 51374 44652
rect 58210 44640 58216 44652
rect 51368 44612 58216 44640
rect 51368 44600 51374 44612
rect 58210 44600 58216 44612
rect 58268 44600 58274 44652
rect 93998 44600 94004 44652
rect 94056 44640 94062 44652
rect 101174 44640 101180 44652
rect 94056 44612 101180 44640
rect 94056 44600 94062 44612
rect 101174 44600 101180 44612
rect 101232 44600 101238 44652
rect 90318 44532 90324 44584
rect 90376 44572 90382 44584
rect 90597 44575 90655 44581
rect 90597 44572 90609 44575
rect 90376 44544 90609 44572
rect 90376 44532 90382 44544
rect 90597 44541 90609 44544
rect 90643 44541 90655 44575
rect 90597 44535 90655 44541
rect 90410 44464 90416 44516
rect 90468 44504 90474 44516
rect 90686 44504 90692 44516
rect 90468 44476 90692 44504
rect 90468 44464 90474 44476
rect 90686 44464 90692 44476
rect 90744 44464 90750 44516
rect 177718 43852 177724 43904
rect 177776 43892 177782 43904
rect 181030 43892 181036 43904
rect 177776 43864 181036 43892
rect 177776 43852 177782 43864
rect 181030 43852 181036 43864
rect 181088 43852 181094 43904
rect 134754 43648 134760 43700
rect 134812 43688 134818 43700
rect 139630 43688 139636 43700
rect 134812 43660 139636 43688
rect 134812 43648 134818 43660
rect 139630 43648 139636 43660
rect 139688 43648 139694 43700
rect 50022 43512 50028 43564
rect 50080 43552 50086 43564
rect 56738 43552 56744 43564
rect 50080 43524 56744 43552
rect 50080 43512 50086 43524
rect 56738 43512 56744 43524
rect 56796 43512 56802 43564
rect 51218 43308 51224 43360
rect 51276 43348 51282 43360
rect 56646 43348 56652 43360
rect 51276 43320 56652 43348
rect 51276 43308 51282 43320
rect 56646 43308 56652 43320
rect 56704 43308 56710 43360
rect 96850 43308 96856 43360
rect 96908 43348 96914 43360
rect 100990 43348 100996 43360
rect 96908 43320 100996 43348
rect 96908 43308 96914 43320
rect 100990 43308 100996 43320
rect 101048 43308 101054 43360
rect 134754 43308 134760 43360
rect 134812 43348 134818 43360
rect 143494 43348 143500 43360
rect 134812 43320 143500 43348
rect 134812 43308 134818 43320
rect 143494 43308 143500 43320
rect 143552 43308 143558 43360
rect 181766 43308 181772 43360
rect 181824 43348 181830 43360
rect 185170 43348 185176 43360
rect 181824 43320 185176 43348
rect 181824 43308 181830 43320
rect 185170 43308 185176 43320
rect 185228 43308 185234 43360
rect 93906 43240 93912 43292
rect 93964 43280 93970 43292
rect 101082 43280 101088 43292
rect 93964 43252 101088 43280
rect 93964 43240 93970 43252
rect 101082 43240 101088 43252
rect 101140 43240 101146 43292
rect 134938 43240 134944 43292
rect 134996 43280 135002 43292
rect 135214 43280 135220 43292
rect 134996 43252 135220 43280
rect 134996 43240 135002 43252
rect 135214 43240 135220 43252
rect 135272 43240 135278 43292
rect 139630 43240 139636 43292
rect 139688 43280 139694 43292
rect 143126 43280 143132 43292
rect 139688 43252 143132 43280
rect 139688 43240 139694 43252
rect 143126 43240 143132 43252
rect 143184 43240 143190 43292
rect 177718 43240 177724 43292
rect 177776 43280 177782 43292
rect 185446 43280 185452 43292
rect 177776 43252 185452 43280
rect 177776 43240 177782 43252
rect 185446 43240 185452 43252
rect 185504 43240 185510 43292
rect 56646 43172 56652 43224
rect 56704 43212 56710 43224
rect 58210 43212 58216 43224
rect 56704 43184 58216 43212
rect 56704 43172 56710 43184
rect 58210 43172 58216 43184
rect 58268 43172 58274 43224
rect 93998 43172 94004 43224
rect 94056 43212 94062 43224
rect 101266 43212 101272 43224
rect 94056 43184 101272 43212
rect 94056 43172 94062 43184
rect 101266 43172 101272 43184
rect 101324 43172 101330 43224
rect 177626 43172 177632 43224
rect 177684 43212 177690 43224
rect 185538 43212 185544 43224
rect 177684 43184 185544 43212
rect 177684 43172 177690 43184
rect 185538 43172 185544 43184
rect 185596 43172 185602 43224
rect 56738 43104 56744 43156
rect 56796 43144 56802 43156
rect 58302 43144 58308 43156
rect 56796 43116 58308 43144
rect 56796 43104 56802 43116
rect 58302 43104 58308 43116
rect 58360 43104 58366 43156
rect 50206 42560 50212 42612
rect 50264 42600 50270 42612
rect 58210 42600 58216 42612
rect 50264 42572 58216 42600
rect 50264 42560 50270 42572
rect 58210 42560 58216 42572
rect 58268 42560 58274 42612
rect 93998 42560 94004 42612
rect 94056 42600 94062 42612
rect 96850 42600 96856 42612
rect 94056 42572 96856 42600
rect 94056 42560 94062 42572
rect 96850 42560 96856 42572
rect 96908 42560 96914 42612
rect 177718 42424 177724 42476
rect 177776 42464 177782 42476
rect 181766 42464 181772 42476
rect 177776 42436 181772 42464
rect 177776 42424 177782 42436
rect 181766 42424 181772 42436
rect 181824 42424 181830 42476
rect 134754 42288 134760 42340
rect 134812 42328 134818 42340
rect 139630 42328 139636 42340
rect 134812 42300 139636 42328
rect 134812 42288 134818 42300
rect 139630 42288 139636 42300
rect 139688 42288 139694 42340
rect 51126 42016 51132 42068
rect 51184 42056 51190 42068
rect 51184 42028 56784 42056
rect 51184 42016 51190 42028
rect 51218 41948 51224 42000
rect 51276 41988 51282 42000
rect 51276 41960 56692 41988
rect 51276 41948 51282 41960
rect 56664 41784 56692 41960
rect 56756 41920 56784 42028
rect 134754 41948 134760 42000
rect 134812 41988 134818 42000
rect 143678 41988 143684 42000
rect 134812 41960 143684 41988
rect 134812 41948 134818 41960
rect 143678 41948 143684 41960
rect 143736 41948 143742 42000
rect 58210 41920 58216 41932
rect 56756 41892 58216 41920
rect 58210 41880 58216 41892
rect 58268 41880 58274 41932
rect 92710 41880 92716 41932
rect 92768 41920 92774 41932
rect 100990 41920 100996 41932
rect 92768 41892 100996 41920
rect 92768 41880 92774 41892
rect 100990 41880 100996 41892
rect 101048 41880 101054 41932
rect 177626 41880 177632 41932
rect 177684 41920 177690 41932
rect 185170 41920 185176 41932
rect 177684 41892 185176 41920
rect 177684 41880 177690 41892
rect 185170 41880 185176 41892
rect 185228 41880 185234 41932
rect 93998 41812 94004 41864
rect 94056 41852 94062 41864
rect 100806 41852 100812 41864
rect 94056 41824 100812 41852
rect 94056 41812 94062 41824
rect 100806 41812 100812 41824
rect 100864 41812 100870 41864
rect 177718 41812 177724 41864
rect 177776 41852 177782 41864
rect 184986 41852 184992 41864
rect 177776 41824 184992 41852
rect 177776 41812 177782 41824
rect 184986 41812 184992 41824
rect 185044 41812 185050 41864
rect 58302 41784 58308 41796
rect 56664 41756 58308 41784
rect 58302 41744 58308 41756
rect 58360 41744 58366 41796
rect 139630 41744 139636 41796
rect 139688 41784 139694 41796
rect 142758 41784 142764 41796
rect 139688 41756 142764 41784
rect 139688 41744 139694 41756
rect 142758 41744 142764 41756
rect 142816 41744 142822 41796
rect 134754 40792 134760 40844
rect 134812 40832 134818 40844
rect 139630 40832 139636 40844
rect 134812 40804 139636 40832
rect 134812 40792 134818 40804
rect 139630 40792 139636 40804
rect 139688 40792 139694 40844
rect 51218 40656 51224 40708
rect 51276 40696 51282 40708
rect 55726 40696 55732 40708
rect 51276 40668 55732 40696
rect 51276 40656 51282 40668
rect 55726 40656 55732 40668
rect 55784 40656 55790 40708
rect 134570 40656 134576 40708
rect 134628 40696 134634 40708
rect 134754 40696 134760 40708
rect 134628 40668 134760 40696
rect 134628 40656 134634 40668
rect 134754 40656 134760 40668
rect 134812 40656 134818 40708
rect 137977 40699 138035 40705
rect 137977 40665 137989 40699
rect 138023 40696 138035 40699
rect 138066 40696 138072 40708
rect 138023 40668 138072 40696
rect 138023 40665 138035 40668
rect 137977 40659 138035 40665
rect 138066 40656 138072 40668
rect 138124 40656 138130 40708
rect 51126 40588 51132 40640
rect 51184 40628 51190 40640
rect 56554 40628 56560 40640
rect 51184 40600 56560 40628
rect 51184 40588 51190 40600
rect 56554 40588 56560 40600
rect 56612 40588 56618 40640
rect 134662 40588 134668 40640
rect 134720 40628 134726 40640
rect 134720 40600 139676 40628
rect 134720 40588 134726 40600
rect 92710 40520 92716 40572
rect 92768 40560 92774 40572
rect 100990 40560 100996 40572
rect 92768 40532 100996 40560
rect 92768 40520 92774 40532
rect 100990 40520 100996 40532
rect 101048 40520 101054 40572
rect 137974 40560 137980 40572
rect 137935 40532 137980 40560
rect 137974 40520 137980 40532
rect 138032 40520 138038 40572
rect 139648 40560 139676 40600
rect 142390 40560 142396 40572
rect 139648 40532 142396 40560
rect 142390 40520 142396 40532
rect 142448 40520 142454 40572
rect 177258 40520 177264 40572
rect 177316 40560 177322 40572
rect 185170 40560 185176 40572
rect 177316 40532 185176 40560
rect 177316 40520 177322 40532
rect 185170 40520 185176 40532
rect 185228 40520 185234 40572
rect 93998 40452 94004 40504
rect 94056 40492 94062 40504
rect 100898 40492 100904 40504
rect 94056 40464 100904 40492
rect 94056 40452 94062 40464
rect 100898 40452 100904 40464
rect 100956 40452 100962 40504
rect 177718 40452 177724 40504
rect 177776 40492 177782 40504
rect 185078 40492 185084 40504
rect 177776 40464 185084 40492
rect 177776 40452 177782 40464
rect 185078 40452 185084 40464
rect 185136 40452 185142 40504
rect 56554 40384 56560 40436
rect 56612 40424 56618 40436
rect 58210 40424 58216 40436
rect 56612 40396 58216 40424
rect 56612 40384 56618 40396
rect 58210 40384 58216 40396
rect 58268 40384 58274 40436
rect 55726 40112 55732 40164
rect 55784 40152 55790 40164
rect 58302 40152 58308 40164
rect 55784 40124 58308 40152
rect 55784 40112 55790 40124
rect 58302 40112 58308 40124
rect 58360 40112 58366 40164
rect 51126 39228 51132 39280
rect 51184 39268 51190 39280
rect 51184 39240 56784 39268
rect 51184 39228 51190 39240
rect 13314 39160 13320 39212
rect 13372 39200 13378 39212
rect 18098 39200 18104 39212
rect 13372 39172 18104 39200
rect 13372 39160 13378 39172
rect 18098 39160 18104 39172
rect 18156 39160 18162 39212
rect 51218 39160 51224 39212
rect 51276 39200 51282 39212
rect 51276 39172 56692 39200
rect 51276 39160 51282 39172
rect 56664 39064 56692 39172
rect 56756 39132 56784 39240
rect 134570 39228 134576 39280
rect 134628 39268 134634 39280
rect 134628 39240 140964 39268
rect 134628 39228 134634 39240
rect 134662 39160 134668 39212
rect 134720 39200 134726 39212
rect 134720 39172 139584 39200
rect 134720 39160 134726 39172
rect 58210 39132 58216 39144
rect 56756 39104 58216 39132
rect 58210 39092 58216 39104
rect 58268 39092 58274 39144
rect 92894 39092 92900 39144
rect 92952 39132 92958 39144
rect 100990 39132 100996 39144
rect 92952 39104 100996 39132
rect 92952 39092 92958 39104
rect 100990 39092 100996 39104
rect 101048 39092 101054 39144
rect 58394 39064 58400 39076
rect 56664 39036 58400 39064
rect 58394 39024 58400 39036
rect 58452 39024 58458 39076
rect 93906 39024 93912 39076
rect 93964 39064 93970 39076
rect 101082 39064 101088 39076
rect 93964 39036 101088 39064
rect 93964 39024 93970 39036
rect 101082 39024 101088 39036
rect 101140 39024 101146 39076
rect 93998 38956 94004 39008
rect 94056 38996 94062 39008
rect 100806 38996 100812 39008
rect 94056 38968 100812 38996
rect 94056 38956 94062 38968
rect 100806 38956 100812 38968
rect 100864 38956 100870 39008
rect 139556 38996 139584 39172
rect 140936 39132 140964 39240
rect 142390 39132 142396 39144
rect 140936 39104 142396 39132
rect 142390 39092 142396 39104
rect 142448 39092 142454 39144
rect 177350 39092 177356 39144
rect 177408 39132 177414 39144
rect 185170 39132 185176 39144
rect 177408 39104 185176 39132
rect 177408 39092 177414 39104
rect 185170 39092 185176 39104
rect 185228 39092 185234 39144
rect 139630 39024 139636 39076
rect 139688 39064 139694 39076
rect 142482 39064 142488 39076
rect 139688 39036 142488 39064
rect 139688 39024 139694 39036
rect 142482 39024 142488 39036
rect 142540 39024 142546 39076
rect 177442 39024 177448 39076
rect 177500 39064 177506 39076
rect 185262 39064 185268 39076
rect 177500 39036 185268 39064
rect 177500 39024 177506 39036
rect 185262 39024 185268 39036
rect 185320 39024 185326 39076
rect 142574 38996 142580 39008
rect 139556 38968 142580 38996
rect 142574 38956 142580 38968
rect 142632 38956 142638 39008
rect 177718 38956 177724 39008
rect 177776 38996 177782 39008
rect 184986 38996 184992 39008
rect 177776 38968 184992 38996
rect 177776 38956 177782 38968
rect 184986 38956 184992 38968
rect 185044 38956 185050 39008
rect 51218 38412 51224 38464
rect 51276 38452 51282 38464
rect 58302 38452 58308 38464
rect 51276 38424 58308 38452
rect 51276 38412 51282 38424
rect 58302 38412 58308 38424
rect 58360 38412 58366 38464
rect 183698 38140 183704 38192
rect 183756 38180 183762 38192
rect 185262 38180 185268 38192
rect 183756 38152 185268 38180
rect 183756 38140 183762 38152
rect 185262 38140 185268 38152
rect 185320 38140 185326 38192
rect 134662 37936 134668 37988
rect 134720 37976 134726 37988
rect 142574 37976 142580 37988
rect 134720 37948 142580 37976
rect 134720 37936 134726 37948
rect 142574 37936 142580 37948
rect 142632 37936 142638 37988
rect 51126 37868 51132 37920
rect 51184 37908 51190 37920
rect 58394 37908 58400 37920
rect 51184 37880 58400 37908
rect 51184 37868 51190 37880
rect 58394 37868 58400 37880
rect 58452 37868 58458 37920
rect 98230 37868 98236 37920
rect 98288 37908 98294 37920
rect 101082 37908 101088 37920
rect 98288 37880 101088 37908
rect 98288 37868 98294 37880
rect 101082 37868 101088 37880
rect 101140 37868 101146 37920
rect 134294 37868 134300 37920
rect 134352 37908 134358 37920
rect 142482 37908 142488 37920
rect 134352 37880 142488 37908
rect 134352 37868 134358 37880
rect 142482 37868 142488 37880
rect 142540 37868 142546 37920
rect 51218 37800 51224 37852
rect 51276 37840 51282 37852
rect 58210 37840 58216 37852
rect 51276 37812 58216 37840
rect 51276 37800 51282 37812
rect 58210 37800 58216 37812
rect 58268 37800 58274 37852
rect 90594 37840 90600 37852
rect 90555 37812 90600 37840
rect 90594 37800 90600 37812
rect 90652 37800 90658 37852
rect 98322 37800 98328 37852
rect 98380 37840 98386 37852
rect 100990 37840 100996 37852
rect 98380 37812 100996 37840
rect 98380 37800 98386 37812
rect 100990 37800 100996 37812
rect 101048 37800 101054 37852
rect 134110 37800 134116 37852
rect 134168 37840 134174 37852
rect 142390 37840 142396 37852
rect 134168 37812 142396 37840
rect 134168 37800 134174 37812
rect 142390 37800 142396 37812
rect 142448 37800 142454 37852
rect 183238 37800 183244 37852
rect 183296 37840 183302 37852
rect 185170 37840 185176 37852
rect 183296 37812 185176 37840
rect 183296 37800 183302 37812
rect 185170 37800 185176 37812
rect 185228 37800 185234 37852
rect 93998 37596 94004 37648
rect 94056 37636 94062 37648
rect 98230 37636 98236 37648
rect 94056 37608 98236 37636
rect 94056 37596 94062 37608
rect 98230 37596 98236 37608
rect 98288 37596 98294 37648
rect 177442 37324 177448 37376
rect 177500 37364 177506 37376
rect 183698 37364 183704 37376
rect 177500 37336 183704 37364
rect 177500 37324 177506 37336
rect 183698 37324 183704 37336
rect 183756 37324 183762 37376
rect 93998 37052 94004 37104
rect 94056 37092 94062 37104
rect 98322 37092 98328 37104
rect 94056 37064 98328 37092
rect 94056 37052 94062 37064
rect 98322 37052 98328 37064
rect 98380 37052 98386 37104
rect 177718 36848 177724 36900
rect 177776 36888 177782 36900
rect 183238 36888 183244 36900
rect 177776 36860 183244 36888
rect 177776 36848 177782 36860
rect 183238 36848 183244 36860
rect 183296 36848 183302 36900
rect 134386 36576 134392 36628
rect 134444 36616 134450 36628
rect 140918 36616 140924 36628
rect 134444 36588 140924 36616
rect 134444 36576 134450 36588
rect 140918 36576 140924 36588
rect 140976 36576 140982 36628
rect 51218 36508 51224 36560
rect 51276 36548 51282 36560
rect 58302 36548 58308 36560
rect 51276 36520 58308 36548
rect 51276 36508 51282 36520
rect 58302 36508 58308 36520
rect 58360 36508 58366 36560
rect 51126 36440 51132 36492
rect 51184 36480 51190 36492
rect 58210 36480 58216 36492
rect 51184 36452 58216 36480
rect 51184 36440 51190 36452
rect 58210 36440 58216 36452
rect 58268 36440 58274 36492
rect 134662 36440 134668 36492
rect 134720 36480 134726 36492
rect 142390 36480 142396 36492
rect 134720 36452 142396 36480
rect 134720 36440 134726 36452
rect 142390 36440 142396 36452
rect 142448 36440 142454 36492
rect 92894 36372 92900 36424
rect 92952 36412 92958 36424
rect 100990 36412 100996 36424
rect 92952 36384 100996 36412
rect 92952 36372 92958 36384
rect 100990 36372 100996 36384
rect 101048 36372 101054 36424
rect 177350 36372 177356 36424
rect 177408 36412 177414 36424
rect 185170 36412 185176 36424
rect 177408 36384 185176 36412
rect 177408 36372 177414 36384
rect 185170 36372 185176 36384
rect 185228 36372 185234 36424
rect 93998 36304 94004 36356
rect 94056 36344 94062 36356
rect 100806 36344 100812 36356
rect 94056 36316 100812 36344
rect 94056 36304 94062 36316
rect 100806 36304 100812 36316
rect 100864 36304 100870 36356
rect 177718 36304 177724 36356
rect 177776 36344 177782 36356
rect 184986 36344 184992 36356
rect 177776 36316 184992 36344
rect 177776 36304 177782 36316
rect 184986 36304 184992 36316
rect 185044 36304 185050 36356
rect 134662 35624 134668 35676
rect 134720 35664 134726 35676
rect 140182 35664 140188 35676
rect 134720 35636 140188 35664
rect 134720 35624 134726 35636
rect 140182 35624 140188 35636
rect 140240 35624 140246 35676
rect 50022 35216 50028 35268
rect 50080 35256 50086 35268
rect 55450 35256 55456 35268
rect 50080 35228 55456 35256
rect 50080 35216 50086 35228
rect 55450 35216 55456 35228
rect 55508 35216 55514 35268
rect 51218 35080 51224 35132
rect 51276 35120 51282 35132
rect 51276 35092 55496 35120
rect 51276 35080 51282 35092
rect 55468 35052 55496 35092
rect 134110 35080 134116 35132
rect 134168 35120 134174 35132
rect 142482 35120 142488 35132
rect 134168 35092 142488 35120
rect 134168 35080 134174 35092
rect 142482 35080 142488 35092
rect 142540 35080 142546 35132
rect 58302 35052 58308 35064
rect 55468 35024 58308 35052
rect 58302 35012 58308 35024
rect 58360 35012 58366 35064
rect 93446 35012 93452 35064
rect 93504 35052 93510 35064
rect 100990 35052 100996 35064
rect 93504 35024 100996 35052
rect 93504 35012 93510 35024
rect 100990 35012 100996 35024
rect 101048 35012 101054 35064
rect 140918 35012 140924 35064
rect 140976 35052 140982 35064
rect 142574 35052 142580 35064
rect 140976 35024 142580 35052
rect 140976 35012 140982 35024
rect 142574 35012 142580 35024
rect 142632 35012 142638 35064
rect 177626 35012 177632 35064
rect 177684 35052 177690 35064
rect 185446 35052 185452 35064
rect 177684 35024 185452 35052
rect 177684 35012 177690 35024
rect 185446 35012 185452 35024
rect 185504 35012 185510 35064
rect 55450 34944 55456 34996
rect 55508 34984 55514 34996
rect 58210 34984 58216 34996
rect 55508 34956 58216 34984
rect 55508 34944 55514 34956
rect 58210 34944 58216 34956
rect 58268 34944 58274 34996
rect 93998 34944 94004 34996
rect 94056 34984 94062 34996
rect 100898 34984 100904 34996
rect 94056 34956 100904 34984
rect 94056 34944 94062 34956
rect 100898 34944 100904 34956
rect 100956 34944 100962 34996
rect 177718 34944 177724 34996
rect 177776 34984 177782 34996
rect 185078 34984 185084 34996
rect 177776 34956 185084 34984
rect 177776 34944 177782 34956
rect 185078 34944 185084 34956
rect 185136 34944 185142 34996
rect 140182 34876 140188 34928
rect 140240 34916 140246 34928
rect 142390 34916 142396 34928
rect 140240 34888 142396 34916
rect 140240 34876 140246 34888
rect 142390 34876 142396 34888
rect 142448 34876 142454 34928
rect 51218 33992 51224 34044
rect 51276 34032 51282 34044
rect 56738 34032 56744 34044
rect 51276 34004 56744 34032
rect 51276 33992 51282 34004
rect 56738 33992 56744 34004
rect 56796 33992 56802 34044
rect 134662 33992 134668 34044
rect 134720 34032 134726 34044
rect 140182 34032 140188 34044
rect 134720 34004 140188 34032
rect 134720 33992 134726 34004
rect 140182 33992 140188 34004
rect 140240 33992 140246 34044
rect 50206 33720 50212 33772
rect 50264 33760 50270 33772
rect 50264 33732 56784 33760
rect 50264 33720 50270 33732
rect 51218 33652 51224 33704
rect 51276 33692 51282 33704
rect 56002 33692 56008 33704
rect 51276 33664 56008 33692
rect 51276 33652 51282 33664
rect 56002 33652 56008 33664
rect 56060 33652 56066 33704
rect 56756 33624 56784 33732
rect 134662 33720 134668 33772
rect 134720 33760 134726 33772
rect 140918 33760 140924 33772
rect 134720 33732 140924 33760
rect 134720 33720 134726 33732
rect 140918 33720 140924 33732
rect 140976 33720 140982 33772
rect 134570 33652 134576 33704
rect 134628 33692 134634 33704
rect 134628 33664 140780 33692
rect 134628 33652 134634 33664
rect 58210 33624 58216 33636
rect 56756 33596 58216 33624
rect 58210 33584 58216 33596
rect 58268 33584 58274 33636
rect 93814 33584 93820 33636
rect 93872 33624 93878 33636
rect 100990 33624 100996 33636
rect 93872 33596 100996 33624
rect 93872 33584 93878 33596
rect 100990 33584 100996 33596
rect 101048 33584 101054 33636
rect 140752 33624 140780 33664
rect 142390 33624 142396 33636
rect 140752 33596 142396 33624
rect 142390 33584 142396 33596
rect 142448 33584 142454 33636
rect 177810 33584 177816 33636
rect 177868 33624 177874 33636
rect 185170 33624 185176 33636
rect 177868 33596 185176 33624
rect 177868 33584 177874 33596
rect 185170 33584 185176 33596
rect 185228 33584 185234 33636
rect 93998 33516 94004 33568
rect 94056 33556 94062 33568
rect 101082 33556 101088 33568
rect 94056 33528 101088 33556
rect 94056 33516 94062 33528
rect 101082 33516 101088 33528
rect 101140 33516 101146 33568
rect 177718 33516 177724 33568
rect 177776 33556 177782 33568
rect 185262 33556 185268 33568
rect 177776 33528 185268 33556
rect 177776 33516 177782 33528
rect 185262 33516 185268 33528
rect 185320 33516 185326 33568
rect 56738 33448 56744 33500
rect 56796 33488 56802 33500
rect 58210 33488 58216 33500
rect 56796 33460 58216 33488
rect 56796 33448 56802 33460
rect 58210 33448 58216 33460
rect 58268 33448 58274 33500
rect 93906 33448 93912 33500
rect 93964 33488 93970 33500
rect 100714 33488 100720 33500
rect 93964 33460 100720 33488
rect 93964 33448 93970 33460
rect 100714 33448 100720 33460
rect 100772 33448 100778 33500
rect 177626 33448 177632 33500
rect 177684 33488 177690 33500
rect 184894 33488 184900 33500
rect 177684 33460 184900 33488
rect 177684 33448 177690 33460
rect 184894 33448 184900 33460
rect 184952 33448 184958 33500
rect 140182 33176 140188 33228
rect 140240 33216 140246 33228
rect 142390 33216 142396 33228
rect 140240 33188 142396 33216
rect 140240 33176 140246 33188
rect 142390 33176 142396 33188
rect 142448 33176 142454 33228
rect 56002 32972 56008 33024
rect 56060 33012 56066 33024
rect 58210 33012 58216 33024
rect 56060 32984 58216 33012
rect 56060 32972 56066 32984
rect 58210 32972 58216 32984
rect 58268 32972 58274 33024
rect 51218 32360 51224 32412
rect 51276 32400 51282 32412
rect 56738 32400 56744 32412
rect 51276 32372 56744 32400
rect 51276 32360 51282 32372
rect 56738 32360 56744 32372
rect 56796 32360 56802 32412
rect 134386 32360 134392 32412
rect 134444 32400 134450 32412
rect 139722 32400 139728 32412
rect 134444 32372 139728 32400
rect 134444 32360 134450 32372
rect 139722 32360 139728 32372
rect 139780 32360 139786 32412
rect 50022 32292 50028 32344
rect 50080 32332 50086 32344
rect 56646 32332 56652 32344
rect 50080 32304 56652 32332
rect 50080 32292 50086 32304
rect 56646 32292 56652 32304
rect 56704 32292 56710 32344
rect 134294 32292 134300 32344
rect 134352 32332 134358 32344
rect 134352 32304 140964 32332
rect 134352 32292 134358 32304
rect 93906 32224 93912 32276
rect 93964 32264 93970 32276
rect 100990 32264 100996 32276
rect 93964 32236 100996 32264
rect 93964 32224 93970 32236
rect 100990 32224 100996 32236
rect 101048 32224 101054 32276
rect 140936 32264 140964 32304
rect 142390 32264 142396 32276
rect 140936 32236 142396 32264
rect 142390 32224 142396 32236
rect 142448 32224 142454 32276
rect 177718 32224 177724 32276
rect 177776 32264 177782 32276
rect 185170 32264 185176 32276
rect 177776 32236 185176 32264
rect 177776 32224 177782 32236
rect 185170 32224 185176 32236
rect 185228 32224 185234 32276
rect 56646 32156 56652 32208
rect 56704 32196 56710 32208
rect 58210 32196 58216 32208
rect 56704 32168 58216 32196
rect 56704 32156 56710 32168
rect 58210 32156 58216 32168
rect 58268 32156 58274 32208
rect 93998 32156 94004 32208
rect 94056 32196 94062 32208
rect 100806 32196 100812 32208
rect 94056 32168 100812 32196
rect 94056 32156 94062 32168
rect 100806 32156 100812 32168
rect 100864 32156 100870 32208
rect 140918 32156 140924 32208
rect 140976 32196 140982 32208
rect 142482 32196 142488 32208
rect 140976 32168 142488 32196
rect 140976 32156 140982 32168
rect 142482 32156 142488 32168
rect 142540 32156 142546 32208
rect 176982 32156 176988 32208
rect 177040 32196 177046 32208
rect 184986 32196 184992 32208
rect 177040 32168 184992 32196
rect 177040 32156 177046 32168
rect 184986 32156 184992 32168
rect 185044 32156 185050 32208
rect 56738 31816 56744 31868
rect 56796 31856 56802 31868
rect 58302 31856 58308 31868
rect 56796 31828 58308 31856
rect 56796 31816 56802 31828
rect 58302 31816 58308 31828
rect 58360 31816 58366 31868
rect 134662 31272 134668 31324
rect 134720 31312 134726 31324
rect 139630 31312 139636 31324
rect 134720 31284 139636 31312
rect 134720 31272 134726 31284
rect 139630 31272 139636 31284
rect 139688 31272 139694 31324
rect 51126 31000 51132 31052
rect 51184 31040 51190 31052
rect 51184 31012 56784 31040
rect 51184 31000 51190 31012
rect 51218 30932 51224 30984
rect 51276 30972 51282 30984
rect 51276 30944 56692 30972
rect 51276 30932 51282 30944
rect 56664 30768 56692 30944
rect 56756 30904 56784 31012
rect 134662 30932 134668 30984
rect 134720 30972 134726 30984
rect 143586 30972 143592 30984
rect 134720 30944 143592 30972
rect 134720 30932 134726 30944
rect 143586 30932 143592 30944
rect 143644 30932 143650 30984
rect 58210 30904 58216 30916
rect 56756 30876 58216 30904
rect 58210 30864 58216 30876
rect 58268 30864 58274 30916
rect 92710 30864 92716 30916
rect 92768 30904 92774 30916
rect 100990 30904 100996 30916
rect 92768 30876 100996 30904
rect 92768 30864 92774 30876
rect 100990 30864 100996 30876
rect 101048 30864 101054 30916
rect 134386 30864 134392 30916
rect 134444 30904 134450 30916
rect 134846 30904 134852 30916
rect 134444 30876 134852 30904
rect 134444 30864 134450 30876
rect 134846 30864 134852 30876
rect 134904 30864 134910 30916
rect 177166 30864 177172 30916
rect 177224 30904 177230 30916
rect 185170 30904 185176 30916
rect 177224 30876 185176 30904
rect 177224 30864 177230 30876
rect 185170 30864 185176 30876
rect 185228 30864 185234 30916
rect 93998 30796 94004 30848
rect 94056 30836 94062 30848
rect 100898 30836 100904 30848
rect 94056 30808 100904 30836
rect 94056 30796 94062 30808
rect 100898 30796 100904 30808
rect 100956 30796 100962 30848
rect 177442 30796 177448 30848
rect 177500 30836 177506 30848
rect 185078 30836 185084 30848
rect 177500 30808 185084 30836
rect 177500 30796 177506 30808
rect 185078 30796 185084 30808
rect 185136 30796 185142 30848
rect 58302 30768 58308 30780
rect 56664 30740 58308 30768
rect 58302 30728 58308 30740
rect 58360 30728 58366 30780
rect 139722 30728 139728 30780
rect 139780 30768 139786 30780
rect 142390 30768 142396 30780
rect 139780 30740 142396 30768
rect 139780 30728 139786 30740
rect 142390 30728 142396 30740
rect 142448 30728 142454 30780
rect 139630 30524 139636 30576
rect 139688 30564 139694 30576
rect 142390 30564 142396 30576
rect 139688 30536 142396 30564
rect 139688 30524 139694 30536
rect 142390 30524 142396 30536
rect 142448 30524 142454 30576
rect 51126 29572 51132 29624
rect 51184 29612 51190 29624
rect 51184 29584 56784 29612
rect 51184 29572 51190 29584
rect 51218 29504 51224 29556
rect 51276 29544 51282 29556
rect 56646 29544 56652 29556
rect 51276 29516 56652 29544
rect 51276 29504 51282 29516
rect 56646 29504 56652 29516
rect 56704 29504 56710 29556
rect 56756 29476 56784 29584
rect 134754 29572 134760 29624
rect 134812 29612 134818 29624
rect 134812 29584 140964 29612
rect 134812 29572 134818 29584
rect 134202 29504 134208 29556
rect 134260 29544 134266 29556
rect 134260 29516 140872 29544
rect 134260 29504 134266 29516
rect 58210 29476 58216 29488
rect 56756 29448 58216 29476
rect 58210 29436 58216 29448
rect 58268 29436 58274 29488
rect 93906 29436 93912 29488
rect 93964 29476 93970 29488
rect 101082 29476 101088 29488
rect 93964 29448 101088 29476
rect 93964 29436 93970 29448
rect 101082 29436 101088 29448
rect 101140 29436 101146 29488
rect 92710 29368 92716 29420
rect 92768 29408 92774 29420
rect 100990 29408 100996 29420
rect 92768 29380 100996 29408
rect 92768 29368 92774 29380
rect 100990 29368 100996 29380
rect 101048 29368 101054 29420
rect 140844 29408 140872 29516
rect 140936 29476 140964 29584
rect 142390 29476 142396 29488
rect 140936 29448 142396 29476
rect 142390 29436 142396 29448
rect 142448 29436 142454 29488
rect 177810 29436 177816 29488
rect 177868 29476 177874 29488
rect 185262 29476 185268 29488
rect 177868 29448 185268 29476
rect 177868 29436 177874 29448
rect 185262 29436 185268 29448
rect 185320 29436 185326 29488
rect 142482 29408 142488 29420
rect 140844 29380 142488 29408
rect 142482 29368 142488 29380
rect 142540 29368 142546 29420
rect 177626 29368 177632 29420
rect 177684 29408 177690 29420
rect 185170 29408 185176 29420
rect 177684 29380 185176 29408
rect 177684 29368 177690 29380
rect 185170 29368 185176 29380
rect 185228 29368 185234 29420
rect 93998 29300 94004 29352
rect 94056 29340 94062 29352
rect 100806 29340 100812 29352
rect 94056 29312 100812 29340
rect 94056 29300 94062 29312
rect 100806 29300 100812 29312
rect 100864 29300 100870 29352
rect 177718 29300 177724 29352
rect 177776 29340 177782 29352
rect 184986 29340 184992 29352
rect 177776 29312 184992 29340
rect 177776 29300 177782 29312
rect 184986 29300 184992 29312
rect 185044 29300 185050 29352
rect 56646 29232 56652 29284
rect 56704 29272 56710 29284
rect 58210 29272 58216 29284
rect 56704 29244 58216 29272
rect 56704 29232 56710 29244
rect 58210 29232 58216 29244
rect 58268 29232 58274 29284
rect 51126 28756 51132 28808
rect 51184 28796 51190 28808
rect 58210 28796 58216 28808
rect 51184 28768 58216 28796
rect 51184 28756 51190 28768
rect 58210 28756 58216 28768
rect 58268 28756 58274 28808
rect 51218 28552 51224 28604
rect 51276 28592 51282 28604
rect 56738 28592 56744 28604
rect 51276 28564 56744 28592
rect 51276 28552 51282 28564
rect 56738 28552 56744 28564
rect 56796 28552 56802 28604
rect 134754 28416 134760 28468
rect 134812 28456 134818 28468
rect 140274 28456 140280 28468
rect 134812 28428 140280 28456
rect 134812 28416 134818 28428
rect 140274 28416 140280 28428
rect 140332 28416 140338 28468
rect 51218 28280 51224 28332
rect 51276 28320 51282 28332
rect 56002 28320 56008 28332
rect 51276 28292 56008 28320
rect 51276 28280 51282 28292
rect 56002 28280 56008 28292
rect 56060 28280 56066 28332
rect 134754 28212 134760 28264
rect 134812 28252 134818 28264
rect 140918 28252 140924 28264
rect 134812 28224 140924 28252
rect 134812 28212 134818 28224
rect 140918 28212 140924 28224
rect 140976 28212 140982 28264
rect 93906 28144 93912 28196
rect 93964 28184 93970 28196
rect 100990 28184 100996 28196
rect 93964 28156 100996 28184
rect 93964 28144 93970 28156
rect 100990 28144 100996 28156
rect 101048 28144 101054 28196
rect 134570 28144 134576 28196
rect 134628 28184 134634 28196
rect 134628 28156 140964 28184
rect 134628 28144 134634 28156
rect 56738 28076 56744 28128
rect 56796 28116 56802 28128
rect 58210 28116 58216 28128
rect 56796 28088 58216 28116
rect 56796 28076 56802 28088
rect 58210 28076 58216 28088
rect 58268 28076 58274 28128
rect 90686 28116 90692 28128
rect 90647 28088 90692 28116
rect 90686 28076 90692 28088
rect 90744 28076 90750 28128
rect 93998 28076 94004 28128
rect 94056 28116 94062 28128
rect 101174 28116 101180 28128
rect 94056 28088 101180 28116
rect 94056 28076 94062 28088
rect 101174 28076 101180 28088
rect 101232 28076 101238 28128
rect 140936 28116 140964 28156
rect 177442 28144 177448 28196
rect 177500 28184 177506 28196
rect 185170 28184 185176 28196
rect 177500 28156 185176 28184
rect 177500 28144 177506 28156
rect 185170 28144 185176 28156
rect 185228 28144 185234 28196
rect 142390 28116 142396 28128
rect 140936 28088 142396 28116
rect 142390 28076 142396 28088
rect 142448 28076 142454 28128
rect 177718 28076 177724 28128
rect 177776 28116 177782 28128
rect 185354 28116 185360 28128
rect 177776 28088 185360 28116
rect 177776 28076 177782 28088
rect 185354 28076 185360 28088
rect 185412 28076 185418 28128
rect 92710 28008 92716 28060
rect 92768 28048 92774 28060
rect 101082 28048 101088 28060
rect 92768 28020 101088 28048
rect 92768 28008 92774 28020
rect 101082 28008 101088 28020
rect 101140 28008 101146 28060
rect 177258 28008 177264 28060
rect 177316 28048 177322 28060
rect 185262 28048 185268 28060
rect 177316 28020 185268 28048
rect 177316 28008 177322 28020
rect 185262 28008 185268 28020
rect 185320 28008 185326 28060
rect 140274 27736 140280 27788
rect 140332 27776 140338 27788
rect 142390 27776 142396 27788
rect 140332 27748 142396 27776
rect 140332 27736 140338 27748
rect 142390 27736 142396 27748
rect 142448 27736 142454 27788
rect 56002 27668 56008 27720
rect 56060 27708 56066 27720
rect 58302 27708 58308 27720
rect 56060 27680 58308 27708
rect 56060 27668 56066 27680
rect 58302 27668 58308 27680
rect 58360 27668 58366 27720
rect 51218 26852 51224 26904
rect 51276 26892 51282 26904
rect 58302 26892 58308 26904
rect 51276 26864 58308 26892
rect 51276 26852 51282 26864
rect 58302 26852 58308 26864
rect 58360 26852 58366 26904
rect 134754 26852 134760 26904
rect 134812 26892 134818 26904
rect 142574 26892 142580 26904
rect 134812 26864 142580 26892
rect 134812 26852 134818 26864
rect 142574 26852 142580 26864
rect 142632 26852 142638 26904
rect 51126 26784 51132 26836
rect 51184 26824 51190 26836
rect 58210 26824 58216 26836
rect 51184 26796 58216 26824
rect 51184 26784 51190 26796
rect 58210 26784 58216 26796
rect 58268 26784 58274 26836
rect 98230 26784 98236 26836
rect 98288 26824 98294 26836
rect 100990 26824 100996 26836
rect 98288 26796 100996 26824
rect 98288 26784 98294 26796
rect 100990 26784 100996 26796
rect 101048 26784 101054 26836
rect 134570 26784 134576 26836
rect 134628 26824 134634 26836
rect 142390 26824 142396 26836
rect 134628 26796 142396 26824
rect 134628 26784 134634 26796
rect 142390 26784 142396 26796
rect 142448 26784 142454 26836
rect 185170 26824 185176 26836
rect 183716 26796 185176 26824
rect 140918 26716 140924 26768
rect 140976 26756 140982 26768
rect 142482 26756 142488 26768
rect 140976 26728 142488 26756
rect 140976 26716 140982 26728
rect 142482 26716 142488 26728
rect 142540 26716 142546 26768
rect 177718 26716 177724 26768
rect 177776 26756 177782 26768
rect 183716 26756 183744 26796
rect 185170 26784 185176 26796
rect 185228 26784 185234 26836
rect 177776 26728 183744 26756
rect 177776 26716 177782 26728
rect 93998 26308 94004 26360
rect 94056 26348 94062 26360
rect 98230 26348 98236 26360
rect 94056 26320 98236 26348
rect 94056 26308 94062 26320
rect 98230 26308 98236 26320
rect 98288 26308 98294 26360
rect 51126 25560 51132 25612
rect 51184 25600 51190 25612
rect 59314 25600 59320 25612
rect 51184 25572 59320 25600
rect 51184 25560 51190 25572
rect 59314 25560 59320 25572
rect 59372 25560 59378 25612
rect 51218 25492 51224 25544
rect 51276 25532 51282 25544
rect 59406 25532 59412 25544
rect 51276 25504 59412 25532
rect 51276 25492 51282 25504
rect 59406 25492 59412 25504
rect 59464 25492 59470 25544
rect 134754 25492 134760 25544
rect 134812 25532 134818 25544
rect 142482 25532 142488 25544
rect 134812 25504 142488 25532
rect 134812 25492 134818 25504
rect 142482 25492 142488 25504
rect 142540 25492 142546 25544
rect 50482 25424 50488 25476
rect 50540 25464 50546 25476
rect 59498 25464 59504 25476
rect 50540 25436 59504 25464
rect 50540 25424 50546 25436
rect 59498 25424 59504 25436
rect 59556 25424 59562 25476
rect 134570 25424 134576 25476
rect 134628 25464 134634 25476
rect 142390 25464 142396 25476
rect 134628 25436 142396 25464
rect 134628 25424 134634 25436
rect 142390 25424 142396 25436
rect 142448 25424 142454 25476
rect 93814 25356 93820 25408
rect 93872 25396 93878 25408
rect 100990 25396 100996 25408
rect 93872 25368 100996 25396
rect 93872 25356 93878 25368
rect 100990 25356 100996 25368
rect 101048 25356 101054 25408
rect 177350 25356 177356 25408
rect 177408 25396 177414 25408
rect 185446 25396 185452 25408
rect 177408 25368 185452 25396
rect 177408 25356 177414 25368
rect 185446 25356 185452 25368
rect 185504 25356 185510 25408
rect 93906 25288 93912 25340
rect 93964 25328 93970 25340
rect 101082 25328 101088 25340
rect 93964 25300 101088 25328
rect 93964 25288 93970 25300
rect 101082 25288 101088 25300
rect 101140 25288 101146 25340
rect 177718 25288 177724 25340
rect 177776 25328 177782 25340
rect 185354 25328 185360 25340
rect 177776 25300 185360 25328
rect 177776 25288 177782 25300
rect 185354 25288 185360 25300
rect 185412 25288 185418 25340
rect 93998 25220 94004 25272
rect 94056 25260 94062 25272
rect 101174 25260 101180 25272
rect 94056 25232 101180 25260
rect 94056 25220 94062 25232
rect 101174 25220 101180 25232
rect 101232 25220 101238 25272
rect 177626 25220 177632 25272
rect 177684 25260 177690 25272
rect 185538 25260 185544 25272
rect 177684 25232 185544 25260
rect 177684 25220 177690 25232
rect 185538 25220 185544 25232
rect 185596 25220 185602 25272
rect 51126 24064 51132 24116
rect 51184 24104 51190 24116
rect 51184 24076 56784 24104
rect 51184 24064 51190 24076
rect 51218 23996 51224 24048
rect 51276 24036 51282 24048
rect 51276 24008 56692 24036
rect 51276 23996 51282 24008
rect 56664 23900 56692 24008
rect 56756 23968 56784 24076
rect 134570 24064 134576 24116
rect 134628 24104 134634 24116
rect 134628 24076 140964 24104
rect 134628 24064 134634 24076
rect 134754 23996 134760 24048
rect 134812 24036 134818 24048
rect 134812 24008 140872 24036
rect 134812 23996 134818 24008
rect 58210 23968 58216 23980
rect 56756 23940 58216 23968
rect 58210 23928 58216 23940
rect 58268 23928 58274 23980
rect 92894 23928 92900 23980
rect 92952 23968 92958 23980
rect 100990 23968 100996 23980
rect 92952 23940 100996 23968
rect 92952 23928 92958 23940
rect 100990 23928 100996 23940
rect 101048 23928 101054 23980
rect 58302 23900 58308 23912
rect 56664 23872 58308 23900
rect 58302 23860 58308 23872
rect 58360 23860 58366 23912
rect 93998 23860 94004 23912
rect 94056 23900 94062 23912
rect 101082 23900 101088 23912
rect 94056 23872 101088 23900
rect 94056 23860 94062 23872
rect 101082 23860 101088 23872
rect 101140 23860 101146 23912
rect 140844 23900 140872 24008
rect 140936 23968 140964 24076
rect 142390 23968 142396 23980
rect 140936 23940 142396 23968
rect 142390 23928 142396 23940
rect 142448 23928 142454 23980
rect 177534 23928 177540 23980
rect 177592 23968 177598 23980
rect 185170 23968 185176 23980
rect 177592 23940 185176 23968
rect 177592 23928 177598 23940
rect 185170 23928 185176 23940
rect 185228 23928 185234 23980
rect 142482 23900 142488 23912
rect 140844 23872 142488 23900
rect 142482 23860 142488 23872
rect 142540 23860 142546 23912
rect 177718 23860 177724 23912
rect 177776 23900 177782 23912
rect 185262 23900 185268 23912
rect 177776 23872 185268 23900
rect 177776 23860 177782 23872
rect 185262 23860 185268 23872
rect 185320 23860 185326 23912
rect 134754 22976 134760 23028
rect 134812 23016 134818 23028
rect 140734 23016 140740 23028
rect 134812 22988 140740 23016
rect 134812 22976 134818 22988
rect 140734 22976 140740 22988
rect 140792 22976 140798 23028
rect 185262 22812 185268 22824
rect 181048 22784 185268 22812
rect 51218 22704 51224 22756
rect 51276 22744 51282 22756
rect 55910 22744 55916 22756
rect 51276 22716 55916 22744
rect 51276 22704 51282 22716
rect 55910 22704 55916 22716
rect 55968 22704 55974 22756
rect 100990 22744 100996 22756
rect 96868 22716 100996 22744
rect 50206 22636 50212 22688
rect 50264 22676 50270 22688
rect 50264 22648 56784 22676
rect 50264 22636 50270 22648
rect 56756 22608 56784 22648
rect 58210 22608 58216 22620
rect 56756 22580 58216 22608
rect 58210 22568 58216 22580
rect 58268 22568 58274 22620
rect 93998 22568 94004 22620
rect 94056 22608 94062 22620
rect 96868 22608 96896 22716
rect 100990 22704 100996 22716
rect 101048 22704 101054 22756
rect 134754 22704 134760 22756
rect 134812 22744 134818 22756
rect 139722 22744 139728 22756
rect 134812 22716 139728 22744
rect 134812 22704 134818 22716
rect 139722 22704 139728 22716
rect 139780 22704 139786 22756
rect 101082 22676 101088 22688
rect 94056 22580 96896 22608
rect 96960 22648 101088 22676
rect 94056 22568 94062 22580
rect 93906 22500 93912 22552
rect 93964 22540 93970 22552
rect 96960 22540 96988 22648
rect 101082 22636 101088 22648
rect 101140 22636 101146 22688
rect 134570 22636 134576 22688
rect 134628 22676 134634 22688
rect 134628 22648 140964 22676
rect 134628 22636 134634 22648
rect 100990 22608 100996 22620
rect 93964 22512 96988 22540
rect 97052 22580 100996 22608
rect 93964 22500 93970 22512
rect 90689 22407 90747 22413
rect 90689 22373 90701 22407
rect 90735 22404 90747 22407
rect 97052 22404 97080 22580
rect 100990 22568 100996 22580
rect 101048 22568 101054 22620
rect 134386 22568 134392 22620
rect 134444 22608 134450 22620
rect 134754 22608 134760 22620
rect 134444 22580 134760 22608
rect 134444 22568 134450 22580
rect 134754 22568 134760 22580
rect 134812 22568 134818 22620
rect 140936 22608 140964 22648
rect 142390 22608 142396 22620
rect 140936 22580 142396 22608
rect 142390 22568 142396 22580
rect 142448 22568 142454 22620
rect 177626 22568 177632 22620
rect 177684 22608 177690 22620
rect 181048 22608 181076 22784
rect 185262 22772 185268 22784
rect 185320 22772 185326 22824
rect 185170 22676 185176 22688
rect 177684 22580 181076 22608
rect 182336 22648 185176 22676
rect 177684 22568 177690 22580
rect 101082 22540 101088 22552
rect 90735 22376 97080 22404
rect 97144 22512 101088 22540
rect 90735 22373 90747 22376
rect 90689 22367 90747 22373
rect 96114 22296 96120 22348
rect 96172 22336 96178 22348
rect 97144 22336 97172 22512
rect 101082 22500 101088 22512
rect 101140 22500 101146 22552
rect 140734 22500 140740 22552
rect 140792 22540 140798 22552
rect 142482 22540 142488 22552
rect 140792 22512 142488 22540
rect 140792 22500 140798 22512
rect 142482 22500 142488 22512
rect 142540 22500 142546 22552
rect 177718 22500 177724 22552
rect 177776 22540 177782 22552
rect 182336 22540 182364 22648
rect 185170 22636 185176 22648
rect 185228 22636 185234 22688
rect 177776 22512 182364 22540
rect 177776 22500 177782 22512
rect 174406 22432 174412 22484
rect 174464 22472 174470 22484
rect 185170 22472 185176 22484
rect 174464 22444 185176 22472
rect 174464 22432 174470 22444
rect 185170 22432 185176 22444
rect 185228 22432 185234 22484
rect 96172 22308 97172 22336
rect 96172 22296 96178 22308
rect 55910 22160 55916 22212
rect 55968 22200 55974 22212
rect 58302 22200 58308 22212
rect 55968 22172 58308 22200
rect 55968 22160 55974 22172
rect 58302 22160 58308 22172
rect 58360 22160 58366 22212
rect 51218 21276 51224 21328
rect 51276 21316 51282 21328
rect 51276 21288 56784 21316
rect 51276 21276 51282 21288
rect 56756 21248 56784 21288
rect 58210 21248 58216 21260
rect 56756 21220 58216 21248
rect 58210 21208 58216 21220
rect 58268 21208 58274 21260
rect 93998 21208 94004 21260
rect 94056 21248 94062 21260
rect 101174 21248 101180 21260
rect 94056 21220 101180 21248
rect 94056 21208 94062 21220
rect 101174 21208 101180 21220
rect 101232 21208 101238 21260
rect 137974 21208 137980 21260
rect 138032 21248 138038 21260
rect 138158 21248 138164 21260
rect 138032 21220 138164 21248
rect 138032 21208 138038 21220
rect 138158 21208 138164 21220
rect 138216 21208 138222 21260
rect 139722 21208 139728 21260
rect 139780 21248 139786 21260
rect 143678 21248 143684 21260
rect 139780 21220 143684 21248
rect 139780 21208 139786 21220
rect 143678 21208 143684 21220
rect 143736 21208 143742 21260
rect 177718 21208 177724 21260
rect 177776 21248 177782 21260
rect 185262 21248 185268 21260
rect 177776 21220 185268 21248
rect 177776 21208 177782 21220
rect 185262 21208 185268 21220
rect 185320 21208 185326 21260
rect 93354 19780 93360 19832
rect 93412 19820 93418 19832
rect 101818 19820 101824 19832
rect 93412 19792 101824 19820
rect 93412 19780 93418 19792
rect 101818 19780 101824 19792
rect 101876 19780 101882 19832
rect 176154 19780 176160 19832
rect 176212 19820 176218 19832
rect 185262 19820 185268 19832
rect 176212 19792 185268 19820
rect 176212 19780 176218 19792
rect 185262 19780 185268 19792
rect 185320 19780 185326 19832
rect 94734 19712 94740 19764
rect 94792 19752 94798 19764
rect 101542 19752 101548 19764
rect 94792 19724 101548 19752
rect 94792 19712 94798 19724
rect 101542 19712 101548 19724
rect 101600 19712 101606 19764
rect 177810 19712 177816 19764
rect 177868 19752 177874 19764
rect 185170 19752 185176 19764
rect 177868 19724 185176 19752
rect 177868 19712 177874 19724
rect 185170 19712 185176 19724
rect 185228 19712 185234 19764
rect 18098 18420 18104 18472
rect 18156 18460 18162 18472
rect 68238 18460 68244 18472
rect 18156 18432 68244 18460
rect 18156 18420 18162 18432
rect 68238 18420 68244 18432
rect 68296 18420 68302 18472
rect 76061 18463 76119 18469
rect 76061 18429 76073 18463
rect 76107 18460 76119 18463
rect 80658 18460 80664 18472
rect 76107 18432 80664 18460
rect 76107 18429 76119 18432
rect 76061 18423 76119 18429
rect 80658 18420 80664 18432
rect 80716 18420 80722 18472
rect 106513 18463 106571 18469
rect 106513 18429 106525 18463
rect 106559 18460 106571 18463
rect 106694 18460 106700 18472
rect 106559 18432 106700 18460
rect 106559 18429 106571 18432
rect 106513 18423 106571 18429
rect 106694 18420 106700 18432
rect 106752 18460 106758 18472
rect 109733 18463 109791 18469
rect 109733 18460 109745 18463
rect 106752 18432 109745 18460
rect 106752 18420 106758 18432
rect 109733 18429 109745 18432
rect 109779 18429 109791 18463
rect 109733 18423 109791 18429
rect 112214 18420 112220 18472
rect 112272 18460 112278 18472
rect 152234 18460 152240 18472
rect 112272 18432 152240 18460
rect 112272 18420 112278 18432
rect 152234 18420 152240 18432
rect 152292 18420 152298 18472
rect 153430 18420 153436 18472
rect 153488 18460 153494 18472
rect 194922 18460 194928 18472
rect 153488 18432 194928 18460
rect 153488 18420 153494 18432
rect 194922 18420 194928 18432
rect 194980 18460 194986 18472
rect 212494 18460 212500 18472
rect 194980 18432 212500 18460
rect 194980 18420 194986 18432
rect 212494 18420 212500 18432
rect 212552 18420 212558 18472
rect 69894 18352 69900 18404
rect 69952 18392 69958 18404
rect 74773 18395 74831 18401
rect 74773 18392 74785 18395
rect 69952 18364 74785 18392
rect 69952 18352 69958 18364
rect 74773 18361 74785 18364
rect 74819 18361 74831 18395
rect 74773 18355 74831 18361
rect 138158 18352 138164 18404
rect 138216 18392 138222 18404
rect 145153 18395 145211 18401
rect 145153 18392 145165 18395
rect 138216 18364 145165 18392
rect 138216 18352 138222 18364
rect 145153 18361 145165 18364
rect 145199 18361 145211 18395
rect 145153 18355 145211 18361
rect 60786 18284 60792 18336
rect 60844 18324 60850 18336
rect 60844 18296 76196 18324
rect 60844 18284 60850 18296
rect 54806 18216 54812 18268
rect 54864 18256 54870 18268
rect 76061 18259 76119 18265
rect 76061 18256 76073 18259
rect 54864 18228 76073 18256
rect 54864 18216 54870 18228
rect 76061 18225 76073 18228
rect 76107 18225 76119 18259
rect 76168 18256 76196 18296
rect 76242 18284 76248 18336
rect 76300 18324 76306 18336
rect 78910 18324 78916 18336
rect 76300 18296 78916 18324
rect 76300 18284 76306 18296
rect 78910 18284 78916 18296
rect 78968 18284 78974 18336
rect 96761 18327 96819 18333
rect 96761 18293 96773 18327
rect 96807 18324 96819 18327
rect 106513 18327 106571 18333
rect 106513 18324 106525 18327
rect 96807 18296 106525 18324
rect 96807 18293 96819 18296
rect 96761 18287 96819 18293
rect 106513 18293 106525 18296
rect 106559 18293 106571 18327
rect 106513 18287 106571 18293
rect 165942 18284 165948 18336
rect 166000 18324 166006 18336
rect 166770 18324 166776 18336
rect 166000 18296 166776 18324
rect 166000 18284 166006 18296
rect 166770 18284 166776 18296
rect 166828 18284 166834 18336
rect 171370 18284 171376 18336
rect 171428 18324 171434 18336
rect 171922 18324 171928 18336
rect 171428 18296 171928 18324
rect 171428 18284 171434 18296
rect 171922 18284 171928 18296
rect 171980 18284 171986 18336
rect 79646 18256 79652 18268
rect 76168 18228 79652 18256
rect 76061 18219 76119 18225
rect 79646 18216 79652 18228
rect 79704 18216 79710 18268
rect 125741 18259 125799 18265
rect 125741 18225 125753 18259
rect 125787 18256 125799 18259
rect 128501 18259 128559 18265
rect 128501 18256 128513 18259
rect 125787 18228 128513 18256
rect 125787 18225 125799 18228
rect 125741 18219 125799 18225
rect 128501 18225 128513 18228
rect 128547 18225 128559 18259
rect 128501 18219 128559 18225
rect 128593 18259 128651 18265
rect 128593 18225 128605 18259
rect 128639 18256 128651 18259
rect 145153 18259 145211 18265
rect 128639 18228 129832 18256
rect 128639 18225 128651 18228
rect 128593 18219 128651 18225
rect 42846 18148 42852 18200
rect 42904 18188 42910 18200
rect 70630 18188 70636 18200
rect 42904 18160 70636 18188
rect 42904 18148 42910 18160
rect 70630 18148 70636 18160
rect 70688 18148 70694 18200
rect 109733 18191 109791 18197
rect 109733 18157 109745 18191
rect 109779 18188 109791 18191
rect 116173 18191 116231 18197
rect 116173 18188 116185 18191
rect 109779 18160 116185 18188
rect 109779 18157 109791 18160
rect 109733 18151 109791 18157
rect 116173 18157 116185 18160
rect 116219 18157 116231 18191
rect 129804 18188 129832 18228
rect 145153 18225 145165 18259
rect 145199 18256 145211 18259
rect 153430 18256 153436 18268
rect 145199 18228 153436 18256
rect 145199 18225 145211 18228
rect 145153 18219 145211 18225
rect 153430 18216 153436 18228
rect 153488 18216 153494 18268
rect 164286 18216 164292 18268
rect 164344 18256 164350 18268
rect 168518 18256 168524 18268
rect 164344 18228 168524 18256
rect 164344 18216 164350 18228
rect 168518 18216 168524 18228
rect 168576 18216 168582 18268
rect 138158 18188 138164 18200
rect 129804 18160 138164 18188
rect 116173 18151 116231 18157
rect 138158 18148 138164 18160
rect 138216 18148 138222 18200
rect 48826 18080 48832 18132
rect 48884 18120 48890 18132
rect 81670 18120 81676 18132
rect 48884 18092 81676 18120
rect 48884 18080 48890 18092
rect 81670 18080 81676 18092
rect 81728 18080 81734 18132
rect 87193 18123 87251 18129
rect 87193 18120 87205 18123
rect 85092 18092 87205 18120
rect 36774 18012 36780 18064
rect 36832 18052 36838 18064
rect 71366 18052 71372 18064
rect 36832 18024 71372 18052
rect 36832 18012 36838 18024
rect 71366 18012 71372 18024
rect 71424 18012 71430 18064
rect 74773 18055 74831 18061
rect 74773 18021 74785 18055
rect 74819 18052 74831 18055
rect 85092 18052 85120 18092
rect 87193 18089 87205 18092
rect 87239 18089 87251 18123
rect 87193 18083 87251 18089
rect 74819 18024 85120 18052
rect 116173 18055 116231 18061
rect 74819 18021 74831 18024
rect 74773 18015 74831 18021
rect 116173 18021 116185 18055
rect 116219 18052 116231 18055
rect 125741 18055 125799 18061
rect 125741 18052 125753 18055
rect 116219 18024 125753 18052
rect 116219 18021 116231 18024
rect 116173 18015 116231 18021
rect 125741 18021 125753 18024
rect 125787 18021 125799 18055
rect 125741 18015 125799 18021
rect 30794 17944 30800 17996
rect 30852 17984 30858 17996
rect 72378 17984 72384 17996
rect 30852 17956 72384 17984
rect 30852 17944 30858 17956
rect 72378 17944 72384 17956
rect 72436 17944 72442 17996
rect 87193 17987 87251 17993
rect 87193 17953 87205 17987
rect 87239 17984 87251 17987
rect 96761 17987 96819 17993
rect 96761 17984 96773 17987
rect 87239 17956 96773 17984
rect 87239 17953 87251 17956
rect 87193 17947 87251 17953
rect 96761 17953 96773 17956
rect 96807 17953 96819 17987
rect 96761 17947 96819 17953
rect 132822 17944 132828 17996
rect 132880 17984 132886 17996
rect 157570 17984 157576 17996
rect 132880 17956 157576 17984
rect 132880 17944 132886 17956
rect 157570 17944 157576 17956
rect 157628 17944 157634 17996
rect 167230 17944 167236 17996
rect 167288 17984 167294 17996
rect 167782 17984 167788 17996
rect 167288 17956 167788 17984
rect 167288 17944 167294 17956
rect 167782 17944 167788 17956
rect 167840 17944 167846 17996
rect 18834 17876 18840 17928
rect 18892 17916 18898 17928
rect 74770 17916 74776 17928
rect 18892 17888 74776 17916
rect 18892 17876 18898 17888
rect 74770 17876 74776 17888
rect 74828 17876 74834 17928
rect 138802 17876 138808 17928
rect 138860 17916 138866 17928
rect 156374 17916 156380 17928
rect 138860 17888 156380 17916
rect 138860 17876 138866 17888
rect 156374 17876 156380 17888
rect 156432 17876 156438 17928
rect 24814 17808 24820 17860
rect 24872 17848 24878 17860
rect 73390 17848 73396 17860
rect 24872 17820 73396 17848
rect 24872 17808 24878 17820
rect 73390 17808 73396 17820
rect 73448 17808 73454 17860
rect 126842 17808 126848 17860
rect 126900 17848 126906 17860
rect 158490 17848 158496 17860
rect 126900 17820 158496 17848
rect 126900 17808 126906 17820
rect 158490 17808 158496 17820
rect 158548 17808 158554 17860
rect 12854 17740 12860 17792
rect 12912 17780 12918 17792
rect 75506 17780 75512 17792
rect 12912 17752 75512 17780
rect 12912 17740 12918 17752
rect 75506 17740 75512 17752
rect 75564 17740 75570 17792
rect 86454 17740 86460 17792
rect 86512 17780 86518 17792
rect 96850 17780 96856 17792
rect 86512 17752 96856 17780
rect 86512 17740 86518 17752
rect 96850 17740 96856 17752
rect 96908 17740 96914 17792
rect 120862 17740 120868 17792
rect 120920 17780 120926 17792
rect 159502 17780 159508 17792
rect 120920 17752 159508 17780
rect 120920 17740 120926 17752
rect 159502 17740 159508 17752
rect 159560 17740 159566 17792
rect 77162 17536 77168 17588
rect 77220 17576 77226 17588
rect 78818 17576 78824 17588
rect 77220 17548 78824 17576
rect 77220 17536 77226 17548
rect 78818 17536 78824 17548
rect 78876 17536 78882 17588
rect 162906 17536 162912 17588
rect 162964 17576 162970 17588
rect 167138 17576 167144 17588
rect 162964 17548 167144 17576
rect 162964 17536 162970 17548
rect 167138 17536 167144 17548
rect 167196 17536 167202 17588
rect 169990 17536 169996 17588
rect 170048 17576 170054 17588
rect 170910 17576 170916 17588
rect 170048 17548 170916 17576
rect 170048 17536 170054 17548
rect 170910 17536 170916 17548
rect 170968 17536 170974 17588
rect 76150 17468 76156 17520
rect 76208 17508 76214 17520
rect 77530 17508 77536 17520
rect 76208 17480 77536 17508
rect 76208 17468 76214 17480
rect 77530 17468 77536 17480
rect 77588 17468 77594 17520
rect 162814 17400 162820 17452
rect 162872 17440 162878 17452
rect 164654 17440 164660 17452
rect 162872 17412 164660 17440
rect 162872 17400 162878 17412
rect 164654 17400 164660 17412
rect 164712 17400 164718 17452
rect 87558 17196 87564 17248
rect 87616 17236 87622 17248
rect 88938 17236 88944 17248
rect 87616 17208 88944 17236
rect 87616 17196 87622 17208
rect 88938 17196 88944 17208
rect 88996 17196 89002 17248
rect 84798 17128 84804 17180
rect 84856 17168 84862 17180
rect 87926 17168 87932 17180
rect 84856 17140 87932 17168
rect 84856 17128 84862 17140
rect 87926 17128 87932 17140
rect 87984 17128 87990 17180
rect 150854 17128 150860 17180
rect 150912 17168 150918 17180
rect 154350 17168 154356 17180
rect 150912 17140 154356 17168
rect 150912 17128 150918 17140
rect 154350 17128 154356 17140
rect 154408 17128 154414 17180
rect 67778 17060 67784 17112
rect 67836 17100 67842 17112
rect 117826 17100 117832 17112
rect 67836 17072 117832 17100
rect 67836 17060 67842 17072
rect 117826 17060 117832 17072
rect 117884 17060 117890 17112
rect 151866 17060 151872 17112
rect 151924 17100 151930 17112
rect 208906 17100 208912 17112
rect 151924 17072 208912 17100
rect 151924 17060 151930 17072
rect 208906 17060 208912 17072
rect 208964 17060 208970 17112
rect 167138 12776 167144 12828
rect 167196 12816 167202 12828
rect 174866 12816 174872 12828
rect 167196 12788 174872 12816
rect 167196 12776 167202 12788
rect 174866 12776 174872 12788
rect 174924 12776 174930 12828
rect 161802 12708 161808 12760
rect 161860 12748 161866 12760
rect 180846 12748 180852 12760
rect 161860 12720 180852 12748
rect 161860 12708 161866 12720
rect 180846 12708 180852 12720
rect 180904 12708 180910 12760
rect 171370 12640 171376 12692
rect 171428 12680 171434 12692
rect 192806 12680 192812 12692
rect 171428 12652 192812 12680
rect 171428 12640 171434 12652
rect 192806 12640 192812 12652
rect 192864 12640 192870 12692
rect 160330 12572 160336 12624
rect 160388 12612 160394 12624
rect 186826 12612 186832 12624
rect 160388 12584 186832 12612
rect 160388 12572 160394 12584
rect 186826 12572 186832 12584
rect 186884 12572 186890 12624
rect 85442 12504 85448 12556
rect 85500 12544 85506 12556
rect 85500 12516 94780 12544
rect 85500 12504 85506 12516
rect 88938 12368 88944 12420
rect 88996 12408 89002 12420
rect 90778 12408 90784 12420
rect 88996 12380 90784 12408
rect 88996 12368 89002 12380
rect 90778 12368 90784 12380
rect 90836 12368 90842 12420
rect 94752 12408 94780 12516
rect 169990 12504 169996 12556
rect 170048 12544 170054 12556
rect 198786 12544 198792 12556
rect 170048 12516 198792 12544
rect 170048 12504 170054 12516
rect 198786 12504 198792 12516
rect 198844 12504 198850 12556
rect 170082 12436 170088 12488
rect 170140 12476 170146 12488
rect 204858 12476 204864 12488
rect 170140 12448 204864 12476
rect 170140 12436 170146 12448
rect 204858 12436 204864 12448
rect 204916 12436 204922 12488
rect 102830 12408 102836 12420
rect 94752 12380 102836 12408
rect 102830 12368 102836 12380
rect 102888 12368 102894 12420
rect 168610 12368 168616 12420
rect 168668 12408 168674 12420
rect 210838 12408 210844 12420
rect 168668 12380 210844 12408
rect 168668 12368 168674 12380
rect 210838 12368 210844 12380
rect 210896 12368 210902 12420
rect 84338 12300 84344 12352
rect 84396 12340 84402 12352
rect 108810 12340 108816 12352
rect 84396 12312 108816 12340
rect 84396 12300 84402 12312
rect 108810 12300 108816 12312
rect 108868 12300 108874 12352
rect 167230 12300 167236 12352
rect 167288 12340 167294 12352
rect 216818 12340 216824 12352
rect 167288 12312 216824 12340
rect 167288 12300 167294 12312
rect 216818 12300 216824 12312
rect 216876 12300 216882 12352
rect 66858 12232 66864 12284
rect 66916 12272 66922 12284
rect 76242 12272 76248 12284
rect 66916 12244 76248 12272
rect 66916 12232 66922 12244
rect 76242 12232 76248 12244
rect 76300 12232 76306 12284
rect 83418 12232 83424 12284
rect 83476 12272 83482 12284
rect 114790 12272 114796 12284
rect 83476 12244 114796 12272
rect 83476 12232 83482 12244
rect 114790 12232 114796 12244
rect 114848 12232 114854 12284
rect 144782 12232 144788 12284
rect 144840 12272 144846 12284
rect 155362 12272 155368 12284
rect 144840 12244 155368 12272
rect 144840 12232 144846 12244
rect 155362 12232 155368 12244
rect 155420 12232 155426 12284
rect 156834 12232 156840 12284
rect 156892 12272 156898 12284
rect 165850 12272 165856 12284
rect 156892 12244 165856 12272
rect 156892 12232 156898 12244
rect 165850 12232 165856 12244
rect 165908 12232 165914 12284
rect 166126 12232 166132 12284
rect 166184 12272 166190 12284
rect 222798 12272 222804 12284
rect 166184 12244 222804 12272
rect 166184 12232 166190 12244
rect 222798 12232 222804 12244
rect 222856 12232 222862 12284
rect 72838 12096 72844 12148
rect 72896 12136 72902 12148
rect 76150 12136 76156 12148
rect 72896 12108 76156 12136
rect 72896 12096 72902 12108
rect 76150 12096 76156 12108
rect 76208 12096 76214 12148
<< via1 >>
rect 99616 244248 99668 244300
rect 99800 244248 99852 244300
rect 89864 241324 89916 241376
rect 171836 241324 171888 241376
rect 174044 241324 174096 241376
rect 207808 241324 207860 241376
rect 27856 241120 27908 241172
rect 29144 241120 29196 241172
rect 135864 240712 135916 240764
rect 136784 240712 136836 240764
rect 12768 236632 12820 236684
rect 30432 236632 30484 236684
rect 62540 236700 62592 236752
rect 107436 236632 107488 236684
rect 146536 236632 146588 236684
rect 23440 236564 23492 236616
rect 72844 236564 72896 236616
rect 121420 236564 121472 236616
rect 208912 236564 208964 236616
rect 218296 236564 218348 236616
rect 29144 235884 29196 235936
rect 82228 235884 82280 235936
rect 86184 235884 86236 235936
rect 99616 235884 99668 235936
rect 136784 235884 136836 235936
rect 169536 235884 169588 235936
rect 63828 235816 63880 235868
rect 166224 235816 166276 235868
rect 114428 235272 114480 235324
rect 159508 235272 159560 235324
rect 173492 235272 173544 235324
rect 174044 235272 174096 235324
rect 47544 235204 47596 235256
rect 65576 235204 65628 235256
rect 156840 235204 156892 235256
rect 215720 235204 215772 235256
rect 37424 235136 37476 235188
rect 75512 235136 75564 235188
rect 146536 235136 146588 235188
rect 216916 235136 216968 235188
rect 135404 233912 135456 233964
rect 142304 233912 142356 233964
rect 49936 233776 49988 233828
rect 58124 233776 58176 233828
rect 177172 233708 177224 233760
rect 185084 233708 185136 233760
rect 92716 233028 92768 233080
rect 100996 233028 101048 233080
rect 135404 232688 135456 232740
rect 142212 232688 142264 232740
rect 134300 232620 134352 232672
rect 142304 232620 142356 232672
rect 51224 232484 51276 232536
rect 58032 232484 58084 232536
rect 182324 232484 182376 232536
rect 185268 232484 185320 232536
rect 50580 232416 50632 232468
rect 58124 232416 58176 232468
rect 94004 232348 94056 232400
rect 100996 232416 101048 232468
rect 177724 232348 177776 232400
rect 185176 232416 185228 232468
rect 218296 232348 218348 232400
rect 222344 232348 222396 232400
rect 177724 231804 177776 231856
rect 182324 231804 182376 231856
rect 92716 231668 92768 231720
rect 100996 231668 101048 231720
rect 134852 231464 134904 231516
rect 139636 231464 139688 231516
rect 51224 231328 51276 231380
rect 56744 231328 56796 231380
rect 51132 231192 51184 231244
rect 51224 231056 51276 231108
rect 52696 231056 52748 231108
rect 95384 231124 95436 231176
rect 100996 231124 101048 231176
rect 135312 231056 135364 231108
rect 136876 231056 136928 231108
rect 178276 231056 178328 231108
rect 185268 231056 185320 231108
rect 94096 230988 94148 231040
rect 101088 230988 101140 231040
rect 135404 230988 135456 231040
rect 58216 230920 58268 230972
rect 92716 230852 92768 230904
rect 95384 230852 95436 230904
rect 177724 230920 177776 230972
rect 185176 230988 185228 231040
rect 143684 230852 143736 230904
rect 56744 230716 56796 230768
rect 58308 230716 58360 230768
rect 139636 230580 139688 230632
rect 142948 230580 143000 230632
rect 135312 229968 135364 230020
rect 139636 229968 139688 230020
rect 51224 229832 51276 229884
rect 56468 229832 56520 229884
rect 51132 229696 51184 229748
rect 56192 229696 56244 229748
rect 135404 229628 135456 229680
rect 52696 229560 52748 229612
rect 58216 229560 58268 229612
rect 92716 229560 92768 229612
rect 101088 229560 101140 229612
rect 143592 229560 143644 229612
rect 177632 229560 177684 229612
rect 185268 229560 185320 229612
rect 93176 229492 93228 229544
rect 100996 229492 101048 229544
rect 136876 229492 136928 229544
rect 143684 229492 143736 229544
rect 177816 229492 177868 229544
rect 185176 229492 185228 229544
rect 139636 229424 139688 229476
rect 143500 229424 143552 229476
rect 177724 229424 177776 229476
rect 185360 229424 185412 229476
rect 56192 229288 56244 229340
rect 58216 229288 58268 229340
rect 56468 229016 56520 229068
rect 58308 229016 58360 229068
rect 92716 228880 92768 228932
rect 100996 228880 101048 228932
rect 50764 228472 50816 228524
rect 55456 228472 55508 228524
rect 135404 228404 135456 228456
rect 51132 228336 51184 228388
rect 51224 228268 51276 228320
rect 52696 228268 52748 228320
rect 135312 228336 135364 228388
rect 135404 228268 135456 228320
rect 138164 228268 138216 228320
rect 58216 228200 58268 228252
rect 93176 228200 93228 228252
rect 101088 228200 101140 228252
rect 92716 228132 92768 228184
rect 100996 228132 101048 228184
rect 181128 228268 181180 228320
rect 185176 228268 185228 228320
rect 143684 228200 143736 228252
rect 177724 228200 177776 228252
rect 185636 228200 185688 228252
rect 143316 228132 143368 228184
rect 177632 228132 177684 228184
rect 185912 228132 185964 228184
rect 55456 227860 55508 227912
rect 58308 227860 58360 227912
rect 50948 227248 51000 227300
rect 56744 227248 56796 227300
rect 135404 226840 135456 226892
rect 52696 226772 52748 226824
rect 58216 226772 58268 226824
rect 93636 226772 93688 226824
rect 100996 226772 101048 226824
rect 182324 226840 182376 226892
rect 185268 226840 185320 226892
rect 143316 226772 143368 226824
rect 177632 226772 177684 226824
rect 185176 226772 185228 226824
rect 92716 226704 92768 226756
rect 101088 226704 101140 226756
rect 138164 226704 138216 226756
rect 143684 226704 143736 226756
rect 56744 226636 56796 226688
rect 58308 226636 58360 226688
rect 177724 226636 177776 226688
rect 181128 226636 181180 226688
rect 50488 225548 50540 225600
rect 58400 225548 58452 225600
rect 134576 225548 134628 225600
rect 143500 225548 143552 225600
rect 50764 225480 50816 225532
rect 58308 225480 58360 225532
rect 135220 225480 135272 225532
rect 143592 225480 143644 225532
rect 51316 225412 51368 225464
rect 58216 225412 58268 225464
rect 92808 225412 92860 225464
rect 101088 225412 101140 225464
rect 135496 225412 135548 225464
rect 143684 225412 143736 225464
rect 177632 225412 177684 225464
rect 185176 225412 185228 225464
rect 92900 225344 92952 225396
rect 100996 225344 101048 225396
rect 177816 225344 177868 225396
rect 185268 225344 185320 225396
rect 92716 225276 92768 225328
rect 101180 225276 101232 225328
rect 177724 225276 177776 225328
rect 182324 225276 182376 225328
rect 51040 224256 51092 224308
rect 52696 224256 52748 224308
rect 135220 224256 135272 224308
rect 136876 224256 136928 224308
rect 51132 224188 51184 224240
rect 51224 224120 51276 224172
rect 135312 224188 135364 224240
rect 135404 224120 135456 224172
rect 58216 224052 58268 224104
rect 93912 224052 93964 224104
rect 100996 224052 101048 224104
rect 58308 223984 58360 224036
rect 93728 223984 93780 224036
rect 101088 223984 101140 224036
rect 143684 224052 143736 224104
rect 177724 224052 177776 224104
rect 185360 224052 185412 224104
rect 143316 223984 143368 224036
rect 177356 223984 177408 224036
rect 185176 223984 185228 224036
rect 50948 223168 51000 223220
rect 56284 223168 56336 223220
rect 51224 223032 51276 223084
rect 52788 223032 52840 223084
rect 135312 223032 135364 223084
rect 137612 223032 137664 223084
rect 135404 222760 135456 222812
rect 52696 222692 52748 222744
rect 58216 222692 58268 222744
rect 92716 222692 92768 222744
rect 101456 222692 101508 222744
rect 143316 222692 143368 222744
rect 177632 222692 177684 222744
rect 185176 222692 185228 222744
rect 92992 222624 93044 222676
rect 101548 222624 101600 222676
rect 136876 222624 136928 222676
rect 143684 222624 143736 222676
rect 177724 222624 177776 222676
rect 185268 222624 185320 222676
rect 56284 222420 56336 222472
rect 58308 222420 58360 222472
rect 134852 222352 134904 222404
rect 139728 222352 139780 222404
rect 134484 221808 134536 221860
rect 139636 221808 139688 221860
rect 51224 221672 51276 221724
rect 56744 221672 56796 221724
rect 51132 221536 51184 221588
rect 55916 221536 55968 221588
rect 51224 221400 51276 221452
rect 52696 221400 52748 221452
rect 135312 221400 135364 221452
rect 136876 221400 136928 221452
rect 52788 221264 52840 221316
rect 58216 221264 58268 221316
rect 93176 221264 93228 221316
rect 101732 221264 101784 221316
rect 137612 221264 137664 221316
rect 143684 221264 143736 221316
rect 177632 221264 177684 221316
rect 185268 221264 185320 221316
rect 93728 221196 93780 221248
rect 101548 221196 101600 221248
rect 177816 221196 177868 221248
rect 185176 221196 185228 221248
rect 92716 221128 92768 221180
rect 101272 221128 101324 221180
rect 139728 221128 139780 221180
rect 143592 221128 143644 221180
rect 177724 221128 177776 221180
rect 185452 221128 185504 221180
rect 55916 220992 55968 221044
rect 58216 220992 58268 221044
rect 56744 220856 56796 220908
rect 58308 220856 58360 220908
rect 139636 220584 139688 220636
rect 143684 220584 143736 220636
rect 50948 220312 51000 220364
rect 56468 220312 56520 220364
rect 135312 220108 135364 220160
rect 138164 220108 138216 220160
rect 50212 219972 50264 220024
rect 52788 219972 52840 220024
rect 135404 219972 135456 220024
rect 52696 219904 52748 219956
rect 58216 219904 58268 219956
rect 92716 219904 92768 219956
rect 101824 219904 101876 219956
rect 143132 219904 143184 219956
rect 177632 219904 177684 219956
rect 185176 219904 185228 219956
rect 92808 219836 92860 219888
rect 101732 219836 101784 219888
rect 136876 219836 136928 219888
rect 143684 219836 143736 219888
rect 177724 219836 177776 219888
rect 185360 219836 185412 219888
rect 56468 219496 56520 219548
rect 58308 219496 58360 219548
rect 50212 218884 50264 218936
rect 53064 218884 53116 218936
rect 135036 218816 135088 218868
rect 137520 218816 137572 218868
rect 51224 218680 51276 218732
rect 52696 218680 52748 218732
rect 135404 218680 135456 218732
rect 50856 218612 50908 218664
rect 55456 218612 55508 218664
rect 135312 218612 135364 218664
rect 137980 218612 138032 218664
rect 52788 218544 52840 218596
rect 58216 218544 58268 218596
rect 92808 218544 92860 218596
rect 101916 218544 101968 218596
rect 185820 218612 185872 218664
rect 186004 218612 186056 218664
rect 143500 218544 143552 218596
rect 177724 218544 177776 218596
rect 185544 218544 185596 218596
rect 93728 218476 93780 218528
rect 101732 218476 101784 218528
rect 138164 218476 138216 218528
rect 143684 218476 143736 218528
rect 177632 218476 177684 218528
rect 185728 218476 185780 218528
rect 55456 218000 55508 218052
rect 58216 218000 58268 218052
rect 51224 217456 51276 217508
rect 52880 217456 52932 217508
rect 135404 217456 135456 217508
rect 137704 217456 137756 217508
rect 51224 217320 51276 217372
rect 52788 217320 52840 217372
rect 135404 217320 135456 217372
rect 137612 217320 137664 217372
rect 97960 217252 98012 217304
rect 101824 217252 101876 217304
rect 181036 217252 181088 217304
rect 185728 217252 185780 217304
rect 98052 217184 98104 217236
rect 101732 217184 101784 217236
rect 181220 217184 181272 217236
rect 185544 217184 185596 217236
rect 52696 217116 52748 217168
rect 58308 217116 58360 217168
rect 92716 217116 92768 217168
rect 101916 217116 101968 217168
rect 137520 217116 137572 217168
rect 143684 217116 143736 217168
rect 177724 217116 177776 217168
rect 185636 217116 185688 217168
rect 53064 217048 53116 217100
rect 58216 217048 58268 217100
rect 93912 217048 93964 217100
rect 102008 217048 102060 217100
rect 137980 217048 138032 217100
rect 143132 217048 143184 217100
rect 177632 217048 177684 217100
rect 185912 217048 185964 217100
rect 51132 215824 51184 215876
rect 56652 215824 56704 215876
rect 98144 215824 98196 215876
rect 101732 215824 101784 215876
rect 135404 215824 135456 215876
rect 52788 215756 52840 215808
rect 58308 215756 58360 215808
rect 93544 215756 93596 215808
rect 101824 215756 101876 215808
rect 181128 215824 181180 215876
rect 185728 215824 185780 215876
rect 143500 215756 143552 215808
rect 177632 215756 177684 215808
rect 185912 215756 185964 215808
rect 52880 215688 52932 215740
rect 58216 215688 58268 215740
rect 92716 215688 92768 215740
rect 97960 215688 98012 215740
rect 137704 215688 137756 215740
rect 143132 215688 143184 215740
rect 92808 215620 92860 215672
rect 98052 215620 98104 215672
rect 137612 215620 137664 215672
rect 142948 215620 143000 215672
rect 177724 215620 177776 215672
rect 181036 215620 181088 215672
rect 177724 215484 177776 215536
rect 181220 215484 181272 215536
rect 56652 215144 56704 215196
rect 58216 215144 58268 215196
rect 50396 214872 50448 214924
rect 52788 214872 52840 214924
rect 134852 214872 134904 214924
rect 137612 214872 137664 214924
rect 51132 214532 51184 214584
rect 52696 214532 52748 214584
rect 135312 214532 135364 214584
rect 136876 214532 136928 214584
rect 181220 214532 181272 214584
rect 185268 214532 185320 214584
rect 51224 214464 51276 214516
rect 58308 214464 58360 214516
rect 98052 214464 98104 214516
rect 101824 214464 101876 214516
rect 135404 214464 135456 214516
rect 143684 214464 143736 214516
rect 181036 214464 181088 214516
rect 185728 214464 185780 214516
rect 51316 214396 51368 214448
rect 58216 214396 58268 214448
rect 92716 214396 92768 214448
rect 100996 214396 101048 214448
rect 135496 214396 135548 214448
rect 142948 214396 143000 214448
rect 177632 214396 177684 214448
rect 185636 214396 185688 214448
rect 92808 214328 92860 214380
rect 98144 214328 98196 214380
rect 177724 214260 177776 214312
rect 181128 214260 181180 214312
rect 50212 213376 50264 213428
rect 52880 213376 52932 213428
rect 135404 213376 135456 213428
rect 137520 213376 137572 213428
rect 50948 213240 51000 213292
rect 52972 213240 53024 213292
rect 97960 213172 98012 213224
rect 101180 213172 101232 213224
rect 181956 213172 182008 213224
rect 185176 213172 185228 213224
rect 98144 213104 98196 213156
rect 101088 213104 101140 213156
rect 134668 213104 134720 213156
rect 136968 213104 137020 213156
rect 181864 213104 181916 213156
rect 185728 213104 185780 213156
rect 52696 213036 52748 213088
rect 58308 213036 58360 213088
rect 93636 213036 93688 213088
rect 100996 213036 101048 213088
rect 137612 213036 137664 213088
rect 143684 213036 143736 213088
rect 177724 213036 177776 213088
rect 181036 213036 181088 213088
rect 52788 212968 52840 213020
rect 58216 212968 58268 213020
rect 92716 212968 92768 213020
rect 98052 212968 98104 213020
rect 136876 212968 136928 213020
rect 143500 212968 143552 213020
rect 177724 212492 177776 212544
rect 181220 212492 181272 212544
rect 51224 212016 51276 212068
rect 52696 212016 52748 212068
rect 135404 212016 135456 212068
rect 137612 212016 137664 212068
rect 50764 211880 50816 211932
rect 56468 211880 56520 211932
rect 134852 211880 134904 211932
rect 139636 211880 139688 211932
rect 98052 211744 98104 211796
rect 101088 211744 101140 211796
rect 182140 211744 182192 211796
rect 185728 211744 185780 211796
rect 52972 211608 53024 211660
rect 58216 211608 58268 211660
rect 93544 211608 93596 211660
rect 100996 211676 101048 211728
rect 181680 211676 181732 211728
rect 185912 211676 185964 211728
rect 136968 211608 137020 211660
rect 143684 211608 143736 211660
rect 177724 211608 177776 211660
rect 181864 211608 181916 211660
rect 52880 211540 52932 211592
rect 58308 211540 58360 211592
rect 92808 211540 92860 211592
rect 98144 211540 98196 211592
rect 92716 211472 92768 211524
rect 97960 211472 98012 211524
rect 137520 211336 137572 211388
rect 143684 211336 143736 211388
rect 177724 211268 177776 211320
rect 181956 211268 182008 211320
rect 56468 211064 56520 211116
rect 58400 211064 58452 211116
rect 177724 210996 177776 211048
rect 182140 210996 182192 211048
rect 139636 210928 139688 210980
rect 143592 210928 143644 210980
rect 51132 210656 51184 210708
rect 56284 210656 56336 210708
rect 94096 210452 94148 210504
rect 101180 210452 101232 210504
rect 178276 210452 178328 210504
rect 185728 210452 185780 210504
rect 94004 210384 94056 210436
rect 101088 210384 101140 210436
rect 178092 210384 178144 210436
rect 185820 210384 185872 210436
rect 92624 210316 92676 210368
rect 100996 210316 101048 210368
rect 135404 210316 135456 210368
rect 52696 210248 52748 210300
rect 58216 210248 58268 210300
rect 92716 210248 92768 210300
rect 98052 210248 98104 210300
rect 176804 210316 176856 210368
rect 186004 210316 186056 210368
rect 143684 210248 143736 210300
rect 137612 210180 137664 210232
rect 142948 210180 143000 210232
rect 177724 210044 177776 210096
rect 181680 210044 181732 210096
rect 56284 209908 56336 209960
rect 58308 209908 58360 209960
rect 91244 209024 91296 209076
rect 101088 209024 101140 209076
rect 175424 209024 175476 209076
rect 185728 209024 185780 209076
rect 83056 208956 83108 209008
rect 84252 208956 84304 209008
rect 90600 208956 90652 209008
rect 100996 208956 101048 209008
rect 174780 208956 174832 209008
rect 185820 208956 185872 209008
rect 51224 207664 51276 207716
rect 56100 207664 56152 207716
rect 135404 207596 135456 207648
rect 140280 207596 140332 207648
rect 50580 207460 50632 207512
rect 61252 207460 61304 207512
rect 87564 207460 87616 207512
rect 101640 207460 101692 207512
rect 134760 207460 134812 207512
rect 145340 207460 145392 207512
rect 171192 207460 171244 207512
rect 185912 207460 185964 207512
rect 174044 207392 174096 207444
rect 187936 207392 187988 207444
rect 172572 206916 172624 206968
rect 177540 206916 177592 206968
rect 148744 206780 148796 206832
rect 149388 206780 149440 206832
rect 90416 206508 90468 206560
rect 91152 206508 91204 206560
rect 63276 206236 63328 206288
rect 65116 206236 65168 206288
rect 64748 206168 64800 206220
rect 65208 206168 65260 206220
rect 66128 206168 66180 206220
rect 66588 206168 66640 206220
rect 72108 206168 72160 206220
rect 72660 206168 72712 206220
rect 73396 206168 73448 206220
rect 74040 206168 74092 206220
rect 74776 206168 74828 206220
rect 75512 206168 75564 206220
rect 76156 206168 76208 206220
rect 76892 206168 76944 206220
rect 77536 206168 77588 206220
rect 78364 206168 78416 206220
rect 85724 206168 85776 206220
rect 100996 206168 101048 206220
rect 147272 206168 147324 206220
rect 149296 206168 149348 206220
rect 150124 206168 150176 206220
rect 150768 206168 150820 206220
rect 152976 206168 153028 206220
rect 153528 206168 153580 206220
rect 156196 206168 156248 206220
rect 156656 206168 156708 206220
rect 157576 206168 157628 206220
rect 158036 206168 158088 206220
rect 158956 206168 159008 206220
rect 159508 206168 159560 206220
rect 160336 206168 160388 206220
rect 160888 206168 160940 206220
rect 169904 206168 169956 206220
rect 185176 206168 185228 206220
rect 205416 204672 205468 204724
rect 208360 204672 208412 204724
rect 22796 204604 22848 204656
rect 26844 204604 26896 204656
rect 121420 204604 121472 204656
rect 124272 204604 124324 204656
rect 23440 204536 23492 204588
rect 26752 204536 26804 204588
rect 208360 204536 208412 204588
rect 211120 204536 211172 204588
rect 26660 204468 26712 204520
rect 27764 204468 27816 204520
rect 208544 204468 208596 204520
rect 212224 204468 212276 204520
rect 24084 204400 24136 204452
rect 28040 204400 28092 204452
rect 98972 204400 99024 204452
rect 104768 204400 104820 204452
rect 120224 204400 120276 204452
rect 121512 204400 121564 204452
rect 208268 204400 208320 204452
rect 210568 204400 210620 204452
rect 22152 204332 22204 204384
rect 26660 204332 26712 204384
rect 24728 204264 24780 204316
rect 28132 204264 28184 204316
rect 99432 204264 99484 204316
rect 107528 204264 107580 204316
rect 121512 204264 121564 204316
rect 123168 204264 123220 204316
rect 121604 204196 121656 204248
rect 123720 204196 123772 204248
rect 208452 204196 208504 204248
rect 211672 204196 211724 204248
rect 99248 204128 99300 204180
rect 106976 204128 107028 204180
rect 183612 204128 183664 204180
rect 191340 204128 191392 204180
rect 20220 204060 20272 204112
rect 41748 204060 41800 204112
rect 99524 204060 99576 204112
rect 108080 204060 108132 204112
rect 183428 204060 183480 204112
rect 190788 204060 190840 204112
rect 191984 204060 192036 204112
rect 214432 204060 214484 204112
rect 99156 203788 99208 203840
rect 106424 203788 106476 203840
rect 124272 203788 124324 203840
rect 128228 203788 128280 203840
rect 123720 203720 123772 203772
rect 125468 203720 125520 203772
rect 187200 203720 187252 203772
rect 191892 203720 191944 203772
rect 21508 203652 21560 203704
rect 26936 203652 26988 203704
rect 36044 203652 36096 203704
rect 37056 203652 37108 203704
rect 124180 203652 124232 203704
rect 127124 203652 127176 203704
rect 183336 203652 183388 203704
rect 190236 203652 190288 203704
rect 40920 203584 40972 203636
rect 43588 203584 43640 203636
rect 45060 203584 45112 203636
rect 46164 203584 46216 203636
rect 99340 203584 99392 203636
rect 105872 203584 105924 203636
rect 120132 203584 120184 203636
rect 122616 203584 122668 203636
rect 123996 203584 124048 203636
rect 126572 203584 126624 203636
rect 127860 203584 127912 203636
rect 129884 203584 129936 203636
rect 183244 203584 183296 203636
rect 189132 203584 189184 203636
rect 201552 203584 201604 203636
rect 202840 203584 202892 203636
rect 204312 203584 204364 203636
rect 206152 203584 206204 203636
rect 39540 203516 39592 203568
rect 41012 203516 41064 203568
rect 41196 203516 41248 203568
rect 42944 203516 42996 203568
rect 99064 203516 99116 203568
rect 105320 203516 105372 203568
rect 118568 203516 118620 203568
rect 119856 203516 119908 203568
rect 120040 203516 120092 203568
rect 122064 203516 122116 203568
rect 123904 203516 123956 203568
rect 126020 203516 126072 203568
rect 128044 203516 128096 203568
rect 130436 203516 130488 203568
rect 183152 203516 183204 203568
rect 188580 203516 188632 203568
rect 37332 203448 37384 203500
rect 39080 203448 39132 203500
rect 41104 203448 41156 203500
rect 42300 203448 42352 203500
rect 20864 203380 20916 203432
rect 24360 203380 24412 203432
rect 25372 203380 25424 203432
rect 26292 203380 26344 203432
rect 27948 203380 28000 203432
rect 29144 203380 29196 203432
rect 29236 203380 29288 203432
rect 30248 203380 30300 203432
rect 31260 203380 31312 203432
rect 31812 203380 31864 203432
rect 37240 203380 37292 203432
rect 38344 203380 38396 203432
rect 39632 203380 39684 203432
rect 40368 203380 40420 203432
rect 41012 203380 41064 203432
rect 41656 203380 41708 203432
rect 33376 203040 33428 203092
rect 34204 203040 34256 203092
rect 34756 203040 34808 203092
rect 35492 203040 35544 203092
rect 45520 203448 45572 203500
rect 98880 203448 98932 203500
rect 104216 203448 104268 203500
rect 110288 203448 110340 203500
rect 111024 203448 111076 203500
rect 116084 203448 116136 203500
rect 117004 203448 117056 203500
rect 117648 203448 117700 203500
rect 118752 203448 118804 203500
rect 118844 203448 118896 203500
rect 120960 203448 121012 203500
rect 123812 203448 123864 203500
rect 124824 203448 124876 203500
rect 127952 203448 128004 203500
rect 129332 203448 129384 203500
rect 183060 203448 183112 203500
rect 188120 203448 188172 203500
rect 204496 203516 204548 203568
rect 205508 203516 205560 203568
rect 207808 203516 207860 203568
rect 207900 203516 207952 203568
rect 209464 203516 209516 203568
rect 204404 203448 204456 203500
rect 205600 203448 205652 203500
rect 205692 203448 205744 203500
rect 207256 203448 207308 203500
rect 208084 203448 208136 203500
rect 210016 203448 210068 203500
rect 43772 203380 43824 203432
rect 44876 203380 44928 203432
rect 108632 203380 108684 203432
rect 109276 203380 109328 203432
rect 109736 203380 109788 203432
rect 110932 203380 110984 203432
rect 111484 203380 111536 203432
rect 112312 203380 112364 203432
rect 115992 203380 116044 203432
rect 116452 203380 116504 203432
rect 117280 203380 117332 203432
rect 118200 203380 118252 203432
rect 118660 203380 118712 203432
rect 119304 203380 119356 203432
rect 118752 203312 118804 203364
rect 120408 203380 120460 203432
rect 124364 203380 124416 203432
rect 127676 203380 127728 203432
rect 128136 203380 128188 203432
rect 128780 203380 128832 203432
rect 183520 203380 183572 203432
rect 189684 203380 189736 203432
rect 192444 203380 192496 203432
rect 193364 203380 193416 203432
rect 193548 203380 193600 203432
rect 194652 203380 194704 203432
rect 201460 203380 201512 203432
rect 202288 203380 202340 203432
rect 202932 203380 202984 203432
rect 203024 203380 203076 203432
rect 203944 203380 203996 203432
rect 204220 203380 204272 203432
rect 205048 203380 205100 203432
rect 205416 203380 205468 203432
rect 205784 203380 205836 203432
rect 206704 203380 206756 203432
rect 207992 203380 208044 203432
rect 208912 203380 208964 203432
rect 205600 203312 205652 203364
rect 199160 203040 199212 203092
rect 199804 203040 199856 203092
rect 212868 203040 212920 203092
rect 213604 203040 213656 203092
rect 43680 202972 43732 203024
rect 30984 202836 31036 202888
rect 31904 202836 31956 202888
rect 197596 199504 197648 199556
rect 198148 199504 198200 199556
rect 122892 196444 122944 196496
rect 123996 196444 124048 196496
rect 194836 196444 194888 196496
rect 196032 196444 196084 196496
rect 26752 196376 26804 196428
rect 27396 196376 27448 196428
rect 30432 196376 30484 196428
rect 31260 196376 31312 196428
rect 31720 196376 31772 196428
rect 32824 196376 32876 196428
rect 39264 196376 39316 196428
rect 41104 196376 41156 196428
rect 115256 196376 115308 196428
rect 115900 196376 115952 196428
rect 119672 196376 119724 196428
rect 120040 196376 120092 196428
rect 123628 196376 123680 196428
rect 124364 196376 124416 196428
rect 125652 196376 125704 196428
rect 128044 196376 128096 196428
rect 194744 196376 194796 196428
rect 195664 196376 195716 196428
rect 203668 196376 203720 196428
rect 204404 196376 204456 196428
rect 24360 196308 24412 196360
rect 26108 196308 26160 196360
rect 26568 196308 26620 196360
rect 26936 196308 26988 196360
rect 27764 196308 27816 196360
rect 29696 196308 29748 196360
rect 30524 196308 30576 196360
rect 31628 196308 31680 196360
rect 31996 196308 32048 196360
rect 32916 196308 32968 196360
rect 33376 196308 33428 196360
rect 34480 196308 34532 196360
rect 34756 196308 34808 196360
rect 35308 196308 35360 196360
rect 36872 196308 36924 196360
rect 37240 196308 37292 196360
rect 37700 196308 37752 196360
rect 39356 196308 39408 196360
rect 40092 196308 40144 196360
rect 40920 196308 40972 196360
rect 41656 196308 41708 196360
rect 45060 196308 45112 196360
rect 56100 196308 56152 196360
rect 57572 196308 57624 196360
rect 67784 196308 67836 196360
rect 68612 196308 68664 196360
rect 80848 196308 80900 196360
rect 81676 196308 81728 196360
rect 81952 196308 82004 196360
rect 83056 196308 83108 196360
rect 89772 196308 89824 196360
rect 90600 196308 90652 196360
rect 93084 196308 93136 196360
rect 94004 196308 94056 196360
rect 109368 196308 109420 196360
rect 110288 196308 110340 196360
rect 114888 196308 114940 196360
rect 115348 196308 115400 196360
rect 116820 196308 116872 196360
rect 117280 196308 117332 196360
rect 119304 196308 119356 196360
rect 120224 196308 120276 196360
rect 120868 196308 120920 196360
rect 121604 196308 121656 196360
rect 123260 196308 123312 196360
rect 124180 196308 124232 196360
rect 125284 196308 125336 196360
rect 127860 196308 127912 196360
rect 140280 196308 140332 196360
rect 141568 196308 141620 196360
rect 163740 196308 163792 196360
rect 164476 196308 164528 196360
rect 164844 196308 164896 196360
rect 165856 196308 165908 196360
rect 173768 196308 173820 196360
rect 174780 196308 174832 196360
rect 175976 196308 176028 196360
rect 176804 196308 176856 196360
rect 177080 196308 177132 196360
rect 178184 196308 178236 196360
rect 194560 196308 194612 196360
rect 195296 196308 195348 196360
rect 196400 196308 196452 196360
rect 197228 196308 197280 196360
rect 197596 196308 197648 196360
rect 198424 196308 198476 196360
rect 199160 196308 199212 196360
rect 199620 196308 199672 196360
rect 202472 196308 202524 196360
rect 203024 196308 203076 196360
rect 203300 196308 203352 196360
rect 204220 196308 204272 196360
rect 204864 196308 204916 196360
rect 205692 196308 205744 196360
rect 206888 196308 206940 196360
rect 208084 196308 208136 196360
rect 27672 196240 27724 196292
rect 30064 196240 30116 196292
rect 165948 196240 166000 196292
rect 167236 196240 167288 196292
rect 122432 196172 122484 196224
rect 123904 196172 123956 196224
rect 29052 196104 29104 196156
rect 30892 196104 30944 196156
rect 51224 196104 51276 196156
rect 59780 196104 59832 196156
rect 202104 196104 202156 196156
rect 202840 196104 202892 196156
rect 207256 196104 207308 196156
rect 208268 196104 208320 196156
rect 38068 196036 38120 196088
rect 39632 196036 39684 196088
rect 51040 196036 51092 196088
rect 58676 196036 58728 196088
rect 122064 196036 122116 196088
rect 123720 196036 123772 196088
rect 135220 196036 135272 196088
rect 142672 196036 142724 196088
rect 38896 195968 38948 196020
rect 41012 195968 41064 196020
rect 50948 195968 51000 196020
rect 60884 195968 60936 196020
rect 117648 195968 117700 196020
rect 118660 195968 118712 196020
rect 121696 195968 121748 196020
rect 123812 195968 123864 196020
rect 134944 195968 134996 196020
rect 144880 195968 144932 196020
rect 193272 195968 193324 196020
rect 194468 195968 194520 196020
rect 200816 195968 200868 196020
rect 201644 195968 201696 196020
rect 39632 195900 39684 195952
rect 41196 195900 41248 195952
rect 50764 195900 50816 195952
rect 61988 195900 62040 195952
rect 88668 195900 88720 195952
rect 102100 195900 102152 195952
rect 135128 195900 135180 195952
rect 145984 195900 146036 195952
rect 172664 195900 172716 195952
rect 186096 195900 186148 195952
rect 204496 195900 204548 195952
rect 205784 195900 205836 195952
rect 206060 195900 206112 195952
rect 207992 195900 208044 195952
rect 209280 195900 209332 195952
rect 213052 195900 213104 195952
rect 50856 195832 50908 195884
rect 63092 195832 63144 195884
rect 91152 195832 91204 195884
rect 94188 195832 94240 195884
rect 134852 195832 134904 195884
rect 147088 195832 147140 195884
rect 171560 195832 171612 195884
rect 186280 195832 186332 195884
rect 208820 195832 208872 195884
rect 212960 195832 213012 195884
rect 26384 195764 26436 195816
rect 29236 195764 29288 195816
rect 50672 195764 50724 195816
rect 64196 195764 64248 195816
rect 86460 195764 86512 195816
rect 101732 195764 101784 195816
rect 124456 195764 124508 195816
rect 128136 195764 128188 195816
rect 135036 195764 135088 195816
rect 148192 195764 148244 195816
rect 170456 195764 170508 195816
rect 185912 195764 185964 195816
rect 209648 195764 209700 195816
rect 212868 195764 212920 195816
rect 38436 195696 38488 195748
rect 39540 195696 39592 195748
rect 41288 195696 41340 195748
rect 43680 195696 43732 195748
rect 87564 195696 87616 195748
rect 101916 195696 101968 195748
rect 110656 195696 110708 195748
rect 111668 195696 111720 195748
rect 118108 195696 118160 195748
rect 118568 195696 118620 195748
rect 135404 195696 135456 195748
rect 143776 195696 143828 195748
rect 26292 195628 26344 195680
rect 28868 195628 28920 195680
rect 40460 195628 40512 195680
rect 43128 195628 43180 195680
rect 33468 195560 33520 195612
rect 34112 195560 34164 195612
rect 36504 195560 36556 195612
rect 37424 195560 37476 195612
rect 40828 195560 40880 195612
rect 43772 195560 43824 195612
rect 116452 195560 116504 195612
rect 117372 195560 117424 195612
rect 124824 195560 124876 195612
rect 127952 195560 128004 195612
rect 135312 195560 135364 195612
rect 140464 195560 140516 195612
rect 120500 195492 120552 195544
rect 121512 195492 121564 195544
rect 51132 195424 51184 195476
rect 56468 195424 56520 195476
rect 112036 195424 112088 195476
rect 112496 195424 112548 195476
rect 29144 195288 29196 195340
rect 30432 195288 30484 195340
rect 31812 195288 31864 195340
rect 32456 195288 32508 195340
rect 177540 195288 177592 195340
rect 179288 195288 179340 195340
rect 206428 195288 206480 195340
rect 207900 195288 207952 195340
rect 182876 193180 182928 193232
rect 187200 193180 187252 193232
rect 18104 190936 18156 190988
rect 22336 190936 22388 190988
rect 187936 188216 187988 188268
rect 191984 188216 192036 188268
rect 99432 186856 99484 186908
rect 106792 186856 106844 186908
rect 13412 185496 13464 185548
rect 16080 185496 16132 185548
rect 104400 184068 104452 184120
rect 106792 184068 106844 184120
rect 13320 184000 13372 184052
rect 22336 184000 22388 184052
rect 99524 184000 99576 184052
rect 105780 184000 105832 184052
rect 182876 184000 182928 184052
rect 187936 184000 187988 184052
rect 104492 182708 104544 182760
rect 107160 182708 107212 182760
rect 128504 182708 128556 182760
rect 137520 182708 137572 182760
rect 98604 182640 98656 182692
rect 106976 182640 107028 182692
rect 183152 182640 183204 182692
rect 191156 182640 191208 182692
rect 183704 181280 183756 181332
rect 191984 181280 192036 181332
rect 105136 180328 105188 180380
rect 106976 180328 107028 180380
rect 98420 179852 98472 179904
rect 104492 179852 104544 179904
rect 182508 179852 182560 179904
rect 190696 179852 190748 179904
rect 212132 179852 212184 179904
rect 222344 179852 222396 179904
rect 183704 179784 183756 179836
rect 190604 179784 190656 179836
rect 99524 179512 99576 179564
rect 104400 179512 104452 179564
rect 44416 178560 44468 178612
rect 49292 178560 49344 178612
rect 182508 178492 182560 178544
rect 191984 178492 192036 178544
rect 99524 177336 99576 177388
rect 105136 177336 105188 177388
rect 16080 177132 16132 177184
rect 22336 177132 22388 177184
rect 98604 177132 98656 177184
rect 106792 177132 106844 177184
rect 183244 176452 183296 176504
rect 191984 176452 192036 176504
rect 211580 175840 211632 175892
rect 216180 175840 216232 175892
rect 98236 175772 98288 175824
rect 106608 175772 106660 175824
rect 183704 175092 183756 175144
rect 191524 175092 191576 175144
rect 49292 174344 49344 174396
rect 52696 174344 52748 174396
rect 99524 173664 99576 173716
rect 106792 173664 106844 173716
rect 183336 173052 183388 173104
rect 191984 173052 192036 173104
rect 99524 171692 99576 171744
rect 106792 171692 106844 171744
rect 183520 171692 183572 171744
rect 191156 171692 191208 171744
rect 182692 171216 182744 171268
rect 185084 171216 185136 171268
rect 99248 170264 99300 170316
rect 106792 170196 106844 170248
rect 99524 168904 99576 168956
rect 106700 168904 106752 168956
rect 182508 168904 182560 168956
rect 191892 168904 191944 168956
rect 185084 168836 185136 168888
rect 191984 168836 192036 168888
rect 99524 167612 99576 167664
rect 106884 167612 106936 167664
rect 44416 167544 44468 167596
rect 53340 167544 53392 167596
rect 99432 167544 99484 167596
rect 106792 167544 106844 167596
rect 183704 167544 183756 167596
rect 191340 167544 191392 167596
rect 182876 166456 182928 166508
rect 187936 166456 187988 166508
rect 99524 166184 99576 166236
rect 107252 166184 107304 166236
rect 183704 164960 183756 165012
rect 190052 164960 190104 165012
rect 99524 164756 99576 164808
rect 107160 164756 107212 164808
rect 211764 163600 211816 163652
rect 217008 163600 217060 163652
rect 99524 163396 99576 163448
rect 104400 163396 104452 163448
rect 128504 163396 128556 163448
rect 137520 163396 137572 163448
rect 183060 163396 183112 163448
rect 189960 163396 190012 163448
rect 13136 163328 13188 163380
rect 22980 163328 23032 163380
rect 183796 162988 183848 163040
rect 191524 162988 191576 163040
rect 187936 161968 187988 162020
rect 191984 161968 192036 162020
rect 212684 157072 212736 157124
rect 216916 157072 216968 157124
rect 216916 156460 216968 156512
rect 218296 156460 218348 156512
rect 182784 155440 182836 155492
rect 188028 155440 188080 155492
rect 104400 155032 104452 155084
rect 106516 155032 106568 155084
rect 212040 153672 212092 153724
rect 222252 153672 222304 153724
rect 32088 152312 32140 152364
rect 32824 152312 32876 152364
rect 33376 152312 33428 152364
rect 34112 152312 34164 152364
rect 36872 152312 36924 152364
rect 37424 152312 37476 152364
rect 37700 152312 37752 152364
rect 38804 152312 38856 152364
rect 41656 152312 41708 152364
rect 43680 152312 43732 152364
rect 110932 152312 110984 152364
rect 111668 152312 111720 152364
rect 113600 152312 113652 152364
rect 114060 152312 114112 152364
rect 117648 152312 117700 152364
rect 118844 152312 118896 152364
rect 119672 152312 119724 152364
rect 121972 152312 122024 152364
rect 124088 152312 124140 152364
rect 127860 152312 127912 152364
rect 197596 152312 197648 152364
rect 198056 152312 198108 152364
rect 200448 152312 200500 152364
rect 201184 152312 201236 152364
rect 201368 152312 201420 152364
rect 201644 152312 201696 152364
rect 203668 152312 203720 152364
rect 205968 152312 206020 152364
rect 35308 152244 35360 152296
rect 35952 152244 36004 152296
rect 36504 152244 36556 152296
rect 37332 152244 37384 152296
rect 38068 152244 38120 152296
rect 38620 152244 38672 152296
rect 118476 152244 118528 152296
rect 120592 152244 120644 152296
rect 124824 152244 124876 152296
rect 129332 152244 129384 152296
rect 203300 152244 203352 152296
rect 205876 152244 205928 152296
rect 207256 152244 207308 152296
rect 210752 152244 210804 152296
rect 39632 152176 39684 152228
rect 43128 152176 43180 152228
rect 118752 152176 118804 152228
rect 120960 152176 121012 152228
rect 196216 152176 196268 152228
rect 197228 152176 197280 152228
rect 204864 152176 204916 152228
rect 207348 152176 207400 152228
rect 39264 152108 39316 152160
rect 43036 152108 43088 152160
rect 120040 152108 120092 152160
rect 123168 152108 123220 152160
rect 204496 152108 204548 152160
rect 207256 152108 207308 152160
rect 41288 152040 41340 152092
rect 45152 152040 45204 152092
rect 109184 152040 109236 152092
rect 110104 152040 110156 152092
rect 119304 152040 119356 152092
rect 121788 152040 121840 152092
rect 124456 152040 124508 152092
rect 128780 152040 128832 152092
rect 205692 152040 205744 152092
rect 207992 152040 208044 152092
rect 40828 151972 40880 152024
rect 45060 151972 45112 152024
rect 122892 151904 122944 151956
rect 123260 151904 123312 151956
rect 127216 151904 127268 151956
rect 205232 151904 205284 151956
rect 207900 151904 207952 151956
rect 31812 151836 31864 151888
rect 32456 151836 32508 151888
rect 112128 151836 112180 151888
rect 112864 151836 112916 151888
rect 31996 151768 32048 151820
rect 33284 151768 33336 151820
rect 40460 151768 40512 151820
rect 44784 151768 44836 151820
rect 79192 151768 79244 151820
rect 96120 151768 96172 151820
rect 120868 151768 120920 151820
rect 123720 151768 123772 151820
rect 72568 151700 72620 151752
rect 98880 151700 98932 151752
rect 156564 151700 156616 151752
rect 69164 151632 69216 151684
rect 92532 151632 92584 151684
rect 96120 151632 96172 151684
rect 163188 151632 163240 151684
rect 40092 151564 40144 151616
rect 43772 151564 43824 151616
rect 123628 151564 123680 151616
rect 127952 151564 128004 151616
rect 127308 151496 127360 151548
rect 25004 151428 25056 151480
rect 28500 151428 28552 151480
rect 204036 151428 204088 151480
rect 206060 151428 206112 151480
rect 206428 151428 206480 151480
rect 210016 151428 210068 151480
rect 24912 151360 24964 151412
rect 28040 151360 28092 151412
rect 121696 151360 121748 151412
rect 124640 151360 124692 151412
rect 202472 151360 202524 151412
rect 203024 151360 203076 151412
rect 206888 151360 206940 151412
rect 210108 151360 210160 151412
rect 26384 151292 26436 151344
rect 29236 151292 29288 151344
rect 122432 151292 122484 151344
rect 125192 151292 125244 151344
rect 125652 151292 125704 151344
rect 131356 151292 131408 151344
rect 207624 151292 207676 151344
rect 210660 151292 210712 151344
rect 25740 151224 25792 151276
rect 27672 151224 27724 151276
rect 116452 151224 116504 151276
rect 117188 151224 117240 151276
rect 118108 151224 118160 151276
rect 120316 151224 120368 151276
rect 120500 151224 120552 151276
rect 123076 151224 123128 151276
rect 200816 151224 200868 151276
rect 201552 151224 201604 151276
rect 208820 151224 208872 151276
rect 212868 151224 212920 151276
rect 26292 151156 26344 151208
rect 28868 151156 28920 151208
rect 29144 151156 29196 151208
rect 30432 151156 30484 151208
rect 208084 151156 208136 151208
rect 210844 151156 210896 151208
rect 25924 151088 25976 151140
rect 27304 151088 27356 151140
rect 29052 151088 29104 151140
rect 30892 151088 30944 151140
rect 208452 151088 208504 151140
rect 210936 151088 210988 151140
rect 25832 151020 25884 151072
rect 26844 151020 26896 151072
rect 27672 151020 27724 151072
rect 30064 151020 30116 151072
rect 30432 151020 30484 151072
rect 31628 151020 31680 151072
rect 109368 151020 109420 151072
rect 110196 151020 110248 151072
rect 121236 151020 121288 151072
rect 123812 151020 123864 151072
rect 125284 151020 125336 151072
rect 129240 151020 129292 151072
rect 193364 151020 193416 151072
rect 194468 151020 194520 151072
rect 209280 151020 209332 151072
rect 214156 151020 214208 151072
rect 26016 150952 26068 151004
rect 26476 150952 26528 151004
rect 27764 150952 27816 151004
rect 29696 150952 29748 151004
rect 30524 150952 30576 151004
rect 31260 150952 31312 151004
rect 38896 150952 38948 151004
rect 41840 150952 41892 151004
rect 111300 150952 111352 151004
rect 115256 150952 115308 151004
rect 115808 150952 115860 151004
rect 122064 150952 122116 151004
rect 125100 150952 125152 151004
rect 193272 150952 193324 151004
rect 194100 150952 194152 151004
rect 195480 150952 195532 151004
rect 196032 150952 196084 151004
rect 196308 150952 196360 151004
rect 196860 150952 196912 151004
rect 202104 150952 202156 151004
rect 202748 150952 202800 151004
rect 206336 150952 206388 151004
rect 208820 150952 208872 151004
rect 209648 150952 209700 151004
rect 214248 150952 214300 151004
rect 110564 150884 110616 150936
rect 196216 148300 196268 148352
rect 197044 148300 197096 148352
rect 33376 147348 33428 147400
rect 34204 147348 34256 147400
rect 59228 146804 59280 146856
rect 59412 146736 59464 146788
rect 123076 146124 123128 146176
rect 123628 146124 123680 146176
rect 127216 146124 127268 146176
rect 127676 146124 127728 146176
rect 197596 146124 197648 146176
rect 198148 146124 198200 146176
rect 59412 144059 59464 144068
rect 59412 144025 59421 144059
rect 59421 144025 59455 144059
rect 59455 144025 59464 144059
rect 59412 144016 59464 144025
rect 118844 144016 118896 144068
rect 119580 144016 119632 144068
rect 120960 144016 121012 144068
rect 121696 144016 121748 144068
rect 123812 144016 123864 144068
rect 124548 144016 124600 144068
rect 125100 144016 125152 144068
rect 126020 144016 126072 144068
rect 127952 144016 128004 144068
rect 128596 144016 128648 144068
rect 129332 144016 129384 144068
rect 130068 144016 130120 144068
rect 183612 144016 183664 144068
rect 187936 144016 187988 144068
rect 198424 144016 198476 144068
rect 199068 144016 199120 144068
rect 201552 144016 201604 144068
rect 202196 144016 202248 144068
rect 203024 144016 203076 144068
rect 204496 144016 204548 144068
rect 207992 144016 208044 144068
rect 208728 144016 208780 144068
rect 210752 144016 210804 144068
rect 211396 144016 211448 144068
rect 21784 143948 21836 144000
rect 26016 143948 26068 144000
rect 41840 143948 41892 144000
rect 42300 143948 42352 144000
rect 123720 143948 123772 144000
rect 124456 143948 124508 144000
rect 125192 143948 125244 144000
rect 126572 143948 126624 144000
rect 127860 143948 127912 144000
rect 128688 143948 128740 144000
rect 129240 143948 129292 144000
rect 130620 143948 130672 144000
rect 183428 143948 183480 144000
rect 189408 143948 189460 144000
rect 198884 143948 198936 144000
rect 199252 143948 199304 144000
rect 201184 143948 201236 144000
rect 201736 143948 201788 144000
rect 202748 143948 202800 144000
rect 203852 143948 203904 144000
rect 207900 143948 207952 144000
rect 208636 143948 208688 144000
rect 210844 143948 210896 144000
rect 212316 143948 212368 144000
rect 117464 143880 117516 143932
rect 119028 143880 119080 143932
rect 183520 143880 183572 143932
rect 190052 143880 190104 143932
rect 202840 143880 202892 143932
rect 204956 143880 205008 143932
rect 210660 143880 210712 143932
rect 211764 143880 211816 143932
rect 38712 143812 38764 143864
rect 41840 143812 41892 143864
rect 183336 143812 183388 143864
rect 189500 143812 189552 143864
rect 201460 143812 201512 143864
rect 202748 143812 202800 143864
rect 210936 143812 210988 143864
rect 212960 143812 213012 143864
rect 201368 143744 201420 143796
rect 203300 143744 203352 143796
rect 24452 143676 24504 143728
rect 24912 143676 24964 143728
rect 23532 143608 23584 143660
rect 25740 143608 25792 143660
rect 26016 143608 26068 143660
rect 26292 143608 26344 143660
rect 27304 143608 27356 143660
rect 27764 143608 27816 143660
rect 28592 143608 28644 143660
rect 29144 143608 29196 143660
rect 30064 143608 30116 143660
rect 30524 143608 30576 143660
rect 31996 143608 32048 143660
rect 32732 143608 32784 143660
rect 34480 143608 34532 143660
rect 34940 143608 34992 143660
rect 35952 143608 36004 143660
rect 36228 143608 36280 143660
rect 37424 143608 37476 143660
rect 38988 143608 39040 143660
rect 43772 143608 43824 143660
rect 44416 143608 44468 143660
rect 110196 143608 110248 143660
rect 110472 143608 110524 143660
rect 112128 143608 112180 143660
rect 112588 143608 112640 143660
rect 114428 143608 114480 143660
rect 114980 143608 115032 143660
rect 115900 143608 115952 143660
rect 116636 143608 116688 143660
rect 192996 143608 193048 143660
rect 193272 143608 193324 143660
rect 194192 143608 194244 143660
rect 194652 143608 194704 143660
rect 20772 143540 20824 143592
rect 25096 143540 25148 143592
rect 34848 143540 34900 143592
rect 35492 143540 35544 143592
rect 35860 143540 35912 143592
rect 37516 143540 37568 143592
rect 43680 143540 43732 143592
rect 47176 143540 47228 143592
rect 99156 143540 99208 143592
rect 106700 143540 106752 143592
rect 114888 143540 114940 143592
rect 115532 143540 115584 143592
rect 116084 143540 116136 143592
rect 117648 143540 117700 143592
rect 99432 143472 99484 143524
rect 106608 143472 106660 143524
rect 113600 143472 113652 143524
rect 114428 143472 114480 143524
rect 183244 143472 183296 143524
rect 190788 143472 190840 143524
rect 38804 143404 38856 143456
rect 40276 143404 40328 143456
rect 99064 143404 99116 143456
rect 107436 143404 107488 143456
rect 183060 143404 183112 143456
rect 192076 143404 192128 143456
rect 22152 143336 22204 143388
rect 25832 143336 25884 143388
rect 20496 143268 20548 143320
rect 44508 143336 44560 143388
rect 98972 143336 99024 143388
rect 107988 143336 108040 143388
rect 183152 143336 183204 143388
rect 191340 143336 191392 143388
rect 191984 143336 192036 143388
rect 215628 143336 215680 143388
rect 37240 143200 37292 143252
rect 39724 143200 39776 143252
rect 45152 143200 45204 143252
rect 46532 143200 46584 143252
rect 35676 143064 35728 143116
rect 36964 143064 37016 143116
rect 117372 143064 117424 143116
rect 118476 143064 118528 143116
rect 31352 142928 31404 142980
rect 31904 142928 31956 142980
rect 38620 142928 38672 142980
rect 41012 142928 41064 142980
rect 45060 142928 45112 142980
rect 45796 142928 45848 142980
rect 98788 142928 98840 142980
rect 103940 142928 103992 142980
rect 117188 142928 117240 142980
rect 117924 142928 117976 142980
rect 99248 142860 99300 142912
rect 105596 142860 105648 142912
rect 23256 142792 23308 142844
rect 25924 142792 25976 142844
rect 37332 142792 37384 142844
rect 38252 142792 38304 142844
rect 99340 142792 99392 142844
rect 105136 142792 105188 142844
rect 200264 142792 200316 142844
rect 200908 142792 200960 142844
rect 99524 142724 99576 142776
rect 104492 142724 104544 142776
rect 68704 142656 68756 142708
rect 69164 142656 69216 142708
rect 167696 142452 167748 142504
rect 169904 142452 169956 142504
rect 49936 140412 49988 140464
rect 53340 140412 53392 140464
rect 134852 140004 134904 140056
rect 143592 140004 143644 140056
rect 49936 139936 49988 139988
rect 58492 139936 58544 139988
rect 135404 139936 135456 139988
rect 143316 139936 143368 139988
rect 135404 138712 135456 138764
rect 139820 138712 139872 138764
rect 49936 138576 49988 138628
rect 58400 138576 58452 138628
rect 134668 138576 134720 138628
rect 139636 138576 139688 138628
rect 92716 138508 92768 138560
rect 100812 138508 100864 138560
rect 177632 138508 177684 138560
rect 185084 138508 185136 138560
rect 49660 138440 49712 138492
rect 58952 138440 59004 138492
rect 92808 138440 92860 138492
rect 100904 138440 100956 138492
rect 177724 138440 177776 138492
rect 184992 138440 185044 138492
rect 97408 137420 97460 137472
rect 101824 137420 101876 137472
rect 134668 137352 134720 137404
rect 139728 137352 139780 137404
rect 49936 137216 49988 137268
rect 58308 137216 58360 137268
rect 98052 137216 98104 137268
rect 101272 137216 101324 137268
rect 181588 137216 181640 137268
rect 185176 137216 185228 137268
rect 50028 137148 50080 137200
rect 58216 137148 58268 137200
rect 135404 137148 135456 137200
rect 143408 137148 143460 137200
rect 182232 137148 182284 137200
rect 185452 137148 185504 137200
rect 92716 137080 92768 137132
rect 101180 137080 101232 137132
rect 177724 137080 177776 137132
rect 185360 137080 185412 137132
rect 92808 137012 92860 137064
rect 101088 137012 101140 137064
rect 139636 137012 139688 137064
rect 143592 137012 143644 137064
rect 177632 137012 177684 137064
rect 185268 137012 185320 137064
rect 92716 136944 92768 136996
rect 97408 136944 97460 136996
rect 139820 136944 139872 136996
rect 143132 136944 143184 136996
rect 139728 136604 139780 136656
rect 143500 136604 143552 136656
rect 177724 136604 177776 136656
rect 181588 136604 181640 136656
rect 51224 135924 51276 135976
rect 56652 135924 56704 135976
rect 135036 135924 135088 135976
rect 143316 135924 143368 135976
rect 51132 135856 51184 135908
rect 56744 135856 56796 135908
rect 97960 135856 98012 135908
rect 101272 135856 101324 135908
rect 135312 135856 135364 135908
rect 143592 135856 143644 135908
rect 182324 135856 182376 135908
rect 185360 135856 185412 135908
rect 51040 135788 51092 135840
rect 56560 135788 56612 135840
rect 98144 135788 98196 135840
rect 101732 135788 101784 135840
rect 135404 135788 135456 135840
rect 143224 135788 143276 135840
rect 181956 135788 182008 135840
rect 185268 135788 185320 135840
rect 92808 135720 92860 135772
rect 101180 135720 101232 135772
rect 177632 135720 177684 135772
rect 185176 135720 185228 135772
rect 92716 135652 92768 135704
rect 98052 135652 98104 135704
rect 177724 135652 177776 135704
rect 182232 135652 182284 135704
rect 56560 135584 56612 135636
rect 58216 135584 58268 135636
rect 56744 135312 56796 135364
rect 58308 135312 58360 135364
rect 134484 134632 134536 134684
rect 136876 134632 136928 134684
rect 51132 134496 51184 134548
rect 59412 134539 59464 134548
rect 51224 134428 51276 134480
rect 56100 134428 56152 134480
rect 59412 134505 59421 134539
rect 59421 134505 59455 134539
rect 59455 134505 59464 134539
rect 59412 134496 59464 134505
rect 134852 134496 134904 134548
rect 139636 134496 139688 134548
rect 58216 134360 58268 134412
rect 92900 134360 92952 134412
rect 101824 134360 101876 134412
rect 177632 134360 177684 134412
rect 185176 134360 185228 134412
rect 92808 134292 92860 134344
rect 98144 134292 98196 134344
rect 177724 134292 177776 134344
rect 181956 134292 182008 134344
rect 56652 134224 56704 134276
rect 58400 134224 58452 134276
rect 92716 134224 92768 134276
rect 97960 134224 98012 134276
rect 177724 134020 177776 134072
rect 182324 134020 182376 134072
rect 139636 133748 139688 133800
rect 142948 133748 143000 133800
rect 56100 133680 56152 133732
rect 58308 133680 58360 133732
rect 50396 133272 50448 133324
rect 56744 133272 56796 133324
rect 51224 133068 51276 133120
rect 55548 133068 55600 133120
rect 135036 133068 135088 133120
rect 138164 133068 138216 133120
rect 51132 133000 51184 133052
rect 135404 133000 135456 133052
rect 58216 132932 58268 132984
rect 59412 132932 59464 132984
rect 92808 132932 92860 132984
rect 101364 132932 101416 132984
rect 143224 132932 143276 132984
rect 177632 132932 177684 132984
rect 185176 132932 185228 132984
rect 56744 132864 56796 132916
rect 58308 132864 58360 132916
rect 92716 132864 92768 132916
rect 100904 132864 100956 132916
rect 177724 132864 177776 132916
rect 185084 132864 185136 132916
rect 136876 132796 136928 132848
rect 143592 132796 143644 132848
rect 135404 131980 135456 132032
rect 138072 131980 138124 132032
rect 135036 131776 135088 131828
rect 137336 131776 137388 131828
rect 51132 131708 51184 131760
rect 55456 131708 55508 131760
rect 51224 131640 51276 131692
rect 58492 131640 58544 131692
rect 135312 131640 135364 131692
rect 92808 131572 92860 131624
rect 101824 131572 101876 131624
rect 142488 131572 142540 131624
rect 177632 131572 177684 131624
rect 185452 131572 185504 131624
rect 92716 131504 92768 131556
rect 101732 131504 101784 131556
rect 138164 131504 138216 131556
rect 143592 131504 143644 131556
rect 177724 131504 177776 131556
rect 185820 131504 185872 131556
rect 55548 131368 55600 131420
rect 58216 131368 58268 131420
rect 55456 131096 55508 131148
rect 58308 131096 58360 131148
rect 135404 130552 135456 130604
rect 137612 130552 137664 130604
rect 51132 130416 51184 130468
rect 56744 130416 56796 130468
rect 51224 130348 51276 130400
rect 56560 130348 56612 130400
rect 50212 130280 50264 130332
rect 135036 130280 135088 130332
rect 137336 130280 137388 130332
rect 92808 130212 92860 130264
rect 101640 130212 101692 130264
rect 138072 130212 138124 130264
rect 143592 130212 143644 130264
rect 177632 130212 177684 130264
rect 185544 130212 185596 130264
rect 58216 130144 58268 130196
rect 92716 130144 92768 130196
rect 101456 130144 101508 130196
rect 137244 130144 137296 130196
rect 143040 130144 143092 130196
rect 177724 130144 177776 130196
rect 185728 130144 185780 130196
rect 135312 129328 135364 129380
rect 137704 129328 137756 129380
rect 51224 128988 51276 129040
rect 56652 128988 56704 129040
rect 51132 128920 51184 128972
rect 56376 128920 56428 128972
rect 135404 128920 135456 128972
rect 92900 128852 92952 128904
rect 101364 128852 101416 128904
rect 143132 128852 143184 128904
rect 177724 128852 177776 128904
rect 185268 128852 185320 128904
rect 56744 128784 56796 128836
rect 58216 128784 58268 128836
rect 92808 128784 92860 128836
rect 101824 128784 101876 128836
rect 137336 128784 137388 128836
rect 142764 128784 142816 128836
rect 177816 128784 177868 128836
rect 185176 128784 185228 128836
rect 56560 128716 56612 128768
rect 58400 128716 58452 128768
rect 92716 128716 92768 128768
rect 101732 128716 101784 128768
rect 137612 128716 137664 128768
rect 143592 128716 143644 128768
rect 177632 128716 177684 128768
rect 185360 128716 185412 128768
rect 56376 128512 56428 128564
rect 58308 128512 58360 128564
rect 135312 127696 135364 127748
rect 137612 127696 137664 127748
rect 50764 127560 50816 127612
rect 58216 127560 58268 127612
rect 134668 127560 134720 127612
rect 137428 127560 137480 127612
rect 51224 127492 51276 127544
rect 58308 127492 58360 127544
rect 135404 127492 135456 127544
rect 56652 127424 56704 127476
rect 58400 127424 58452 127476
rect 92808 127424 92860 127476
rect 100996 127424 101048 127476
rect 143316 127424 143368 127476
rect 177724 127424 177776 127476
rect 185176 127424 185228 127476
rect 216180 127424 216232 127476
rect 222344 127424 222396 127476
rect 92716 127356 92768 127408
rect 101272 127356 101324 127408
rect 137704 127356 137756 127408
rect 142488 127356 142540 127408
rect 177172 127356 177224 127408
rect 185452 127356 185504 127408
rect 50396 126336 50448 126388
rect 56744 126336 56796 126388
rect 51224 126200 51276 126252
rect 56100 126200 56152 126252
rect 98052 126200 98104 126252
rect 101272 126200 101324 126252
rect 182232 126200 182284 126252
rect 185452 126200 185504 126252
rect 50212 126132 50264 126184
rect 58216 126132 58268 126184
rect 98144 126132 98196 126184
rect 100996 126132 101048 126184
rect 182324 126132 182376 126184
rect 185176 126132 185228 126184
rect 92716 126064 92768 126116
rect 101180 126064 101232 126116
rect 137612 126064 137664 126116
rect 143500 126064 143552 126116
rect 177724 126064 177776 126116
rect 185360 126064 185412 126116
rect 92808 125996 92860 126048
rect 101088 125996 101140 126048
rect 137428 125996 137480 126048
rect 143592 125996 143644 126048
rect 177632 125996 177684 126048
rect 185268 125996 185320 126048
rect 135404 125384 135456 125436
rect 137612 125384 137664 125436
rect 51132 124840 51184 124892
rect 55456 124840 55508 124892
rect 135404 124840 135456 124892
rect 136876 124840 136928 124892
rect 51224 124772 51276 124824
rect 58400 124772 58452 124824
rect 135220 124772 135272 124824
rect 142764 124772 142816 124824
rect 55456 124704 55508 124756
rect 58216 124704 58268 124756
rect 92900 124704 92952 124756
rect 100996 124704 101048 124756
rect 135588 124704 135640 124756
rect 143592 124704 143644 124756
rect 177632 124704 177684 124756
rect 185176 124704 185228 124756
rect 56744 124636 56796 124688
rect 58308 124636 58360 124688
rect 92716 124636 92768 124688
rect 98052 124636 98104 124688
rect 177724 124636 177776 124688
rect 182232 124636 182284 124688
rect 56100 124568 56152 124620
rect 58492 124568 58544 124620
rect 92808 124568 92860 124620
rect 98144 124568 98196 124620
rect 135496 124364 135548 124416
rect 142488 124364 142540 124416
rect 177172 124364 177224 124416
rect 182324 124364 182376 124416
rect 51224 123616 51276 123668
rect 55548 123616 55600 123668
rect 135036 123616 135088 123668
rect 137428 123616 137480 123668
rect 51224 123480 51276 123532
rect 55456 123480 55508 123532
rect 50212 123344 50264 123396
rect 134116 123344 134168 123396
rect 138164 123344 138216 123396
rect 92808 123276 92860 123328
rect 101088 123276 101140 123328
rect 137612 123276 137664 123328
rect 143592 123276 143644 123328
rect 177632 123276 177684 123328
rect 185360 123276 185412 123328
rect 58216 123208 58268 123260
rect 92716 123208 92768 123260
rect 101272 123208 101324 123260
rect 177724 123208 177776 123260
rect 185452 123208 185504 123260
rect 136876 122800 136928 122852
rect 143592 122800 143644 122852
rect 135220 122528 135272 122580
rect 137888 122528 137940 122580
rect 135220 122188 135272 122240
rect 137796 122188 137848 122240
rect 51224 122120 51276 122172
rect 55732 122120 55784 122172
rect 51132 121984 51184 122036
rect 55640 121984 55692 122036
rect 92808 121916 92860 121968
rect 100996 121916 101048 121968
rect 137428 121916 137480 121968
rect 142764 121916 142816 121968
rect 177724 121916 177776 121968
rect 185820 121916 185872 121968
rect 92716 121848 92768 121900
rect 101180 121848 101232 121900
rect 138164 121848 138216 121900
rect 143040 121848 143092 121900
rect 177356 121848 177408 121900
rect 185268 121848 185320 121900
rect 55548 121780 55600 121832
rect 58216 121780 58268 121832
rect 55456 121508 55508 121560
rect 58216 121508 58268 121560
rect 97500 120760 97552 120812
rect 100996 120760 101048 120812
rect 134852 120760 134904 120812
rect 137336 120760 137388 120812
rect 182048 120760 182100 120812
rect 185360 120760 185412 120812
rect 51224 120692 51276 120744
rect 58492 120692 58544 120744
rect 97960 120692 98012 120744
rect 101180 120692 101232 120744
rect 134668 120692 134720 120744
rect 137612 120692 137664 120744
rect 182324 120692 182376 120744
rect 185268 120692 185320 120744
rect 51132 120624 51184 120676
rect 58308 120624 58360 120676
rect 98144 120624 98196 120676
rect 100996 120624 101048 120676
rect 135404 120624 135456 120676
rect 136876 120624 136928 120676
rect 181588 120624 181640 120676
rect 185176 120624 185228 120676
rect 55640 120556 55692 120608
rect 58216 120556 58268 120608
rect 92808 120556 92860 120608
rect 101088 120556 101140 120608
rect 137888 120556 137940 120608
rect 142948 120556 143000 120608
rect 177632 120556 177684 120608
rect 185912 120556 185964 120608
rect 55732 120488 55784 120540
rect 58400 120488 58452 120540
rect 92716 120488 92768 120540
rect 101272 120488 101324 120540
rect 137796 120488 137848 120540
rect 143592 120488 143644 120540
rect 177724 120488 177776 120540
rect 185636 120488 185688 120540
rect 134300 120080 134352 120132
rect 136968 120080 137020 120132
rect 51224 119536 51276 119588
rect 56744 119536 56796 119588
rect 135404 119536 135456 119588
rect 137704 119536 137756 119588
rect 51224 119400 51276 119452
rect 56284 119400 56336 119452
rect 97868 119332 97920 119384
rect 101088 119332 101140 119384
rect 182140 119332 182192 119384
rect 185268 119332 185320 119384
rect 50212 119264 50264 119316
rect 98052 119264 98104 119316
rect 100996 119264 101048 119316
rect 182232 119264 182284 119316
rect 185176 119264 185228 119316
rect 92900 119196 92952 119248
rect 98144 119196 98196 119248
rect 137336 119196 137388 119248
rect 143592 119196 143644 119248
rect 58216 119128 58268 119180
rect 92808 119128 92860 119180
rect 97960 119128 98012 119180
rect 137612 119128 137664 119180
rect 143040 119128 143092 119180
rect 92716 119060 92768 119112
rect 97500 119060 97552 119112
rect 136876 119060 136928 119112
rect 143316 119060 143368 119112
rect 177724 119060 177776 119112
rect 182048 119060 182100 119112
rect 177724 118924 177776 118976
rect 181588 118924 181640 118976
rect 177632 118788 177684 118840
rect 182324 118788 182376 118840
rect 134484 118176 134536 118228
rect 137612 118176 137664 118228
rect 51224 118040 51276 118092
rect 56560 118040 56612 118092
rect 50580 117904 50632 117956
rect 55548 117904 55600 117956
rect 97960 117904 98012 117956
rect 101088 117904 101140 117956
rect 134852 117904 134904 117956
rect 137428 117904 137480 117956
rect 182048 117904 182100 117956
rect 185268 117904 185320 117956
rect 98144 117836 98196 117888
rect 100996 117836 101048 117888
rect 182324 117836 182376 117888
rect 185176 117836 185228 117888
rect 56744 117768 56796 117820
rect 58216 117768 58268 117820
rect 92808 117768 92860 117820
rect 98052 117768 98104 117820
rect 136968 117768 137020 117820
rect 142580 117768 142632 117820
rect 56284 117700 56336 117752
rect 58308 117700 58360 117752
rect 92716 117700 92768 117752
rect 97868 117700 97920 117752
rect 137704 117700 137756 117752
rect 143224 117700 143276 117752
rect 177724 117700 177776 117752
rect 182140 117700 182192 117752
rect 177172 117428 177224 117480
rect 182232 117428 182284 117480
rect 94004 116544 94056 116596
rect 101088 116544 101140 116596
rect 178184 116544 178236 116596
rect 185268 116544 185320 116596
rect 50028 116476 50080 116528
rect 58216 116476 58268 116528
rect 92624 116476 92676 116528
rect 100996 116476 101048 116528
rect 134852 116476 134904 116528
rect 55548 116408 55600 116460
rect 58308 116408 58360 116460
rect 92900 116408 92952 116460
rect 101180 116408 101232 116460
rect 176804 116476 176856 116528
rect 185176 116476 185228 116528
rect 142764 116408 142816 116460
rect 177080 116408 177132 116460
rect 185360 116408 185412 116460
rect 56560 116340 56612 116392
rect 58400 116340 58452 116392
rect 92808 116340 92860 116392
rect 98144 116340 98196 116392
rect 137428 116340 137480 116392
rect 142948 116340 143000 116392
rect 177724 116340 177776 116392
rect 182048 116340 182100 116392
rect 92716 116272 92768 116324
rect 97960 116272 98012 116324
rect 137612 116272 137664 116324
rect 143592 116272 143644 116324
rect 177724 116068 177776 116120
rect 182324 116068 182376 116120
rect 91244 115184 91296 115236
rect 101088 115184 101140 115236
rect 175424 115184 175476 115236
rect 185268 115184 185320 115236
rect 59320 115159 59372 115168
rect 59320 115125 59329 115159
rect 59329 115125 59363 115159
rect 59363 115125 59372 115159
rect 59320 115116 59372 115125
rect 90600 115116 90652 115168
rect 100996 115116 101048 115168
rect 174780 115116 174832 115168
rect 185176 115116 185228 115168
rect 135404 113688 135456 113740
rect 141568 113688 141620 113740
rect 18012 113280 18064 113332
rect 64104 113280 64156 113332
rect 147272 113280 147324 113332
rect 218388 113280 218440 113332
rect 51224 112736 51276 112788
rect 54720 112736 54772 112788
rect 85724 112328 85776 112380
rect 100996 112328 101048 112380
rect 169904 112328 169956 112380
rect 185176 112328 185228 112380
rect 90416 112192 90468 112244
rect 93360 112192 93412 112244
rect 82320 111580 82372 111632
rect 85448 111580 85500 111632
rect 129976 111580 130028 111632
rect 148100 111580 148152 111632
rect 83700 111512 83752 111564
rect 87196 111512 87248 111564
rect 80940 111444 80992 111496
rect 84068 111444 84120 111496
rect 79560 111104 79612 111156
rect 82596 111104 82648 111156
rect 163832 111104 163884 111156
rect 166592 111104 166644 111156
rect 167880 111104 167932 111156
rect 170916 111104 170968 111156
rect 74040 111036 74092 111088
rect 75512 111036 75564 111088
rect 77444 111036 77496 111088
rect 79744 111036 79796 111088
rect 158864 111036 158916 111088
rect 160888 111036 160940 111088
rect 166500 111036 166552 111088
rect 169444 111036 169496 111088
rect 74684 110968 74736 111020
rect 76892 110968 76944 111020
rect 79652 110968 79704 111020
rect 81216 110968 81268 111020
rect 156840 110968 156892 111020
rect 158036 110968 158088 111020
rect 158312 110968 158364 111020
rect 159508 110968 159560 111020
rect 161624 110968 161676 111020
rect 163740 110968 163792 111020
rect 165120 110968 165172 111020
rect 168064 110968 168116 111020
rect 172664 110968 172716 111020
rect 176160 110968 176212 111020
rect 61436 110900 61488 110952
rect 108448 110900 108500 110952
rect 109000 110900 109052 110952
rect 129976 110900 130028 110952
rect 137520 110900 137572 110952
rect 145340 110900 145392 110952
rect 63276 110832 63328 110884
rect 109552 110832 109604 110884
rect 113140 110492 113192 110544
rect 114520 110492 114572 110544
rect 114612 110492 114664 110544
rect 115624 110492 115676 110544
rect 115992 110492 116044 110544
rect 117280 110492 117332 110544
rect 117464 110492 117516 110544
rect 118844 110492 118896 110544
rect 99524 110424 99576 110476
rect 107344 110424 107396 110476
rect 183612 110356 183664 110408
rect 191616 110356 191668 110408
rect 99432 110288 99484 110340
rect 106792 110288 106844 110340
rect 183704 110288 183756 110340
rect 192168 110288 192220 110340
rect 208268 110288 208320 110340
rect 213236 110288 213288 110340
rect 20220 110220 20272 110272
rect 41748 110220 41800 110272
rect 53340 110220 53392 110272
rect 61436 110220 61488 110272
rect 98788 110220 98840 110272
rect 107896 110220 107948 110272
rect 108448 110220 108500 110272
rect 133380 110220 133432 110272
rect 137520 110220 137572 110272
rect 183520 110220 183572 110272
rect 191064 110220 191116 110272
rect 191984 110220 192036 110272
rect 215536 110220 215588 110272
rect 113048 110152 113100 110204
rect 113968 110152 114020 110204
rect 115716 110152 115768 110204
rect 116728 110152 116780 110204
rect 115808 110016 115860 110068
rect 118292 110016 118344 110068
rect 25924 109948 25976 110000
rect 26292 109948 26344 110000
rect 29052 109948 29104 110000
rect 30892 109948 30944 110000
rect 24912 109880 24964 109932
rect 22888 109812 22940 109864
rect 27304 109812 27356 109864
rect 27672 109880 27724 109932
rect 30064 109880 30116 109932
rect 28500 109812 28552 109864
rect 99248 109812 99300 109864
rect 106240 109812 106292 109864
rect 119764 109812 119816 109864
rect 121604 109812 121656 109864
rect 183336 109812 183388 109864
rect 190420 109812 190472 109864
rect 203760 109812 203812 109864
rect 205324 109812 205376 109864
rect 23624 109744 23676 109796
rect 27672 109744 27724 109796
rect 99156 109744 99208 109796
rect 105688 109744 105740 109796
rect 118936 109744 118988 109796
rect 119948 109744 120000 109796
rect 126664 109744 126716 109796
rect 129332 109744 129384 109796
rect 183244 109744 183296 109796
rect 189868 109744 189920 109796
rect 21508 109676 21560 109728
rect 26476 109676 26528 109728
rect 42944 109676 42996 109728
rect 47452 109676 47504 109728
rect 99064 109676 99116 109728
rect 104584 109676 104636 109728
rect 115900 109676 115952 109728
rect 117832 109676 117884 109728
rect 119580 109676 119632 109728
rect 121052 109676 121104 109728
rect 183152 109676 183204 109728
rect 188764 109676 188816 109728
rect 205324 109676 205376 109728
rect 206428 109676 206480 109728
rect 208176 109676 208228 109728
rect 212132 109676 212184 109728
rect 22244 109608 22296 109660
rect 26568 109608 26620 109660
rect 27028 109608 27080 109660
rect 29696 109608 29748 109660
rect 38252 109608 38304 109660
rect 40000 109608 40052 109660
rect 45060 109608 45112 109660
rect 46808 109608 46860 109660
rect 98972 109608 99024 109660
rect 104124 109608 104176 109660
rect 119948 109608 120000 109660
rect 122156 109608 122208 109660
rect 126572 109608 126624 109660
rect 128780 109608 128832 109660
rect 129332 109608 129384 109660
rect 130988 109608 131040 109660
rect 183060 109608 183112 109660
rect 188212 109608 188264 109660
rect 201460 109608 201512 109660
rect 203024 109608 203076 109660
rect 205140 109608 205192 109660
rect 205876 109608 205928 109660
rect 208544 109608 208596 109660
rect 212684 109608 212736 109660
rect 213512 109608 213564 109660
rect 214984 109608 215036 109660
rect 20864 109540 20916 109592
rect 22980 109540 23032 109592
rect 24268 109540 24320 109592
rect 28132 109540 28184 109592
rect 28316 109540 28368 109592
rect 29144 109540 29196 109592
rect 31076 109540 31128 109592
rect 31812 109540 31864 109592
rect 38160 109540 38212 109592
rect 39264 109540 39316 109592
rect 45152 109540 45204 109592
rect 46072 109540 46124 109592
rect 99340 109540 99392 109592
rect 105136 109540 105188 109592
rect 119856 109540 119908 109592
rect 120500 109540 120552 109592
rect 120960 109540 121012 109592
rect 122708 109540 122760 109592
rect 126480 109540 126532 109592
rect 128228 109540 128280 109592
rect 129240 109540 129292 109592
rect 130436 109540 130488 109592
rect 183428 109540 183480 109592
rect 189316 109540 189368 109592
rect 193916 109540 193968 109592
rect 194744 109540 194796 109592
rect 201644 109540 201696 109592
rect 202472 109540 202524 109592
rect 203852 109540 203904 109592
rect 204680 109540 204732 109592
rect 205416 109540 205468 109592
rect 206980 109540 207032 109592
rect 208360 109540 208412 109592
rect 211580 109540 211632 109592
rect 213420 109540 213472 109592
rect 214432 109540 214484 109592
rect 59320 108180 59372 108232
rect 59412 108112 59464 108164
rect 208636 107500 208688 107552
rect 209556 107500 209608 107552
rect 210016 107500 210068 107552
rect 210660 107500 210712 107552
rect 194928 102672 194980 102724
rect 195112 102672 195164 102724
rect 199068 102672 199120 102724
rect 30248 102604 30300 102656
rect 31260 102604 31312 102656
rect 31996 102604 32048 102656
rect 32824 102604 32876 102656
rect 33468 102604 33520 102656
rect 34112 102604 34164 102656
rect 35124 102604 35176 102656
rect 35492 102604 35544 102656
rect 35676 102604 35728 102656
rect 36596 102604 36648 102656
rect 37700 102604 37752 102656
rect 40276 102604 40328 102656
rect 54720 102604 54772 102656
rect 56468 102604 56520 102656
rect 111300 102604 111352 102656
rect 111760 102604 111812 102656
rect 112496 102604 112548 102656
rect 113324 102604 113376 102656
rect 113692 102604 113744 102656
rect 114704 102604 114756 102656
rect 115624 102604 115676 102656
rect 115900 102604 115952 102656
rect 193272 102604 193324 102656
rect 194100 102604 194152 102656
rect 196308 102604 196360 102656
rect 196860 102604 196912 102656
rect 198424 102604 198476 102656
rect 199620 102604 199672 102656
rect 200356 102604 200408 102656
rect 200816 102604 200868 102656
rect 201644 102604 201696 102656
rect 202840 102604 202892 102656
rect 203760 102604 203812 102656
rect 204864 102604 204916 102656
rect 207348 102604 207400 102656
rect 32088 102536 32140 102588
rect 33284 102536 33336 102588
rect 36504 102536 36556 102588
rect 38068 102536 38120 102588
rect 111668 102536 111720 102588
rect 112312 102536 112364 102588
rect 114060 102536 114112 102588
rect 114612 102536 114664 102588
rect 114888 102536 114940 102588
rect 115716 102536 115768 102588
rect 199252 102536 199304 102588
rect 199712 102536 199764 102588
rect 202472 102536 202524 102588
rect 203852 102536 203904 102588
rect 204036 102536 204088 102588
rect 205416 102536 205468 102588
rect 115256 102468 115308 102520
rect 115992 102468 116044 102520
rect 120500 102468 120552 102520
rect 124364 102468 124416 102520
rect 201644 102468 201696 102520
rect 203116 102468 203168 102520
rect 203300 102468 203352 102520
rect 205140 102468 205192 102520
rect 22980 102400 23032 102452
rect 26108 102400 26160 102452
rect 36872 102400 36924 102452
rect 38160 102400 38212 102452
rect 50948 102400 51000 102452
rect 57572 102400 57624 102452
rect 93360 102400 93412 102452
rect 94188 102400 94240 102452
rect 120040 102400 120092 102452
rect 123812 102400 123864 102452
rect 205232 102400 205284 102452
rect 208820 102400 208872 102452
rect 38068 102332 38120 102384
rect 40828 102332 40880 102384
rect 51132 102332 51184 102384
rect 59780 102332 59832 102384
rect 119672 102332 119724 102384
rect 123260 102332 123312 102384
rect 135128 102332 135180 102384
rect 143776 102332 143828 102384
rect 206428 102332 206480 102384
rect 210108 102332 210160 102384
rect 143684 102264 143736 102316
rect 167144 102264 167196 102316
rect 50856 102196 50908 102248
rect 60884 102196 60936 102248
rect 114428 102196 114480 102248
rect 116176 102196 116228 102248
rect 122432 102196 122484 102248
rect 127124 102196 127176 102248
rect 135036 102196 135088 102248
rect 144880 102196 144932 102248
rect 208820 102196 208872 102248
rect 212868 102196 212920 102248
rect 50672 102128 50724 102180
rect 61988 102128 62040 102180
rect 121696 102128 121748 102180
rect 126020 102128 126072 102180
rect 134852 102128 134904 102180
rect 145984 102128 146036 102180
rect 203668 102128 203720 102180
rect 205324 102128 205376 102180
rect 50764 102060 50816 102112
rect 63092 102060 63144 102112
rect 88668 102060 88720 102112
rect 102008 102060 102060 102112
rect 122892 102060 122944 102112
rect 127676 102060 127728 102112
rect 134760 102060 134812 102112
rect 147088 102060 147140 102112
rect 172664 102060 172716 102112
rect 186004 102060 186056 102112
rect 209280 102060 209332 102112
rect 213420 102060 213472 102112
rect 26292 101992 26344 102044
rect 28868 101992 28920 102044
rect 29144 101992 29196 102044
rect 30432 101992 30484 102044
rect 37240 101992 37292 102044
rect 38252 101992 38304 102044
rect 41656 101992 41708 102044
rect 42944 101992 42996 102044
rect 50580 101992 50632 102044
rect 64196 101992 64248 102044
rect 87564 101992 87616 102044
rect 101640 101992 101692 102044
rect 122064 101992 122116 102044
rect 126112 101992 126164 102044
rect 134944 101992 134996 102044
rect 148192 101992 148244 102044
rect 161532 101992 161584 102044
rect 164476 101992 164528 102044
rect 171560 101992 171612 102044
rect 185820 101992 185872 102044
rect 202104 101992 202156 102044
rect 203208 101992 203260 102044
rect 50488 101924 50540 101976
rect 58676 101924 58728 101976
rect 59412 101924 59464 101976
rect 83148 101924 83200 101976
rect 86460 101924 86512 101976
rect 101824 101924 101876 101976
rect 112036 101924 112088 101976
rect 112864 101924 112916 101976
rect 121236 101924 121288 101976
rect 125468 101924 125520 101976
rect 135312 101924 135364 101976
rect 142672 101924 142724 101976
rect 170456 101924 170508 101976
rect 186188 101924 186240 101976
rect 209648 101924 209700 101976
rect 213512 101924 213564 101976
rect 40092 101856 40144 101908
rect 44416 101856 44468 101908
rect 200448 101856 200500 101908
rect 201552 101856 201604 101908
rect 30524 101788 30576 101840
rect 31628 101788 31680 101840
rect 40828 101788 40880 101840
rect 45152 101788 45204 101840
rect 116452 101788 116504 101840
rect 117464 101788 117516 101840
rect 124456 101788 124508 101840
rect 129884 101788 129936 101840
rect 206888 101788 206940 101840
rect 210016 101788 210068 101840
rect 26384 101720 26436 101772
rect 29236 101720 29288 101772
rect 39632 101720 39684 101772
rect 43588 101720 43640 101772
rect 120868 101720 120920 101772
rect 124916 101720 124968 101772
rect 35308 101652 35360 101704
rect 36136 101652 36188 101704
rect 39264 101652 39316 101704
rect 43036 101652 43088 101704
rect 117648 101652 117700 101704
rect 119856 101652 119908 101704
rect 123260 101652 123312 101704
rect 126480 101652 126532 101704
rect 204496 101652 204548 101704
rect 207256 101652 207308 101704
rect 36044 101584 36096 101636
rect 37516 101584 37568 101636
rect 38436 101584 38488 101636
rect 41840 101584 41892 101636
rect 116820 101584 116872 101636
rect 119396 101584 119448 101636
rect 123628 101584 123680 101636
rect 126572 101584 126624 101636
rect 159324 101584 159376 101636
rect 161716 101584 161768 101636
rect 205692 101584 205744 101636
rect 208912 101584 208964 101636
rect 40460 101516 40512 101568
rect 44876 101516 44928 101568
rect 75328 101516 75380 101568
rect 77536 101516 77588 101568
rect 118844 101516 118896 101568
rect 119948 101516 120000 101568
rect 124824 101516 124876 101568
rect 129240 101516 129292 101568
rect 207624 101516 207676 101568
rect 208176 101516 208228 101568
rect 38896 101448 38948 101500
rect 42300 101448 42352 101500
rect 118476 101448 118528 101500
rect 119764 101448 119816 101500
rect 124088 101448 124140 101500
rect 126664 101448 126716 101500
rect 206060 101448 206112 101500
rect 208636 101448 208688 101500
rect 41288 101380 41340 101432
rect 45060 101380 45112 101432
rect 72384 101380 72436 101432
rect 73488 101380 73540 101432
rect 77536 101380 77588 101432
rect 79652 101380 79704 101432
rect 80848 101380 80900 101432
rect 82320 101380 82372 101432
rect 117280 101380 117332 101432
rect 118936 101380 118988 101432
rect 119304 101380 119356 101432
rect 120960 101380 121012 101432
rect 125652 101380 125704 101432
rect 131540 101380 131592 101432
rect 154908 101380 154960 101432
rect 156196 101380 156248 101432
rect 158220 101380 158272 101432
rect 158864 101380 158916 101432
rect 163740 101380 163792 101432
rect 165120 101380 165172 101432
rect 165948 101380 166000 101432
rect 167880 101380 167932 101432
rect 176160 101380 176212 101432
rect 179288 101380 179340 101432
rect 193364 101380 193416 101432
rect 194468 101380 194520 101432
rect 207256 101380 207308 101432
rect 208360 101380 208412 101432
rect 68612 101312 68664 101364
rect 69256 101312 69308 101364
rect 69808 101312 69860 101364
rect 70636 101312 70688 101364
rect 70912 101312 70964 101364
rect 72016 101312 72068 101364
rect 73120 101312 73172 101364
rect 74040 101312 74092 101364
rect 76432 101312 76484 101364
rect 77444 101312 77496 101364
rect 78640 101312 78692 101364
rect 79560 101312 79612 101364
rect 79744 101312 79796 101364
rect 80940 101312 80992 101364
rect 81952 101312 82004 101364
rect 83700 101312 83752 101364
rect 89772 101312 89824 101364
rect 90600 101312 90652 101364
rect 91980 101312 92032 101364
rect 92624 101312 92676 101364
rect 93084 101312 93136 101364
rect 94004 101312 94056 101364
rect 118108 101312 118160 101364
rect 119580 101312 119632 101364
rect 125284 101312 125336 101364
rect 129332 101312 129384 101364
rect 135220 101312 135272 101364
rect 140464 101312 140516 101364
rect 152608 101312 152660 101364
rect 153436 101312 153488 101364
rect 153804 101312 153856 101364
rect 154816 101312 154868 101364
rect 156012 101312 156064 101364
rect 156840 101312 156892 101364
rect 157116 101312 157168 101364
rect 158312 101312 158364 101364
rect 160428 101312 160480 101364
rect 161624 101312 161676 101364
rect 162636 101312 162688 101364
rect 163832 101312 163884 101364
rect 164844 101312 164896 101364
rect 166500 101312 166552 101364
rect 173768 101312 173820 101364
rect 174780 101312 174832 101364
rect 175976 101312 176028 101364
rect 176804 101312 176856 101364
rect 177080 101312 177132 101364
rect 178184 101312 178236 101364
rect 194652 101312 194704 101364
rect 194928 101312 194980 101364
rect 196032 101312 196084 101364
rect 208084 101312 208136 101364
rect 208544 101312 208596 101364
rect 194928 101176 194980 101228
rect 98788 97164 98840 97216
rect 106792 97164 106844 97216
rect 18104 97096 18156 97148
rect 22336 97096 22388 97148
rect 212316 97096 212368 97148
rect 220964 97096 221016 97148
rect 99524 95804 99576 95856
rect 106792 95804 106844 95856
rect 188580 94376 188632 94428
rect 191984 94376 192036 94428
rect 98696 93016 98748 93068
rect 106516 93016 106568 93068
rect 105044 90228 105096 90280
rect 106792 90228 106844 90280
rect 13320 90160 13372 90212
rect 22336 90160 22388 90212
rect 182876 90160 182928 90212
rect 188580 90160 188632 90212
rect 104952 88868 105004 88920
rect 106792 88868 106844 88920
rect 128504 88868 128556 88920
rect 132000 88868 132052 88920
rect 183520 88800 183572 88852
rect 191156 88800 191208 88852
rect 183704 87440 183756 87492
rect 190788 87440 190840 87492
rect 183704 86012 183756 86064
rect 191708 86012 191760 86064
rect 99524 85196 99576 85248
rect 105044 85196 105096 85248
rect 44416 84720 44468 84772
rect 52696 84720 52748 84772
rect 99432 84652 99484 84704
rect 106792 84652 106844 84704
rect 182508 84652 182560 84704
rect 191984 84652 192036 84704
rect 99524 84584 99576 84636
rect 104952 84584 105004 84636
rect 183704 84584 183756 84636
rect 191616 84584 191668 84636
rect 13412 83292 13464 83344
rect 22336 83292 22388 83344
rect 99524 83292 99576 83344
rect 107804 83292 107856 83344
rect 183704 82612 183756 82664
rect 191984 82612 192036 82664
rect 99524 81932 99576 81984
rect 106792 82068 106844 82120
rect 183244 81252 183296 81304
rect 191892 81252 191944 81304
rect 132000 80504 132052 80556
rect 136876 80504 136928 80556
rect 99524 79824 99576 79876
rect 106792 79824 106844 79876
rect 183704 79212 183756 79264
rect 191984 79144 192036 79196
rect 99524 77852 99576 77904
rect 106516 77852 106568 77904
rect 183520 77852 183572 77904
rect 191984 77852 192036 77904
rect 13504 77784 13556 77836
rect 22336 77784 22388 77836
rect 99524 76424 99576 76476
rect 100996 76424 101048 76476
rect 183060 76424 183112 76476
rect 185176 76424 185228 76476
rect 98236 75064 98288 75116
rect 183244 75064 183296 75116
rect 186188 75064 186240 75116
rect 100996 74996 101048 75048
rect 106792 74996 106844 75048
rect 185176 74996 185228 75048
rect 191524 74996 191576 75048
rect 212132 74996 212184 75048
rect 222344 74996 222396 75048
rect 100996 74860 101048 74912
rect 44416 74316 44468 74368
rect 53340 74316 53392 74368
rect 99524 73840 99576 73892
rect 105136 73840 105188 73892
rect 183704 73840 183756 73892
rect 99432 73704 99484 73756
rect 106700 73704 106752 73756
rect 183704 73704 183756 73756
rect 188488 73704 188540 73756
rect 190788 73704 190840 73756
rect 100996 73636 101048 73688
rect 106792 73636 106844 73688
rect 186188 73636 186240 73688
rect 191984 73636 192036 73688
rect 99524 72344 99576 72396
rect 106516 72344 106568 72396
rect 99524 70984 99576 71036
rect 104492 70984 104544 71036
rect 183704 70916 183756 70968
rect 191524 70916 191576 70968
rect 128504 70168 128556 70220
rect 133380 70168 133432 70220
rect 136876 70168 136928 70220
rect 182876 69896 182928 69948
rect 189960 69896 190012 69948
rect 212684 69760 212736 69812
rect 215628 69760 215680 69812
rect 99524 69556 99576 69608
rect 104400 69556 104452 69608
rect 188488 69488 188540 69540
rect 190972 69488 191024 69540
rect 105136 68128 105188 68180
rect 106608 68128 106660 68180
rect 183796 68128 183848 68180
rect 191340 68128 191392 68180
rect 104492 63640 104544 63692
rect 106608 63640 106660 63692
rect 183704 61464 183756 61516
rect 188028 61464 188080 61516
rect 99524 61328 99576 61380
rect 105320 61328 105372 61380
rect 104400 61192 104452 61244
rect 107160 61192 107212 61244
rect 182692 60376 182744 60428
rect 184440 60376 184492 60428
rect 26752 59968 26804 60020
rect 26936 59968 26988 60020
rect 137980 59832 138032 59884
rect 138164 59832 138216 59884
rect 112404 58540 112456 58592
rect 112864 58540 112916 58592
rect 36136 58472 36188 58524
rect 37608 58472 37660 58524
rect 79192 58472 79244 58524
rect 96120 58472 96172 58524
rect 163188 58472 163240 58524
rect 199620 58472 199672 58524
rect 200356 58472 200408 58524
rect 208084 58472 208136 58524
rect 210660 58472 210712 58524
rect 41288 58404 41340 58456
rect 45888 58404 45940 58456
rect 72568 58404 72620 58456
rect 98880 58404 98932 58456
rect 156564 58404 156616 58456
rect 209648 58404 209700 58456
rect 212316 58404 212368 58456
rect 41656 58336 41708 58388
rect 46440 58336 46492 58388
rect 121236 58336 121288 58388
rect 123720 58336 123772 58388
rect 207624 58336 207676 58388
rect 210752 58336 210804 58388
rect 122432 58268 122484 58320
rect 125100 58268 125152 58320
rect 208820 58268 208872 58320
rect 212224 58268 212276 58320
rect 123260 58200 123312 58252
rect 127308 58200 127360 58252
rect 207256 58200 207308 58252
rect 210844 58200 210896 58252
rect 120500 58064 120552 58116
rect 123260 58064 123312 58116
rect 209280 58064 209332 58116
rect 212132 58064 212184 58116
rect 120868 57928 120920 57980
rect 123444 57928 123496 57980
rect 70544 57860 70596 57912
rect 92532 57860 92584 57912
rect 13320 57792 13372 57844
rect 72568 57792 72620 57844
rect 122064 57792 122116 57844
rect 125192 57792 125244 57844
rect 156104 57792 156156 57844
rect 169904 57792 169956 57844
rect 208452 57792 208504 57844
rect 212868 57792 212920 57844
rect 40828 57724 40880 57776
rect 45796 57724 45848 57776
rect 114060 57724 114112 57776
rect 114980 57724 115032 57776
rect 116820 57656 116872 57708
rect 118384 57656 118436 57708
rect 125284 57656 125336 57708
rect 129976 57656 130028 57708
rect 116084 57588 116136 57640
rect 117740 57588 117792 57640
rect 206428 57588 206480 57640
rect 210108 57588 210160 57640
rect 40092 57520 40144 57572
rect 43772 57520 43824 57572
rect 118844 57520 118896 57572
rect 121236 57520 121288 57572
rect 122892 57520 122944 57572
rect 125284 57520 125336 57572
rect 204496 57520 204548 57572
rect 207256 57520 207308 57572
rect 39264 57452 39316 57504
rect 43036 57452 43088 57504
rect 118108 57452 118160 57504
rect 120500 57452 120552 57504
rect 124088 57452 124140 57504
rect 128780 57452 128832 57504
rect 205232 57452 205284 57504
rect 207992 57452 208044 57504
rect 39632 57384 39684 57436
rect 43128 57384 43180 57436
rect 118476 57384 118528 57436
rect 120776 57384 120828 57436
rect 121696 57384 121748 57436
rect 124916 57384 124968 57436
rect 203300 57384 203352 57436
rect 205324 57384 205376 57436
rect 206888 57384 206940 57436
rect 210016 57384 210068 57436
rect 29144 57316 29196 57368
rect 30432 57316 30484 57368
rect 37700 57316 37752 57368
rect 40276 57316 40328 57368
rect 124456 57316 124508 57368
rect 128872 57316 128924 57368
rect 200724 57316 200776 57368
rect 201828 57316 201880 57368
rect 202472 57316 202524 57368
rect 204588 57316 204640 57368
rect 204864 57316 204916 57368
rect 207348 57316 207400 57368
rect 36872 57248 36924 57300
rect 38252 57248 38304 57300
rect 38896 57248 38948 57300
rect 41840 57248 41892 57300
rect 115256 57248 115308 57300
rect 116268 57248 116320 57300
rect 117648 57248 117700 57300
rect 118844 57248 118896 57300
rect 119304 57248 119356 57300
rect 121052 57248 121104 57300
rect 123628 57248 123680 57300
rect 127216 57248 127268 57300
rect 194652 57248 194704 57300
rect 195296 57248 195348 57300
rect 198884 57248 198936 57300
rect 199160 57248 199212 57300
rect 201276 57248 201328 57300
rect 202196 57248 202248 57300
rect 203668 57248 203720 57300
rect 205232 57248 205284 57300
rect 30432 57180 30484 57232
rect 31260 57180 31312 57232
rect 37240 57180 37292 57232
rect 38160 57180 38212 57232
rect 38436 57180 38488 57232
rect 40920 57180 40972 57232
rect 109276 57180 109328 57232
rect 110472 57180 110524 57232
rect 114428 57180 114480 57232
rect 115348 57180 115400 57232
rect 116452 57180 116504 57232
rect 118108 57180 118160 57232
rect 120040 57180 120092 57232
rect 121144 57180 121196 57232
rect 124824 57180 124876 57232
rect 129516 57180 129568 57232
rect 193364 57180 193416 57232
rect 194468 57180 194520 57232
rect 195112 57180 195164 57232
rect 196032 57180 196084 57232
rect 196400 57180 196452 57232
rect 196860 57180 196912 57232
rect 201644 57180 201696 57232
rect 202380 57180 202432 57232
rect 202840 57180 202892 57232
rect 204496 57180 204548 57232
rect 205692 57180 205744 57232
rect 207900 57180 207952 57232
rect 26568 57112 26620 57164
rect 27028 57112 27080 57164
rect 27856 57112 27908 57164
rect 28592 57112 28644 57164
rect 29328 57112 29380 57164
rect 29604 57112 29656 57164
rect 30524 57112 30576 57164
rect 31628 57112 31680 57164
rect 26476 57044 26528 57096
rect 27396 57044 27448 57096
rect 29420 57044 29472 57096
rect 29788 57044 29840 57096
rect 33284 57112 33336 57164
rect 33468 57112 33520 57164
rect 34112 57112 34164 57164
rect 35308 57112 35360 57164
rect 36044 57112 36096 57164
rect 36504 57112 36556 57164
rect 37516 57112 37568 57164
rect 38068 57112 38120 57164
rect 40368 57112 40420 57164
rect 40460 57112 40512 57164
rect 43680 57112 43732 57164
rect 109184 57112 109236 57164
rect 110104 57112 110156 57164
rect 111116 57112 111168 57164
rect 111668 57112 111720 57164
rect 114888 57112 114940 57164
rect 115532 57112 115584 57164
rect 115992 57112 116044 57164
rect 116636 57112 116688 57164
rect 117280 57112 117332 57164
rect 118200 57112 118252 57164
rect 119672 57112 119724 57164
rect 120960 57112 121012 57164
rect 125652 57112 125704 57164
rect 130068 57112 130120 57164
rect 193272 57112 193324 57164
rect 194100 57112 194152 57164
rect 194928 57112 194980 57164
rect 195664 57112 195716 57164
rect 196308 57112 196360 57164
rect 197228 57112 197280 57164
rect 200816 57112 200868 57164
rect 201920 57112 201972 57164
rect 202104 57112 202156 57164
rect 203024 57112 203076 57164
rect 204036 57112 204088 57164
rect 205140 57112 205192 57164
rect 206060 57112 206112 57164
rect 207164 57112 207216 57164
rect 32088 56772 32140 56824
rect 138164 55684 138216 55736
rect 138348 55684 138400 55736
rect 194192 54324 194244 54376
rect 194744 54324 194796 54376
rect 198976 54324 199028 54376
rect 199252 54324 199304 54376
rect 210660 50516 210712 50568
rect 210936 50516 210988 50568
rect 127216 50380 127268 50432
rect 127860 50380 127912 50432
rect 196216 50380 196268 50432
rect 197044 50380 197096 50432
rect 197688 50380 197740 50432
rect 198148 50380 198200 50432
rect 199068 50380 199120 50432
rect 199804 50380 199856 50432
rect 204496 50380 204548 50432
rect 204956 50380 205008 50432
rect 210016 50380 210068 50432
rect 210660 50380 210712 50432
rect 212132 50312 212184 50364
rect 33468 50244 33520 50296
rect 34296 50244 34348 50296
rect 112312 50244 112364 50296
rect 112496 50244 112548 50296
rect 199068 50244 199120 50296
rect 199252 50244 199304 50296
rect 25648 50176 25700 50228
rect 27856 50176 27908 50228
rect 28316 50176 28368 50228
rect 29144 50176 29196 50228
rect 29696 50176 29748 50228
rect 30432 50176 30484 50228
rect 31076 50176 31128 50228
rect 31812 50176 31864 50228
rect 38252 50176 38304 50228
rect 39264 50176 39316 50228
rect 40920 50176 40972 50228
rect 42024 50176 42076 50228
rect 43772 50176 43824 50228
rect 44692 50176 44744 50228
rect 46440 50176 46492 50228
rect 47452 50176 47504 50228
rect 100260 50176 100312 50228
rect 104768 50176 104820 50228
rect 118200 50176 118252 50228
rect 119304 50176 119356 50228
rect 120960 50176 121012 50228
rect 122616 50176 122668 50228
rect 123720 50176 123772 50228
rect 124824 50176 124876 50228
rect 184440 50176 184492 50228
rect 188212 50176 188264 50228
rect 205324 50176 205376 50228
rect 205876 50176 205928 50228
rect 207992 50176 208044 50228
rect 208728 50176 208780 50228
rect 210752 50176 210804 50228
rect 212132 50176 212184 50228
rect 214432 50176 214484 50228
rect 29052 50108 29104 50160
rect 30708 50108 30760 50160
rect 38160 50108 38212 50160
rect 40000 50108 40052 50160
rect 99340 50108 99392 50160
rect 105872 50108 105924 50160
rect 205232 50108 205284 50160
rect 206428 50108 206480 50160
rect 207900 50108 207952 50160
rect 209280 50108 209332 50160
rect 210936 50108 210988 50160
rect 212684 50108 212736 50160
rect 22244 50040 22296 50092
rect 26660 50040 26712 50092
rect 37516 50040 37568 50092
rect 38252 50040 38304 50092
rect 99524 50040 99576 50092
rect 106424 50040 106476 50092
rect 121144 50040 121196 50092
rect 123168 50040 123220 50092
rect 202380 50040 202432 50092
rect 203576 50040 203628 50092
rect 205140 50040 205192 50092
rect 206980 50040 207032 50092
rect 21508 49972 21560 50024
rect 26936 49972 26988 50024
rect 125192 49904 125244 49956
rect 126020 49904 126072 49956
rect 20864 49836 20916 49888
rect 25096 49836 25148 49888
rect 23624 49700 23676 49752
rect 26476 49836 26528 49888
rect 24268 49632 24320 49684
rect 27948 49768 28000 49820
rect 43680 49768 43732 49820
rect 45428 49768 45480 49820
rect 99248 49768 99300 49820
rect 106976 49768 107028 49820
rect 26292 49700 26344 49752
rect 29512 49700 29564 49752
rect 121052 49700 121104 49752
rect 122064 49700 122116 49752
rect 99156 49632 99208 49684
rect 107528 49632 107580 49684
rect 183244 49632 183296 49684
rect 191064 49632 191116 49684
rect 212224 49632 212276 49684
rect 213880 49632 213932 49684
rect 99064 49564 99116 49616
rect 108080 49564 108132 49616
rect 183060 49564 183112 49616
rect 192168 49564 192220 49616
rect 20220 49496 20272 49548
rect 44416 49496 44468 49548
rect 98972 49496 99024 49548
rect 108632 49496 108684 49548
rect 125100 49496 125152 49548
rect 126572 49496 126624 49548
rect 183152 49496 183204 49548
rect 191616 49496 191668 49548
rect 191984 49496 192036 49548
rect 215536 49564 215588 49616
rect 210844 49496 210896 49548
rect 211580 49496 211632 49548
rect 212316 49496 212368 49548
rect 214984 49496 215036 49548
rect 24912 49360 24964 49412
rect 28040 49360 28092 49412
rect 183428 49292 183480 49344
rect 189316 49292 189368 49344
rect 22888 49224 22940 49276
rect 26568 49224 26620 49276
rect 27672 49224 27724 49276
rect 29420 49224 29472 49276
rect 183612 49224 183664 49276
rect 189868 49224 189920 49276
rect 125284 49156 125336 49208
rect 127124 49156 127176 49208
rect 207164 49156 207216 49208
rect 209832 49156 209884 49208
rect 118844 49088 118896 49140
rect 119856 49088 119908 49140
rect 183336 49088 183388 49140
rect 190420 49088 190472 49140
rect 203024 49088 203076 49140
rect 204128 49088 204180 49140
rect 27028 49020 27080 49072
rect 29328 49020 29380 49072
rect 36136 48884 36188 48936
rect 37240 48884 37292 48936
rect 90692 48884 90744 48936
rect 104216 48884 104268 48936
rect 212040 48816 212092 48868
rect 222252 48816 222304 48868
rect 50396 47048 50448 47100
rect 53340 47048 53392 47100
rect 110748 46912 110800 46964
rect 110932 46912 110984 46964
rect 134576 46504 134628 46556
rect 145340 46504 145392 46556
rect 50580 46436 50632 46488
rect 61344 46436 61396 46488
rect 134760 46436 134812 46488
rect 142580 46436 142632 46488
rect 50764 46368 50816 46420
rect 62816 46368 62868 46420
rect 135220 46368 135272 46420
rect 146812 46368 146864 46420
rect 50856 46300 50908 46352
rect 64288 46300 64340 46352
rect 135036 46300 135088 46352
rect 148284 46300 148336 46352
rect 51040 46232 51092 46284
rect 65760 46232 65812 46284
rect 82964 46232 83016 46284
rect 93360 46232 93412 46284
rect 134944 46232 134996 46284
rect 149756 46232 149808 46284
rect 50672 46164 50724 46216
rect 67324 46164 67376 46216
rect 84068 46164 84120 46216
rect 94740 46164 94792 46216
rect 135128 46164 135180 46216
rect 151320 46164 151372 46216
rect 168432 46164 168484 46216
rect 177540 46164 177592 46216
rect 50948 46096 51000 46148
rect 68796 46096 68848 46148
rect 88944 46096 88996 46148
rect 96120 46096 96172 46148
rect 135312 46096 135364 46148
rect 152792 46096 152844 46148
rect 166960 46096 167012 46148
rect 176160 46096 176212 46148
rect 181036 45280 181088 45332
rect 185176 45280 185228 45332
rect 134760 44872 134812 44924
rect 142672 44872 142724 44924
rect 134300 44804 134352 44856
rect 142488 44804 142540 44856
rect 51224 44736 51276 44788
rect 134852 44736 134904 44788
rect 58308 44668 58360 44720
rect 93912 44668 93964 44720
rect 100996 44668 101048 44720
rect 142396 44668 142448 44720
rect 177724 44668 177776 44720
rect 185820 44668 185872 44720
rect 51316 44600 51368 44652
rect 58216 44600 58268 44652
rect 94004 44600 94056 44652
rect 101180 44600 101232 44652
rect 90324 44532 90376 44584
rect 90416 44464 90468 44516
rect 90692 44464 90744 44516
rect 177724 43852 177776 43904
rect 181036 43852 181088 43904
rect 134760 43648 134812 43700
rect 139636 43648 139688 43700
rect 50028 43512 50080 43564
rect 56744 43512 56796 43564
rect 51224 43308 51276 43360
rect 56652 43308 56704 43360
rect 96856 43308 96908 43360
rect 100996 43308 101048 43360
rect 134760 43308 134812 43360
rect 143500 43308 143552 43360
rect 181772 43308 181824 43360
rect 185176 43308 185228 43360
rect 93912 43240 93964 43292
rect 101088 43240 101140 43292
rect 134944 43240 134996 43292
rect 135220 43240 135272 43292
rect 139636 43240 139688 43292
rect 143132 43240 143184 43292
rect 177724 43240 177776 43292
rect 185452 43240 185504 43292
rect 56652 43172 56704 43224
rect 58216 43172 58268 43224
rect 94004 43172 94056 43224
rect 101272 43172 101324 43224
rect 177632 43172 177684 43224
rect 185544 43172 185596 43224
rect 56744 43104 56796 43156
rect 58308 43104 58360 43156
rect 50212 42560 50264 42612
rect 58216 42560 58268 42612
rect 94004 42560 94056 42612
rect 96856 42560 96908 42612
rect 177724 42424 177776 42476
rect 181772 42424 181824 42476
rect 134760 42288 134812 42340
rect 139636 42288 139688 42340
rect 51132 42016 51184 42068
rect 51224 41948 51276 42000
rect 134760 41948 134812 42000
rect 143684 41948 143736 42000
rect 58216 41880 58268 41932
rect 92716 41880 92768 41932
rect 100996 41880 101048 41932
rect 177632 41880 177684 41932
rect 185176 41880 185228 41932
rect 94004 41812 94056 41864
rect 100812 41812 100864 41864
rect 177724 41812 177776 41864
rect 184992 41812 185044 41864
rect 58308 41744 58360 41796
rect 139636 41744 139688 41796
rect 142764 41744 142816 41796
rect 134760 40792 134812 40844
rect 139636 40792 139688 40844
rect 51224 40656 51276 40708
rect 55732 40656 55784 40708
rect 134576 40656 134628 40708
rect 134760 40656 134812 40708
rect 138072 40656 138124 40708
rect 51132 40588 51184 40640
rect 56560 40588 56612 40640
rect 134668 40588 134720 40640
rect 92716 40520 92768 40572
rect 100996 40520 101048 40572
rect 137980 40563 138032 40572
rect 137980 40529 137989 40563
rect 137989 40529 138023 40563
rect 138023 40529 138032 40563
rect 137980 40520 138032 40529
rect 142396 40520 142448 40572
rect 177264 40520 177316 40572
rect 185176 40520 185228 40572
rect 94004 40452 94056 40504
rect 100904 40452 100956 40504
rect 177724 40452 177776 40504
rect 185084 40452 185136 40504
rect 56560 40384 56612 40436
rect 58216 40384 58268 40436
rect 55732 40112 55784 40164
rect 58308 40112 58360 40164
rect 51132 39228 51184 39280
rect 13320 39160 13372 39212
rect 18104 39160 18156 39212
rect 51224 39160 51276 39212
rect 134576 39228 134628 39280
rect 134668 39160 134720 39212
rect 58216 39092 58268 39144
rect 92900 39092 92952 39144
rect 100996 39092 101048 39144
rect 58400 39024 58452 39076
rect 93912 39024 93964 39076
rect 101088 39024 101140 39076
rect 94004 38956 94056 39008
rect 100812 38956 100864 39008
rect 142396 39092 142448 39144
rect 177356 39092 177408 39144
rect 185176 39092 185228 39144
rect 139636 39024 139688 39076
rect 142488 39024 142540 39076
rect 177448 39024 177500 39076
rect 185268 39024 185320 39076
rect 142580 38956 142632 39008
rect 177724 38956 177776 39008
rect 184992 38956 185044 39008
rect 51224 38412 51276 38464
rect 58308 38412 58360 38464
rect 183704 38140 183756 38192
rect 185268 38140 185320 38192
rect 134668 37936 134720 37988
rect 142580 37936 142632 37988
rect 51132 37868 51184 37920
rect 58400 37868 58452 37920
rect 98236 37868 98288 37920
rect 101088 37868 101140 37920
rect 134300 37868 134352 37920
rect 142488 37868 142540 37920
rect 51224 37800 51276 37852
rect 58216 37800 58268 37852
rect 90600 37843 90652 37852
rect 90600 37809 90609 37843
rect 90609 37809 90643 37843
rect 90643 37809 90652 37843
rect 90600 37800 90652 37809
rect 98328 37800 98380 37852
rect 100996 37800 101048 37852
rect 134116 37800 134168 37852
rect 142396 37800 142448 37852
rect 183244 37800 183296 37852
rect 185176 37800 185228 37852
rect 94004 37596 94056 37648
rect 98236 37596 98288 37648
rect 177448 37324 177500 37376
rect 183704 37324 183756 37376
rect 94004 37052 94056 37104
rect 98328 37052 98380 37104
rect 177724 36848 177776 36900
rect 183244 36848 183296 36900
rect 134392 36576 134444 36628
rect 140924 36576 140976 36628
rect 51224 36508 51276 36560
rect 58308 36508 58360 36560
rect 51132 36440 51184 36492
rect 58216 36440 58268 36492
rect 134668 36440 134720 36492
rect 142396 36440 142448 36492
rect 92900 36372 92952 36424
rect 100996 36372 101048 36424
rect 177356 36372 177408 36424
rect 185176 36372 185228 36424
rect 94004 36304 94056 36356
rect 100812 36304 100864 36356
rect 177724 36304 177776 36356
rect 184992 36304 185044 36356
rect 134668 35624 134720 35676
rect 140188 35624 140240 35676
rect 50028 35216 50080 35268
rect 55456 35216 55508 35268
rect 51224 35080 51276 35132
rect 134116 35080 134168 35132
rect 142488 35080 142540 35132
rect 58308 35012 58360 35064
rect 93452 35012 93504 35064
rect 100996 35012 101048 35064
rect 140924 35012 140976 35064
rect 142580 35012 142632 35064
rect 177632 35012 177684 35064
rect 185452 35012 185504 35064
rect 55456 34944 55508 34996
rect 58216 34944 58268 34996
rect 94004 34944 94056 34996
rect 100904 34944 100956 34996
rect 177724 34944 177776 34996
rect 185084 34944 185136 34996
rect 140188 34876 140240 34928
rect 142396 34876 142448 34928
rect 51224 33992 51276 34044
rect 56744 33992 56796 34044
rect 134668 33992 134720 34044
rect 140188 33992 140240 34044
rect 50212 33720 50264 33772
rect 51224 33652 51276 33704
rect 56008 33652 56060 33704
rect 134668 33720 134720 33772
rect 140924 33720 140976 33772
rect 134576 33652 134628 33704
rect 58216 33584 58268 33636
rect 93820 33584 93872 33636
rect 100996 33584 101048 33636
rect 142396 33584 142448 33636
rect 177816 33584 177868 33636
rect 185176 33584 185228 33636
rect 94004 33516 94056 33568
rect 101088 33516 101140 33568
rect 177724 33516 177776 33568
rect 185268 33516 185320 33568
rect 56744 33448 56796 33500
rect 58216 33448 58268 33500
rect 93912 33448 93964 33500
rect 100720 33448 100772 33500
rect 177632 33448 177684 33500
rect 184900 33448 184952 33500
rect 140188 33176 140240 33228
rect 142396 33176 142448 33228
rect 56008 32972 56060 33024
rect 58216 32972 58268 33024
rect 51224 32360 51276 32412
rect 56744 32360 56796 32412
rect 134392 32360 134444 32412
rect 139728 32360 139780 32412
rect 50028 32292 50080 32344
rect 56652 32292 56704 32344
rect 134300 32292 134352 32344
rect 93912 32224 93964 32276
rect 100996 32224 101048 32276
rect 142396 32224 142448 32276
rect 177724 32224 177776 32276
rect 185176 32224 185228 32276
rect 56652 32156 56704 32208
rect 58216 32156 58268 32208
rect 94004 32156 94056 32208
rect 100812 32156 100864 32208
rect 140924 32156 140976 32208
rect 142488 32156 142540 32208
rect 176988 32156 177040 32208
rect 184992 32156 185044 32208
rect 56744 31816 56796 31868
rect 58308 31816 58360 31868
rect 134668 31272 134720 31324
rect 139636 31272 139688 31324
rect 51132 31000 51184 31052
rect 51224 30932 51276 30984
rect 134668 30932 134720 30984
rect 143592 30932 143644 30984
rect 58216 30864 58268 30916
rect 92716 30864 92768 30916
rect 100996 30864 101048 30916
rect 134392 30864 134444 30916
rect 134852 30864 134904 30916
rect 177172 30864 177224 30916
rect 185176 30864 185228 30916
rect 94004 30796 94056 30848
rect 100904 30796 100956 30848
rect 177448 30796 177500 30848
rect 185084 30796 185136 30848
rect 58308 30728 58360 30780
rect 139728 30728 139780 30780
rect 142396 30728 142448 30780
rect 139636 30524 139688 30576
rect 142396 30524 142448 30576
rect 51132 29572 51184 29624
rect 51224 29504 51276 29556
rect 56652 29504 56704 29556
rect 134760 29572 134812 29624
rect 134208 29504 134260 29556
rect 58216 29436 58268 29488
rect 93912 29436 93964 29488
rect 101088 29436 101140 29488
rect 92716 29368 92768 29420
rect 100996 29368 101048 29420
rect 142396 29436 142448 29488
rect 177816 29436 177868 29488
rect 185268 29436 185320 29488
rect 142488 29368 142540 29420
rect 177632 29368 177684 29420
rect 185176 29368 185228 29420
rect 94004 29300 94056 29352
rect 100812 29300 100864 29352
rect 177724 29300 177776 29352
rect 184992 29300 185044 29352
rect 56652 29232 56704 29284
rect 58216 29232 58268 29284
rect 51132 28756 51184 28808
rect 58216 28756 58268 28808
rect 51224 28552 51276 28604
rect 56744 28552 56796 28604
rect 134760 28416 134812 28468
rect 140280 28416 140332 28468
rect 51224 28280 51276 28332
rect 56008 28280 56060 28332
rect 134760 28212 134812 28264
rect 140924 28212 140976 28264
rect 93912 28144 93964 28196
rect 100996 28144 101048 28196
rect 134576 28144 134628 28196
rect 56744 28076 56796 28128
rect 58216 28076 58268 28128
rect 90692 28119 90744 28128
rect 90692 28085 90701 28119
rect 90701 28085 90735 28119
rect 90735 28085 90744 28119
rect 90692 28076 90744 28085
rect 94004 28076 94056 28128
rect 101180 28076 101232 28128
rect 177448 28144 177500 28196
rect 185176 28144 185228 28196
rect 142396 28076 142448 28128
rect 177724 28076 177776 28128
rect 185360 28076 185412 28128
rect 92716 28008 92768 28060
rect 101088 28008 101140 28060
rect 177264 28008 177316 28060
rect 185268 28008 185320 28060
rect 140280 27736 140332 27788
rect 142396 27736 142448 27788
rect 56008 27668 56060 27720
rect 58308 27668 58360 27720
rect 51224 26852 51276 26904
rect 58308 26852 58360 26904
rect 134760 26852 134812 26904
rect 142580 26852 142632 26904
rect 51132 26784 51184 26836
rect 58216 26784 58268 26836
rect 98236 26784 98288 26836
rect 100996 26784 101048 26836
rect 134576 26784 134628 26836
rect 142396 26784 142448 26836
rect 140924 26716 140976 26768
rect 142488 26716 142540 26768
rect 177724 26716 177776 26768
rect 185176 26784 185228 26836
rect 94004 26308 94056 26360
rect 98236 26308 98288 26360
rect 51132 25560 51184 25612
rect 59320 25560 59372 25612
rect 51224 25492 51276 25544
rect 59412 25492 59464 25544
rect 134760 25492 134812 25544
rect 142488 25492 142540 25544
rect 50488 25424 50540 25476
rect 59504 25424 59556 25476
rect 134576 25424 134628 25476
rect 142396 25424 142448 25476
rect 93820 25356 93872 25408
rect 100996 25356 101048 25408
rect 177356 25356 177408 25408
rect 185452 25356 185504 25408
rect 93912 25288 93964 25340
rect 101088 25288 101140 25340
rect 177724 25288 177776 25340
rect 185360 25288 185412 25340
rect 94004 25220 94056 25272
rect 101180 25220 101232 25272
rect 177632 25220 177684 25272
rect 185544 25220 185596 25272
rect 51132 24064 51184 24116
rect 51224 23996 51276 24048
rect 134576 24064 134628 24116
rect 134760 23996 134812 24048
rect 58216 23928 58268 23980
rect 92900 23928 92952 23980
rect 100996 23928 101048 23980
rect 58308 23860 58360 23912
rect 94004 23860 94056 23912
rect 101088 23860 101140 23912
rect 142396 23928 142448 23980
rect 177540 23928 177592 23980
rect 185176 23928 185228 23980
rect 142488 23860 142540 23912
rect 177724 23860 177776 23912
rect 185268 23860 185320 23912
rect 134760 22976 134812 23028
rect 140740 22976 140792 23028
rect 51224 22704 51276 22756
rect 55916 22704 55968 22756
rect 50212 22636 50264 22688
rect 58216 22568 58268 22620
rect 94004 22568 94056 22620
rect 100996 22704 101048 22756
rect 134760 22704 134812 22756
rect 139728 22704 139780 22756
rect 93912 22500 93964 22552
rect 101088 22636 101140 22688
rect 134576 22636 134628 22688
rect 100996 22568 101048 22620
rect 134392 22568 134444 22620
rect 134760 22568 134812 22620
rect 142396 22568 142448 22620
rect 177632 22568 177684 22620
rect 185268 22772 185320 22824
rect 96120 22296 96172 22348
rect 101088 22500 101140 22552
rect 140740 22500 140792 22552
rect 142488 22500 142540 22552
rect 177724 22500 177776 22552
rect 185176 22636 185228 22688
rect 174412 22432 174464 22484
rect 185176 22432 185228 22484
rect 55916 22160 55968 22212
rect 58308 22160 58360 22212
rect 51224 21276 51276 21328
rect 58216 21208 58268 21260
rect 94004 21208 94056 21260
rect 101180 21208 101232 21260
rect 137980 21208 138032 21260
rect 138164 21208 138216 21260
rect 139728 21208 139780 21260
rect 143684 21208 143736 21260
rect 177724 21208 177776 21260
rect 185268 21208 185320 21260
rect 93360 19780 93412 19832
rect 101824 19780 101876 19832
rect 176160 19780 176212 19832
rect 185268 19780 185320 19832
rect 94740 19712 94792 19764
rect 101548 19712 101600 19764
rect 177816 19712 177868 19764
rect 185176 19712 185228 19764
rect 18104 18420 18156 18472
rect 68244 18420 68296 18472
rect 80664 18420 80716 18472
rect 106700 18420 106752 18472
rect 112220 18420 112272 18472
rect 152240 18420 152292 18472
rect 153436 18420 153488 18472
rect 194928 18420 194980 18472
rect 212500 18420 212552 18472
rect 69900 18352 69952 18404
rect 138164 18352 138216 18404
rect 60792 18284 60844 18336
rect 54812 18216 54864 18268
rect 76248 18284 76300 18336
rect 78916 18284 78968 18336
rect 165948 18284 166000 18336
rect 166776 18284 166828 18336
rect 171376 18284 171428 18336
rect 171928 18284 171980 18336
rect 79652 18216 79704 18268
rect 42852 18148 42904 18200
rect 70636 18148 70688 18200
rect 153436 18216 153488 18268
rect 164292 18216 164344 18268
rect 168524 18216 168576 18268
rect 138164 18148 138216 18200
rect 48832 18080 48884 18132
rect 81676 18080 81728 18132
rect 36780 18012 36832 18064
rect 71372 18012 71424 18064
rect 30800 17944 30852 17996
rect 72384 17944 72436 17996
rect 132828 17944 132880 17996
rect 157576 17944 157628 17996
rect 167236 17944 167288 17996
rect 167788 17944 167840 17996
rect 18840 17876 18892 17928
rect 74776 17876 74828 17928
rect 138808 17876 138860 17928
rect 156380 17876 156432 17928
rect 24820 17808 24872 17860
rect 73396 17808 73448 17860
rect 126848 17808 126900 17860
rect 158496 17808 158548 17860
rect 12860 17740 12912 17792
rect 75512 17740 75564 17792
rect 86460 17740 86512 17792
rect 96856 17740 96908 17792
rect 120868 17740 120920 17792
rect 159508 17740 159560 17792
rect 77168 17536 77220 17588
rect 78824 17536 78876 17588
rect 162912 17536 162964 17588
rect 167144 17536 167196 17588
rect 169996 17536 170048 17588
rect 170916 17536 170968 17588
rect 76156 17468 76208 17520
rect 77536 17468 77588 17520
rect 162820 17400 162872 17452
rect 164660 17400 164712 17452
rect 87564 17196 87616 17248
rect 88944 17196 88996 17248
rect 84804 17128 84856 17180
rect 87932 17128 87984 17180
rect 150860 17128 150912 17180
rect 154356 17128 154408 17180
rect 67784 17060 67836 17112
rect 117832 17060 117884 17112
rect 151872 17060 151924 17112
rect 208912 17060 208964 17112
rect 167144 12776 167196 12828
rect 174872 12776 174924 12828
rect 161808 12708 161860 12760
rect 180852 12708 180904 12760
rect 171376 12640 171428 12692
rect 192812 12640 192864 12692
rect 160336 12572 160388 12624
rect 186832 12572 186884 12624
rect 85448 12504 85500 12556
rect 88944 12368 88996 12420
rect 90784 12368 90836 12420
rect 169996 12504 170048 12556
rect 198792 12504 198844 12556
rect 170088 12436 170140 12488
rect 204864 12436 204916 12488
rect 102836 12368 102888 12420
rect 168616 12368 168668 12420
rect 210844 12368 210896 12420
rect 84344 12300 84396 12352
rect 108816 12300 108868 12352
rect 167236 12300 167288 12352
rect 216824 12300 216876 12352
rect 66864 12232 66916 12284
rect 76248 12232 76300 12284
rect 83424 12232 83476 12284
rect 114796 12232 114848 12284
rect 144788 12232 144840 12284
rect 155368 12232 155420 12284
rect 156840 12232 156892 12284
rect 165856 12232 165908 12284
rect 166132 12232 166184 12284
rect 222804 12232 222856 12284
rect 72844 12096 72896 12148
rect 76156 12096 76208 12148
<< metal2 >>
rect 27854 244344 27910 244824
rect 63826 244344 63882 244824
rect 99798 244344 99854 244824
rect 135862 244344 135918 244824
rect 171834 244344 171890 244824
rect 207806 244344 207862 244824
rect 27868 241178 27896 244344
rect 27856 241172 27908 241178
rect 27856 241114 27908 241120
rect 29144 241172 29196 241178
rect 29144 241114 29196 241120
rect 12768 236684 12820 236690
rect 12768 236626 12820 236632
rect 12780 232921 12808 236626
rect 23440 236616 23492 236622
rect 23440 236558 23492 236564
rect 23452 234788 23480 236558
rect 29156 235942 29184 241114
rect 62540 236752 62592 236758
rect 62540 236694 62592 236700
rect 30432 236684 30484 236690
rect 30432 236626 30484 236632
rect 29144 235936 29196 235942
rect 29144 235878 29196 235884
rect 30444 234788 30472 236626
rect 47544 235256 47596 235262
rect 47544 235198 47596 235204
rect 37424 235188 37476 235194
rect 37424 235130 37476 235136
rect 37436 234788 37464 235130
rect 12766 232912 12822 232921
rect 12766 232847 12822 232856
rect 18102 220944 18158 220953
rect 18102 220879 18158 220888
rect 13318 209384 13374 209393
rect 13318 209319 13374 209328
rect 13332 184058 13360 209319
rect 18116 190994 18144 220879
rect 47556 207194 47584 235198
rect 50670 234544 50726 234553
rect 50670 234479 50726 234488
rect 49934 234000 49990 234009
rect 49934 233935 49990 233944
rect 49948 233834 49976 233935
rect 49936 233828 49988 233834
rect 49936 233770 49988 233776
rect 50578 233456 50634 233465
rect 50578 233391 50634 233400
rect 50592 232474 50620 233391
rect 50580 232468 50632 232474
rect 50580 232410 50632 232416
rect 50684 228274 50712 234479
rect 58124 233828 58176 233834
rect 58124 233770 58176 233776
rect 58136 233057 58164 233770
rect 58122 233048 58178 233057
rect 58122 232983 58178 232992
rect 51222 232912 51278 232921
rect 51222 232847 51278 232856
rect 51236 232542 51264 232847
rect 62552 232762 62580 236694
rect 63840 235874 63868 244344
rect 99812 244306 99840 244344
rect 99616 244300 99668 244306
rect 99616 244242 99668 244248
rect 99800 244300 99852 244306
rect 99800 244242 99852 244248
rect 89864 241376 89916 241382
rect 89864 241318 89916 241324
rect 72844 236616 72896 236622
rect 72844 236558 72896 236564
rect 63828 235868 63880 235874
rect 63828 235810 63880 235816
rect 65576 235256 65628 235262
rect 65576 235198 65628 235204
rect 65588 232762 65616 235198
rect 72856 232762 72884 236558
rect 82228 235936 82280 235942
rect 82228 235878 82280 235884
rect 86184 235936 86236 235942
rect 86184 235878 86236 235884
rect 79558 235224 79614 235233
rect 75512 235188 75564 235194
rect 79558 235159 79614 235168
rect 75512 235130 75564 235136
rect 62552 232734 62612 232762
rect 65588 232734 65924 232762
rect 72548 232734 72884 232762
rect 75524 232762 75552 235130
rect 79572 232762 79600 235159
rect 75524 232734 75860 232762
rect 79264 232734 79600 232762
rect 82240 232762 82268 235878
rect 86196 232762 86224 235878
rect 89876 232898 89904 241318
rect 99628 235942 99656 244242
rect 135876 240770 135904 244344
rect 171848 241382 171876 244344
rect 207820 241382 207848 244344
rect 171836 241376 171888 241382
rect 171836 241318 171888 241324
rect 174044 241376 174096 241382
rect 174044 241318 174096 241324
rect 207808 241376 207860 241382
rect 207808 241318 207860 241324
rect 135864 240764 135916 240770
rect 135864 240706 135916 240712
rect 136784 240764 136836 240770
rect 136784 240706 136836 240712
rect 107436 236684 107488 236690
rect 107436 236626 107488 236632
rect 99616 235936 99668 235942
rect 99616 235878 99668 235884
rect 107448 234788 107476 236626
rect 121420 236616 121472 236622
rect 121420 236558 121472 236564
rect 114428 235324 114480 235330
rect 114428 235266 114480 235272
rect 114440 234788 114468 235266
rect 121432 234788 121460 236558
rect 136796 235942 136824 240706
rect 146536 236684 146588 236690
rect 146536 236626 146588 236632
rect 136784 235936 136836 235942
rect 136784 235878 136836 235884
rect 146548 235194 146576 236626
rect 169536 235936 169588 235942
rect 169536 235878 169588 235884
rect 166224 235868 166276 235874
rect 166224 235810 166276 235816
rect 159508 235324 159560 235330
rect 159508 235266 159560 235272
rect 156840 235256 156892 235262
rect 156840 235198 156892 235204
rect 146536 235188 146588 235194
rect 146536 235130 146588 235136
rect 134758 234544 134814 234553
rect 134758 234479 134814 234488
rect 101638 234136 101694 234145
rect 101638 234071 101694 234080
rect 100994 233184 101050 233193
rect 100994 233119 101050 233128
rect 101008 233086 101036 233119
rect 92716 233080 92768 233086
rect 92716 233022 92768 233028
rect 100996 233080 101048 233086
rect 100996 233022 101048 233028
rect 89508 232870 89904 232898
rect 89508 232762 89536 232870
rect 82240 232734 82576 232762
rect 85888 232734 86224 232762
rect 89200 232734 89536 232762
rect 51224 232536 51276 232542
rect 51224 232478 51276 232484
rect 58032 232536 58084 232542
rect 92728 232513 92756 233022
rect 100994 232640 101050 232649
rect 100994 232575 101050 232584
rect 58032 232478 58084 232484
rect 92714 232504 92770 232513
rect 51130 232232 51186 232241
rect 51130 232167 51186 232176
rect 51144 231250 51172 232167
rect 51222 231688 51278 231697
rect 51222 231623 51278 231632
rect 51236 231386 51264 231623
rect 51224 231380 51276 231386
rect 51224 231322 51276 231328
rect 56744 231380 56796 231386
rect 56744 231322 56796 231328
rect 51132 231244 51184 231250
rect 51132 231186 51184 231192
rect 51222 231144 51278 231153
rect 51222 231079 51224 231088
rect 51276 231079 51278 231088
rect 52696 231108 52748 231114
rect 51224 231050 51276 231056
rect 52696 231050 52748 231056
rect 51130 230600 51186 230609
rect 51130 230535 51186 230544
rect 51144 229754 51172 230535
rect 51222 230056 51278 230065
rect 51222 229991 51278 230000
rect 51236 229890 51264 229991
rect 51224 229884 51276 229890
rect 51224 229826 51276 229832
rect 51132 229748 51184 229754
rect 51132 229690 51184 229696
rect 52708 229618 52736 231050
rect 56756 230774 56784 231322
rect 58044 231289 58072 232478
rect 58124 232468 58176 232474
rect 101008 232474 101036 232575
rect 92714 232439 92770 232448
rect 100996 232468 101048 232474
rect 58124 232410 58176 232416
rect 100996 232410 101048 232416
rect 58136 231969 58164 232410
rect 94004 232400 94056 232406
rect 94004 232342 94056 232348
rect 94016 231969 94044 232342
rect 100994 232096 101050 232105
rect 100994 232031 101050 232040
rect 58122 231960 58178 231969
rect 58122 231895 58178 231904
rect 94002 231960 94058 231969
rect 94002 231895 94058 231904
rect 101008 231726 101036 232031
rect 92716 231720 92768 231726
rect 92716 231662 92768 231668
rect 100996 231720 101048 231726
rect 100996 231662 101048 231668
rect 92728 231289 92756 231662
rect 100994 231552 101050 231561
rect 100994 231487 101050 231496
rect 58030 231280 58086 231289
rect 58030 231215 58086 231224
rect 92714 231280 92770 231289
rect 92714 231215 92770 231224
rect 101008 231182 101036 231487
rect 95384 231176 95436 231182
rect 95384 231118 95436 231124
rect 100996 231176 101048 231182
rect 100996 231118 101048 231124
rect 101086 231144 101142 231153
rect 94096 231040 94148 231046
rect 94096 230982 94148 230988
rect 58216 230972 58268 230978
rect 58216 230914 58268 230920
rect 56744 230768 56796 230774
rect 58228 230745 58256 230914
rect 92716 230904 92768 230910
rect 92716 230846 92768 230852
rect 58308 230768 58360 230774
rect 56744 230710 56796 230716
rect 58214 230736 58270 230745
rect 92728 230745 92756 230846
rect 58308 230710 58360 230716
rect 92714 230736 92770 230745
rect 58214 230671 58270 230680
rect 58320 230201 58348 230710
rect 92714 230671 92770 230680
rect 94108 230201 94136 230982
rect 95396 230910 95424 231118
rect 101086 231079 101142 231088
rect 101100 231046 101128 231079
rect 101088 231040 101140 231046
rect 101088 230982 101140 230988
rect 95384 230904 95436 230910
rect 95384 230846 95436 230852
rect 58306 230192 58362 230201
rect 58306 230127 58362 230136
rect 94094 230192 94150 230201
rect 94094 230127 94150 230136
rect 101086 230192 101142 230201
rect 101086 230127 101142 230136
rect 56468 229884 56520 229890
rect 56468 229826 56520 229832
rect 56192 229748 56244 229754
rect 56192 229690 56244 229696
rect 52696 229612 52748 229618
rect 52696 229554 52748 229560
rect 51130 229376 51186 229385
rect 56204 229346 56232 229690
rect 51130 229311 51186 229320
rect 56192 229340 56244 229346
rect 50762 228832 50818 228841
rect 50762 228767 50818 228776
rect 50776 228530 50804 228767
rect 50764 228524 50816 228530
rect 50764 228466 50816 228472
rect 51144 228394 51172 229311
rect 56192 229282 56244 229288
rect 56480 229074 56508 229826
rect 100994 229784 101050 229793
rect 100994 229719 101050 229728
rect 58216 229612 58268 229618
rect 58216 229554 58268 229560
rect 92716 229612 92768 229618
rect 92716 229554 92768 229560
rect 58228 229521 58256 229554
rect 92728 229521 92756 229554
rect 101008 229550 101036 229719
rect 101100 229618 101128 230127
rect 101088 229612 101140 229618
rect 101088 229554 101140 229560
rect 93176 229544 93228 229550
rect 58214 229512 58270 229521
rect 58214 229447 58270 229456
rect 92714 229512 92770 229521
rect 93176 229486 93228 229492
rect 100996 229544 101048 229550
rect 100996 229486 101048 229492
rect 92714 229447 92770 229456
rect 58216 229340 58268 229346
rect 58216 229282 58268 229288
rect 56468 229068 56520 229074
rect 56468 229010 56520 229016
rect 58228 228977 58256 229282
rect 58308 229068 58360 229074
rect 58308 229010 58360 229016
rect 58214 228968 58270 228977
rect 58214 228903 58270 228912
rect 55456 228524 55508 228530
rect 55456 228466 55508 228472
rect 51132 228388 51184 228394
rect 51132 228330 51184 228336
rect 51224 228320 51276 228326
rect 50592 228246 50712 228274
rect 51222 228288 51224 228297
rect 52696 228320 52748 228326
rect 51276 228288 51278 228297
rect 50486 225976 50542 225985
rect 50486 225911 50542 225920
rect 50500 225606 50528 225911
rect 50488 225600 50540 225606
rect 50488 225542 50540 225548
rect 50210 220264 50266 220273
rect 50210 220199 50266 220208
rect 50224 220030 50252 220199
rect 50212 220024 50264 220030
rect 50212 219966 50264 219972
rect 50210 219176 50266 219185
rect 50210 219111 50266 219120
rect 50224 218942 50252 219111
rect 50212 218936 50264 218942
rect 50212 218878 50264 218884
rect 50394 215096 50450 215105
rect 50394 215031 50450 215040
rect 50408 214930 50436 215031
rect 50396 214924 50448 214930
rect 50396 214866 50448 214872
rect 50210 213464 50266 213473
rect 50210 213399 50212 213408
rect 50264 213399 50266 213408
rect 50212 213370 50264 213376
rect 50592 207518 50620 228246
rect 52696 228262 52748 228268
rect 51222 228223 51278 228232
rect 50946 227744 51002 227753
rect 50946 227679 51002 227688
rect 50960 227306 50988 227679
rect 50948 227300 51000 227306
rect 50948 227242 51000 227248
rect 51222 227200 51278 227209
rect 51278 227158 51356 227186
rect 51222 227135 51278 227144
rect 50762 226520 50818 226529
rect 50762 226455 50818 226464
rect 50776 225538 50804 226455
rect 50764 225532 50816 225538
rect 50764 225474 50816 225480
rect 51328 225470 51356 227158
rect 52708 226830 52736 228262
rect 55468 227918 55496 228466
rect 58320 228297 58348 229010
rect 93188 228977 93216 229486
rect 100994 229240 101050 229249
rect 100994 229175 101050 229184
rect 93174 228968 93230 228977
rect 92716 228932 92768 228938
rect 101008 228938 101036 229175
rect 93174 228903 93230 228912
rect 100996 228932 101048 228938
rect 92716 228874 92768 228880
rect 100996 228874 101048 228880
rect 92728 228297 92756 228874
rect 101086 228696 101142 228705
rect 101086 228631 101142 228640
rect 58306 228288 58362 228297
rect 58216 228252 58268 228258
rect 58306 228223 58362 228232
rect 92714 228288 92770 228297
rect 100994 228288 101050 228297
rect 92714 228223 92770 228232
rect 93176 228252 93228 228258
rect 58216 228194 58268 228200
rect 101100 228258 101128 228631
rect 100994 228223 101050 228232
rect 101088 228252 101140 228258
rect 93176 228194 93228 228200
rect 55456 227912 55508 227918
rect 55456 227854 55508 227860
rect 58228 227753 58256 228194
rect 92716 228184 92768 228190
rect 92716 228126 92768 228132
rect 58308 227912 58360 227918
rect 58308 227854 58360 227860
rect 58214 227744 58270 227753
rect 58214 227679 58270 227688
rect 56744 227300 56796 227306
rect 56744 227242 56796 227248
rect 52696 226824 52748 226830
rect 52696 226766 52748 226772
rect 56756 226694 56784 227242
rect 58320 227209 58348 227854
rect 92728 227209 92756 228126
rect 93188 227753 93216 228194
rect 101008 228190 101036 228223
rect 101088 228194 101140 228200
rect 100996 228184 101048 228190
rect 100996 228126 101048 228132
rect 93174 227744 93230 227753
rect 93174 227679 93230 227688
rect 101086 227472 101142 227481
rect 101086 227407 101142 227416
rect 58306 227200 58362 227209
rect 58306 227135 58362 227144
rect 92714 227200 92770 227209
rect 92714 227135 92770 227144
rect 100994 227064 101050 227073
rect 100994 226999 101050 227008
rect 101008 226830 101036 226999
rect 58216 226824 58268 226830
rect 58216 226766 58268 226772
rect 93636 226824 93688 226830
rect 93636 226766 93688 226772
rect 100996 226824 101048 226830
rect 100996 226766 101048 226772
rect 56744 226688 56796 226694
rect 56744 226630 56796 226636
rect 58228 226529 58256 226766
rect 92716 226756 92768 226762
rect 92716 226698 92768 226704
rect 58308 226688 58360 226694
rect 58308 226630 58360 226636
rect 58214 226520 58270 226529
rect 58214 226455 58270 226464
rect 58320 225985 58348 226630
rect 92728 226529 92756 226698
rect 92714 226520 92770 226529
rect 92714 226455 92770 226464
rect 93648 225985 93676 226766
rect 101100 226762 101128 227407
rect 101088 226756 101140 226762
rect 101088 226698 101140 226704
rect 101086 226384 101142 226393
rect 101086 226319 101142 226328
rect 58306 225976 58362 225985
rect 58306 225911 58362 225920
rect 93634 225976 93690 225985
rect 93634 225911 93690 225920
rect 58400 225600 58452 225606
rect 58400 225542 58452 225548
rect 100994 225568 101050 225577
rect 58308 225532 58360 225538
rect 58308 225474 58360 225480
rect 51316 225464 51368 225470
rect 51130 225432 51186 225441
rect 51316 225406 51368 225412
rect 58216 225464 58268 225470
rect 58216 225406 58268 225412
rect 51130 225367 51186 225376
rect 51038 224344 51094 224353
rect 51038 224279 51040 224288
rect 51092 224279 51094 224288
rect 51040 224250 51092 224256
rect 51144 224246 51172 225367
rect 58228 225305 58256 225406
rect 58214 225296 58270 225305
rect 58214 225231 58270 225240
rect 51222 224888 51278 224897
rect 51222 224823 51278 224832
rect 51132 224240 51184 224246
rect 51132 224182 51184 224188
rect 51236 224178 51264 224823
rect 58320 224761 58348 225474
rect 58306 224752 58362 224761
rect 58306 224687 58362 224696
rect 52696 224308 52748 224314
rect 52696 224250 52748 224256
rect 51224 224172 51276 224178
rect 51224 224114 51276 224120
rect 50946 223664 51002 223673
rect 50946 223599 51002 223608
rect 50960 223226 50988 223599
rect 50948 223220 51000 223226
rect 50948 223162 51000 223168
rect 51222 223120 51278 223129
rect 51222 223055 51224 223064
rect 51276 223055 51278 223064
rect 51224 223026 51276 223032
rect 52708 222750 52736 224250
rect 58412 224217 58440 225542
rect 100994 225503 101050 225512
rect 92808 225464 92860 225470
rect 92808 225406 92860 225412
rect 92716 225328 92768 225334
rect 92820 225305 92848 225406
rect 101008 225402 101036 225503
rect 101100 225470 101128 226319
rect 101178 225704 101234 225713
rect 101178 225639 101234 225648
rect 101088 225464 101140 225470
rect 101088 225406 101140 225412
rect 92900 225396 92952 225402
rect 92900 225338 92952 225344
rect 100996 225396 101048 225402
rect 100996 225338 101048 225344
rect 92716 225270 92768 225276
rect 92806 225296 92862 225305
rect 92728 224761 92756 225270
rect 92806 225231 92862 225240
rect 92714 224752 92770 224761
rect 92714 224687 92770 224696
rect 92912 224217 92940 225338
rect 101192 225334 101220 225639
rect 101180 225328 101232 225334
rect 101180 225270 101232 225276
rect 101086 224616 101142 224625
rect 101086 224551 101142 224560
rect 58398 224208 58454 224217
rect 58398 224143 58454 224152
rect 92898 224208 92954 224217
rect 92898 224143 92954 224152
rect 100994 224208 101050 224217
rect 100994 224143 101050 224152
rect 101008 224110 101036 224143
rect 58216 224104 58268 224110
rect 58216 224046 58268 224052
rect 93912 224104 93964 224110
rect 93912 224046 93964 224052
rect 100996 224104 101048 224110
rect 100996 224046 101048 224052
rect 58228 223537 58256 224046
rect 58308 224036 58360 224042
rect 58308 223978 58360 223984
rect 93728 224036 93780 224042
rect 93728 223978 93780 223984
rect 58214 223528 58270 223537
rect 58214 223463 58270 223472
rect 56284 223220 56336 223226
rect 56284 223162 56336 223168
rect 52788 223084 52840 223090
rect 52788 223026 52840 223032
rect 52696 222744 52748 222750
rect 52696 222686 52748 222692
rect 51130 222576 51186 222585
rect 51130 222511 51186 222520
rect 51144 221594 51172 222511
rect 51222 222032 51278 222041
rect 51222 221967 51278 221976
rect 51236 221730 51264 221967
rect 51224 221724 51276 221730
rect 51224 221666 51276 221672
rect 51132 221588 51184 221594
rect 51132 221530 51184 221536
rect 51222 221488 51278 221497
rect 51222 221423 51224 221432
rect 51276 221423 51278 221432
rect 52696 221452 52748 221458
rect 51224 221394 51276 221400
rect 52696 221394 52748 221400
rect 50946 220808 51002 220817
rect 50946 220743 51002 220752
rect 50960 220370 50988 220743
rect 50948 220364 51000 220370
rect 50948 220306 51000 220312
rect 52708 219962 52736 221394
rect 52800 221322 52828 223026
rect 56296 222478 56324 223162
rect 58320 222993 58348 223978
rect 93740 223537 93768 223978
rect 93726 223528 93782 223537
rect 93726 223463 93782 223472
rect 93924 222993 93952 224046
rect 101100 224042 101128 224551
rect 101088 224036 101140 224042
rect 101088 223978 101140 223984
rect 101454 223528 101510 223537
rect 101454 223463 101510 223472
rect 58306 222984 58362 222993
rect 58306 222919 58362 222928
rect 93910 222984 93966 222993
rect 93910 222919 93966 222928
rect 101270 222848 101326 222857
rect 101270 222783 101326 222792
rect 58216 222744 58268 222750
rect 58216 222686 58268 222692
rect 92716 222744 92768 222750
rect 92716 222686 92768 222692
rect 56284 222472 56336 222478
rect 56284 222414 56336 222420
rect 58228 222313 58256 222686
rect 58308 222472 58360 222478
rect 58308 222414 58360 222420
rect 58214 222304 58270 222313
rect 58214 222239 58270 222248
rect 58320 221769 58348 222414
rect 92728 222313 92756 222686
rect 92992 222676 93044 222682
rect 92992 222618 93044 222624
rect 92714 222304 92770 222313
rect 92714 222239 92770 222248
rect 93004 221769 93032 222618
rect 58306 221760 58362 221769
rect 56744 221724 56796 221730
rect 58306 221695 58362 221704
rect 92990 221760 93046 221769
rect 92990 221695 93046 221704
rect 56744 221666 56796 221672
rect 55916 221588 55968 221594
rect 55916 221530 55968 221536
rect 52788 221316 52840 221322
rect 52788 221258 52840 221264
rect 55928 221050 55956 221530
rect 55916 221044 55968 221050
rect 55916 220986 55968 220992
rect 56756 220914 56784 221666
rect 58216 221316 58268 221322
rect 58216 221258 58268 221264
rect 93176 221316 93228 221322
rect 93176 221258 93228 221264
rect 58228 221225 58256 221258
rect 58214 221216 58270 221225
rect 58214 221151 58270 221160
rect 92714 221216 92770 221225
rect 92714 221151 92716 221160
rect 92768 221151 92770 221160
rect 92716 221122 92768 221128
rect 58216 221044 58268 221050
rect 58216 220986 58268 220992
rect 56744 220908 56796 220914
rect 56744 220850 56796 220856
rect 58228 220545 58256 220986
rect 58308 220908 58360 220914
rect 58308 220850 58360 220856
rect 58214 220536 58270 220545
rect 58214 220471 58270 220480
rect 56468 220364 56520 220370
rect 56468 220306 56520 220312
rect 52788 220024 52840 220030
rect 52788 219966 52840 219972
rect 52696 219956 52748 219962
rect 52696 219898 52748 219904
rect 50854 219720 50910 219729
rect 50854 219655 50910 219664
rect 50868 218670 50896 219655
rect 51224 218732 51276 218738
rect 51224 218674 51276 218680
rect 52696 218732 52748 218738
rect 52696 218674 52748 218680
rect 50856 218664 50908 218670
rect 51236 218641 51264 218674
rect 50856 218606 50908 218612
rect 51222 218632 51278 218641
rect 51222 218567 51278 218576
rect 51222 217952 51278 217961
rect 51222 217887 51278 217896
rect 51236 217514 51264 217887
rect 51224 217508 51276 217514
rect 51224 217450 51276 217456
rect 51222 217408 51278 217417
rect 51222 217343 51224 217352
rect 51276 217343 51278 217352
rect 51224 217314 51276 217320
rect 52708 217174 52736 218674
rect 52800 218602 52828 219966
rect 56480 219554 56508 220306
rect 58320 220001 58348 220850
rect 93188 220001 93216 221258
rect 93728 221248 93780 221254
rect 93728 221190 93780 221196
rect 93740 220545 93768 221190
rect 101284 221186 101312 222783
rect 101468 222750 101496 223463
rect 101546 223120 101602 223129
rect 101546 223055 101602 223064
rect 101456 222744 101508 222750
rect 101456 222686 101508 222692
rect 101560 222682 101588 223055
rect 101548 222676 101600 222682
rect 101548 222618 101600 222624
rect 101546 221896 101602 221905
rect 101546 221831 101602 221840
rect 101560 221254 101588 221831
rect 101548 221248 101600 221254
rect 101548 221190 101600 221196
rect 101272 221180 101324 221186
rect 101272 221122 101324 221128
rect 93726 220536 93782 220545
rect 93726 220471 93782 220480
rect 58306 219992 58362 220001
rect 58216 219956 58268 219962
rect 93174 219992 93230 220001
rect 58306 219927 58362 219936
rect 92716 219956 92768 219962
rect 58216 219898 58268 219904
rect 93174 219927 93230 219936
rect 92716 219898 92768 219904
rect 56468 219548 56520 219554
rect 56468 219490 56520 219496
rect 58228 219321 58256 219898
rect 58308 219548 58360 219554
rect 58308 219490 58360 219496
rect 58214 219312 58270 219321
rect 58214 219247 58270 219256
rect 53064 218936 53116 218942
rect 53064 218878 53116 218884
rect 52788 218596 52840 218602
rect 52788 218538 52840 218544
rect 52880 217508 52932 217514
rect 52880 217450 52932 217456
rect 52788 217372 52840 217378
rect 52788 217314 52840 217320
rect 52696 217168 52748 217174
rect 52696 217110 52748 217116
rect 51130 216864 51186 216873
rect 51130 216799 51186 216808
rect 51144 215882 51172 216799
rect 51222 216320 51278 216329
rect 51278 216278 51356 216306
rect 51222 216255 51278 216264
rect 51132 215876 51184 215882
rect 51132 215818 51184 215824
rect 51222 215776 51278 215785
rect 51222 215711 51278 215720
rect 51132 214584 51184 214590
rect 51130 214552 51132 214561
rect 51184 214552 51186 214561
rect 51236 214522 51264 215711
rect 51130 214487 51186 214496
rect 51224 214516 51276 214522
rect 51224 214458 51276 214464
rect 51328 214454 51356 216278
rect 52800 215814 52828 217314
rect 52788 215808 52840 215814
rect 52788 215750 52840 215756
rect 52892 215746 52920 217450
rect 53076 217106 53104 218878
rect 58320 218777 58348 219490
rect 92728 218777 92756 219898
rect 92808 219888 92860 219894
rect 92808 219830 92860 219836
rect 92820 219321 92848 219830
rect 92806 219312 92862 219321
rect 92806 219247 92862 219256
rect 58306 218768 58362 218777
rect 58306 218703 58362 218712
rect 92714 218768 92770 218777
rect 92714 218703 92770 218712
rect 55456 218664 55508 218670
rect 55456 218606 55508 218612
rect 55468 218058 55496 218606
rect 58216 218596 58268 218602
rect 58216 218538 58268 218544
rect 92808 218596 92860 218602
rect 92808 218538 92860 218544
rect 58228 218233 58256 218538
rect 92820 218233 92848 218538
rect 93728 218528 93780 218534
rect 93728 218470 93780 218476
rect 58214 218224 58270 218233
rect 58214 218159 58270 218168
rect 92806 218224 92862 218233
rect 92806 218159 92862 218168
rect 55456 218052 55508 218058
rect 55456 217994 55508 218000
rect 58216 218052 58268 218058
rect 58216 217994 58268 218000
rect 58228 217553 58256 217994
rect 93740 217553 93768 218470
rect 58214 217544 58270 217553
rect 58214 217479 58270 217488
rect 93726 217544 93782 217553
rect 93726 217479 93782 217488
rect 97960 217304 98012 217310
rect 97960 217246 98012 217252
rect 58308 217168 58360 217174
rect 58308 217110 58360 217116
rect 92716 217168 92768 217174
rect 92716 217110 92768 217116
rect 53064 217100 53116 217106
rect 53064 217042 53116 217048
rect 58216 217100 58268 217106
rect 58216 217042 58268 217048
rect 58228 217009 58256 217042
rect 58214 217000 58270 217009
rect 58214 216935 58270 216944
rect 58320 216329 58348 217110
rect 92728 216329 92756 217110
rect 93912 217100 93964 217106
rect 93912 217042 93964 217048
rect 93924 217009 93952 217042
rect 93910 217000 93966 217009
rect 93910 216935 93966 216944
rect 58306 216320 58362 216329
rect 58306 216255 58362 216264
rect 92714 216320 92770 216329
rect 92714 216255 92770 216264
rect 56652 215876 56704 215882
rect 56652 215818 56704 215824
rect 52880 215740 52932 215746
rect 52880 215682 52932 215688
rect 56664 215202 56692 215818
rect 58308 215808 58360 215814
rect 58214 215776 58270 215785
rect 93544 215808 93596 215814
rect 58308 215750 58360 215756
rect 92714 215776 92770 215785
rect 58214 215711 58216 215720
rect 58268 215711 58270 215720
rect 58216 215682 58268 215688
rect 58320 215241 58348 215750
rect 93544 215750 93596 215756
rect 92714 215711 92716 215720
rect 92768 215711 92770 215720
rect 92716 215682 92768 215688
rect 92808 215672 92860 215678
rect 92808 215614 92860 215620
rect 92820 215241 92848 215614
rect 58306 215232 58362 215241
rect 56652 215196 56704 215202
rect 56652 215138 56704 215144
rect 58216 215196 58268 215202
rect 58306 215167 58362 215176
rect 92806 215232 92862 215241
rect 92806 215167 92862 215176
rect 58216 215138 58268 215144
rect 52788 214924 52840 214930
rect 52788 214866 52840 214872
rect 52696 214584 52748 214590
rect 52696 214526 52748 214532
rect 51316 214448 51368 214454
rect 51316 214390 51368 214396
rect 50946 214008 51002 214017
rect 50946 213943 51002 213952
rect 50960 213298 50988 213943
rect 50948 213292 51000 213298
rect 50948 213234 51000 213240
rect 52708 213094 52736 214526
rect 52696 213088 52748 213094
rect 52696 213030 52748 213036
rect 52800 213026 52828 214866
rect 58228 214561 58256 215138
rect 93556 214561 93584 215750
rect 97972 215746 98000 217246
rect 98052 217236 98104 217242
rect 98052 217178 98104 217184
rect 97960 215740 98012 215746
rect 97960 215682 98012 215688
rect 98064 215678 98092 217178
rect 98144 215876 98196 215882
rect 98144 215818 98196 215824
rect 98052 215672 98104 215678
rect 98052 215614 98104 215620
rect 58214 214552 58270 214561
rect 93542 214552 93598 214561
rect 58214 214487 58270 214496
rect 58308 214516 58360 214522
rect 93542 214487 93598 214496
rect 98052 214516 98104 214522
rect 58308 214458 58360 214464
rect 98052 214458 98104 214464
rect 58216 214448 58268 214454
rect 58216 214390 58268 214396
rect 58228 214017 58256 214390
rect 58214 214008 58270 214017
rect 58214 213943 58270 213952
rect 52880 213428 52932 213434
rect 52880 213370 52932 213376
rect 52788 213020 52840 213026
rect 52788 212962 52840 212968
rect 50762 212920 50818 212929
rect 50762 212855 50818 212864
rect 50776 211938 50804 212855
rect 51222 212240 51278 212249
rect 51222 212175 51278 212184
rect 51236 212074 51264 212175
rect 51224 212068 51276 212074
rect 51224 212010 51276 212016
rect 52696 212068 52748 212074
rect 52696 212010 52748 212016
rect 50764 211932 50816 211938
rect 50764 211874 50816 211880
rect 51130 211696 51186 211705
rect 51130 211631 51186 211640
rect 50670 211152 50726 211161
rect 50670 211087 50726 211096
rect 50580 207512 50632 207518
rect 50580 207454 50632 207460
rect 47478 207166 47584 207194
rect 20232 204118 20260 206908
rect 20220 204112 20272 204118
rect 20220 204054 20272 204060
rect 20876 203438 20904 206908
rect 21520 203710 21548 206908
rect 22164 204390 22192 206908
rect 22808 204662 22836 206908
rect 22796 204656 22848 204662
rect 22796 204598 22848 204604
rect 23452 204594 23480 206908
rect 23440 204588 23492 204594
rect 23440 204530 23492 204536
rect 24096 204458 24124 206908
rect 24084 204452 24136 204458
rect 24084 204394 24136 204400
rect 22152 204384 22204 204390
rect 22152 204326 22204 204332
rect 24740 204322 24768 206908
rect 24728 204316 24780 204322
rect 24728 204258 24780 204264
rect 21508 203704 21560 203710
rect 21508 203646 21560 203652
rect 25384 203438 25412 206908
rect 26042 206894 26424 206922
rect 20864 203432 20916 203438
rect 20864 203374 20916 203380
rect 24360 203432 24412 203438
rect 24360 203374 24412 203380
rect 25372 203432 25424 203438
rect 25372 203374 25424 203380
rect 26292 203432 26344 203438
rect 26292 203374 26344 203380
rect 24372 196366 24400 203374
rect 24360 196360 24412 196366
rect 24360 196302 24412 196308
rect 26108 196360 26160 196366
rect 26108 196302 26160 196308
rect 26120 193716 26148 196302
rect 26304 195686 26332 203374
rect 26396 195822 26424 206894
rect 26672 204526 26700 206908
rect 27330 206894 27712 206922
rect 26844 204656 26896 204662
rect 26844 204598 26896 204604
rect 26752 204588 26804 204594
rect 26752 204530 26804 204536
rect 26660 204520 26712 204526
rect 26660 204462 26712 204468
rect 26660 204384 26712 204390
rect 26660 204326 26712 204332
rect 26568 196360 26620 196366
rect 26568 196302 26620 196308
rect 26384 195816 26436 195822
rect 26384 195758 26436 195764
rect 26292 195680 26344 195686
rect 26292 195622 26344 195628
rect 26580 193730 26608 196302
rect 26502 193702 26608 193730
rect 26672 193730 26700 204326
rect 26764 196434 26792 204530
rect 26752 196428 26804 196434
rect 26752 196370 26804 196376
rect 26856 194138 26884 204598
rect 26936 203704 26988 203710
rect 26936 203646 26988 203652
rect 26948 196366 26976 203646
rect 27396 196428 27448 196434
rect 27396 196370 27448 196376
rect 26936 196360 26988 196366
rect 26936 196302 26988 196308
rect 26856 194110 26976 194138
rect 26948 193730 26976 194110
rect 27408 193730 27436 196370
rect 27684 196298 27712 206894
rect 27764 204520 27816 204526
rect 27764 204462 27816 204468
rect 27776 196366 27804 204462
rect 27960 203438 27988 206908
rect 28618 206894 29092 206922
rect 28040 204452 28092 204458
rect 28040 204394 28092 204400
rect 27948 203432 28000 203438
rect 27948 203374 28000 203380
rect 27764 196360 27816 196366
rect 27764 196302 27816 196308
rect 27672 196292 27724 196298
rect 27672 196234 27724 196240
rect 26672 193702 26870 193730
rect 26948 193702 27330 193730
rect 27408 193702 27698 193730
rect 28052 193716 28080 204394
rect 28132 204316 28184 204322
rect 28132 204258 28184 204264
rect 28144 193730 28172 204258
rect 29064 196162 29092 206894
rect 29248 203438 29276 206908
rect 29998 206894 30472 206922
rect 30642 206894 31024 206922
rect 29144 203432 29196 203438
rect 29144 203374 29196 203380
rect 29236 203432 29288 203438
rect 29236 203374 29288 203380
rect 30248 203432 30300 203438
rect 30248 203374 30300 203380
rect 29052 196156 29104 196162
rect 29052 196098 29104 196104
rect 28868 195680 28920 195686
rect 28868 195622 28920 195628
rect 28144 193702 28526 193730
rect 28880 193716 28908 195622
rect 29156 195346 29184 203374
rect 30260 199306 30288 203374
rect 30444 203114 30472 206894
rect 30444 203086 30564 203114
rect 30260 199278 30472 199306
rect 30444 196434 30472 199278
rect 30432 196428 30484 196434
rect 30432 196370 30484 196376
rect 30536 196366 30564 203086
rect 30996 202894 31024 206894
rect 31272 203438 31300 206908
rect 31732 206894 31930 206922
rect 32008 206894 32574 206922
rect 33218 206894 33324 206922
rect 31260 203432 31312 203438
rect 31260 203374 31312 203380
rect 30984 202888 31036 202894
rect 30984 202830 31036 202836
rect 31732 196434 31760 206894
rect 31812 203432 31864 203438
rect 31812 203374 31864 203380
rect 31260 196428 31312 196434
rect 31260 196370 31312 196376
rect 31720 196428 31772 196434
rect 31720 196370 31772 196376
rect 29696 196360 29748 196366
rect 29696 196302 29748 196308
rect 30524 196360 30576 196366
rect 30524 196302 30576 196308
rect 29236 195816 29288 195822
rect 29236 195758 29288 195764
rect 29144 195340 29196 195346
rect 29144 195282 29196 195288
rect 29248 193716 29276 195758
rect 29708 193716 29736 196302
rect 30064 196292 30116 196298
rect 30064 196234 30116 196240
rect 30076 193716 30104 196234
rect 30892 196156 30944 196162
rect 30892 196098 30944 196104
rect 30432 195340 30484 195346
rect 30432 195282 30484 195288
rect 30444 193716 30472 195282
rect 30904 193716 30932 196098
rect 31272 193716 31300 196370
rect 31628 196360 31680 196366
rect 31628 196302 31680 196308
rect 31640 193716 31668 196302
rect 31824 195346 31852 203374
rect 31904 202888 31956 202894
rect 31904 202830 31956 202836
rect 31812 195340 31864 195346
rect 31812 195282 31864 195288
rect 31916 195226 31944 202830
rect 32008 196366 32036 206894
rect 32824 196428 32876 196434
rect 32824 196370 32876 196376
rect 31996 196360 32048 196366
rect 31996 196302 32048 196308
rect 32456 195340 32508 195346
rect 32456 195282 32508 195288
rect 31916 195198 32036 195226
rect 32008 193730 32036 195198
rect 32008 193702 32114 193730
rect 32468 193716 32496 195282
rect 32836 193716 32864 196370
rect 32916 196360 32968 196366
rect 32916 196302 32968 196308
rect 32928 193730 32956 196302
rect 33296 195226 33324 206894
rect 33480 206894 33862 206922
rect 34216 206894 34506 206922
rect 34860 206894 35150 206922
rect 35504 206894 35794 206922
rect 36148 206894 36438 206922
rect 33376 203092 33428 203098
rect 33376 203034 33428 203040
rect 33388 196366 33416 203034
rect 33376 196360 33428 196366
rect 33376 196302 33428 196308
rect 33480 195618 33508 206894
rect 34216 203098 34244 206894
rect 34204 203092 34256 203098
rect 34204 203034 34256 203040
rect 34756 203092 34808 203098
rect 34756 203034 34808 203040
rect 34768 196366 34796 203034
rect 34480 196360 34532 196366
rect 34480 196302 34532 196308
rect 34756 196360 34808 196366
rect 34756 196302 34808 196308
rect 33468 195612 33520 195618
rect 33468 195554 33520 195560
rect 34112 195612 34164 195618
rect 34112 195554 34164 195560
rect 33296 195198 33416 195226
rect 33388 193730 33416 195198
rect 32928 193702 33310 193730
rect 33388 193702 33678 193730
rect 34124 193716 34152 195554
rect 34492 193716 34520 196302
rect 34860 193716 34888 206894
rect 35504 203098 35532 206894
rect 36148 204474 36176 206894
rect 35964 204446 36176 204474
rect 35492 203092 35544 203098
rect 35492 203034 35544 203040
rect 35308 196360 35360 196366
rect 35308 196302 35360 196308
rect 35320 193716 35348 196302
rect 35964 193730 35992 204446
rect 37068 203710 37096 206908
rect 37528 206894 37726 206922
rect 36044 203704 36096 203710
rect 36044 203646 36096 203652
rect 37056 203704 37108 203710
rect 37056 203646 37108 203652
rect 35702 193702 35992 193730
rect 36056 193716 36084 203646
rect 37528 203522 37556 206894
rect 37332 203500 37384 203506
rect 37332 203442 37384 203448
rect 37436 203494 37556 203522
rect 37240 203432 37292 203438
rect 37240 203374 37292 203380
rect 37252 196366 37280 203374
rect 36872 196360 36924 196366
rect 36872 196302 36924 196308
rect 37240 196360 37292 196366
rect 37240 196302 37292 196308
rect 36504 195612 36556 195618
rect 36504 195554 36556 195560
rect 36516 193716 36544 195554
rect 36884 193716 36912 196302
rect 37344 193730 37372 203442
rect 37436 195618 37464 203494
rect 38356 203438 38384 206908
rect 39092 203506 39120 206908
rect 39368 206894 39750 206922
rect 39080 203500 39132 203506
rect 39080 203442 39132 203448
rect 38344 203432 38396 203438
rect 38344 203374 38396 203380
rect 39264 196428 39316 196434
rect 39264 196370 39316 196376
rect 37700 196360 37752 196366
rect 37700 196302 37752 196308
rect 37424 195612 37476 195618
rect 37424 195554 37476 195560
rect 37266 193702 37372 193730
rect 37712 193716 37740 196302
rect 38068 196088 38120 196094
rect 38068 196030 38120 196036
rect 38080 193716 38108 196030
rect 38896 196020 38948 196026
rect 38896 195962 38948 195968
rect 38436 195748 38488 195754
rect 38436 195690 38488 195696
rect 38448 193716 38476 195690
rect 38908 193716 38936 195962
rect 39276 193716 39304 196370
rect 39368 196366 39396 206894
rect 39540 203568 39592 203574
rect 39540 203510 39592 203516
rect 39356 196360 39408 196366
rect 39356 196302 39408 196308
rect 39552 195754 39580 203510
rect 40380 203438 40408 206908
rect 40920 203636 40972 203642
rect 40920 203578 40972 203584
rect 39632 203432 39684 203438
rect 39632 203374 39684 203380
rect 40368 203432 40420 203438
rect 40368 203374 40420 203380
rect 39644 196094 39672 203374
rect 40932 196366 40960 203578
rect 41024 203574 41052 206908
rect 41012 203568 41064 203574
rect 41012 203510 41064 203516
rect 41196 203568 41248 203574
rect 41196 203510 41248 203516
rect 41104 203500 41156 203506
rect 41104 203442 41156 203448
rect 41012 203432 41064 203438
rect 41012 203374 41064 203380
rect 40092 196360 40144 196366
rect 40092 196302 40144 196308
rect 40920 196360 40972 196366
rect 40920 196302 40972 196308
rect 39632 196088 39684 196094
rect 39632 196030 39684 196036
rect 39632 195952 39684 195958
rect 39632 195894 39684 195900
rect 39540 195748 39592 195754
rect 39540 195690 39592 195696
rect 39644 193716 39672 195894
rect 40104 193716 40132 196302
rect 41024 196026 41052 203374
rect 41116 196434 41144 203442
rect 41104 196428 41156 196434
rect 41104 196370 41156 196376
rect 41012 196020 41064 196026
rect 41012 195962 41064 195968
rect 41208 195958 41236 203510
rect 41668 203438 41696 206908
rect 41748 204112 41800 204118
rect 41748 204054 41800 204060
rect 41656 203432 41708 203438
rect 41656 203374 41708 203380
rect 41656 196360 41708 196366
rect 41656 196302 41708 196308
rect 41196 195952 41248 195958
rect 41196 195894 41248 195900
rect 41288 195748 41340 195754
rect 41288 195690 41340 195696
rect 40460 195680 40512 195686
rect 40460 195622 40512 195628
rect 40472 193716 40500 195622
rect 40828 195612 40880 195618
rect 40828 195554 40880 195560
rect 40840 193716 40868 195554
rect 41300 193716 41328 195690
rect 41668 193716 41696 196302
rect 18104 190988 18156 190994
rect 18104 190930 18156 190936
rect 22336 190988 22388 190994
rect 22336 190930 22388 190936
rect 22348 190489 22376 190930
rect 22334 190480 22390 190489
rect 22334 190415 22390 190424
rect 41760 189242 41788 204054
rect 42312 203506 42340 206908
rect 42956 203574 42984 206908
rect 43600 203642 43628 206908
rect 43692 206894 44258 206922
rect 43588 203636 43640 203642
rect 43588 203578 43640 203584
rect 42944 203568 42996 203574
rect 42944 203510 42996 203516
rect 42300 203500 42352 203506
rect 42300 203442 42352 203448
rect 43692 203114 43720 206894
rect 44888 203438 44916 206908
rect 45060 203636 45112 203642
rect 45060 203578 45112 203584
rect 43772 203432 43824 203438
rect 43772 203374 43824 203380
rect 44876 203432 44928 203438
rect 44876 203374 44928 203380
rect 43140 203086 43720 203114
rect 43140 195686 43168 203086
rect 43680 203024 43732 203030
rect 43680 202966 43732 202972
rect 43692 195754 43720 202966
rect 43680 195748 43732 195754
rect 43680 195690 43732 195696
rect 43128 195680 43180 195686
rect 43128 195622 43180 195628
rect 43784 195618 43812 203374
rect 45072 196366 45100 203578
rect 45532 203506 45560 206908
rect 46176 203642 46204 206908
rect 46164 203636 46216 203642
rect 46164 203578 46216 203584
rect 45520 203500 45572 203506
rect 45520 203442 45572 203448
rect 45060 196360 45112 196366
rect 45060 196302 45112 196308
rect 50684 195822 50712 211087
rect 51144 210714 51172 211631
rect 51132 210708 51184 210714
rect 51132 210650 51184 210656
rect 50854 210608 50910 210617
rect 50854 210543 50910 210552
rect 50762 210064 50818 210073
rect 50762 209999 50818 210008
rect 50776 195958 50804 209999
rect 50764 195952 50816 195958
rect 50764 195894 50816 195900
rect 50868 195890 50896 210543
rect 52708 210306 52736 212010
rect 52892 211598 52920 213370
rect 58320 213337 58348 214458
rect 92716 214448 92768 214454
rect 92716 214390 92768 214396
rect 92728 213337 92756 214390
rect 92808 214380 92860 214386
rect 92808 214322 92860 214328
rect 92820 214017 92848 214322
rect 92806 214008 92862 214017
rect 92806 213943 92862 213952
rect 58306 213328 58362 213337
rect 52972 213292 53024 213298
rect 58306 213263 58362 213272
rect 92714 213328 92770 213337
rect 92714 213263 92770 213272
rect 52972 213234 53024 213240
rect 52984 211666 53012 213234
rect 97960 213224 98012 213230
rect 97960 213166 98012 213172
rect 58308 213088 58360 213094
rect 58308 213030 58360 213036
rect 93636 213088 93688 213094
rect 93636 213030 93688 213036
rect 58216 213020 58268 213026
rect 58216 212962 58268 212968
rect 58228 212793 58256 212962
rect 58214 212784 58270 212793
rect 58214 212719 58270 212728
rect 58320 212249 58348 213030
rect 92716 213020 92768 213026
rect 92716 212962 92768 212968
rect 92728 212793 92756 212962
rect 92714 212784 92770 212793
rect 92714 212719 92770 212728
rect 93648 212249 93676 213030
rect 58306 212240 58362 212249
rect 58306 212175 58362 212184
rect 93634 212240 93690 212249
rect 93634 212175 93690 212184
rect 56468 211932 56520 211938
rect 56468 211874 56520 211880
rect 52972 211660 53024 211666
rect 52972 211602 53024 211608
rect 52880 211592 52932 211598
rect 52880 211534 52932 211540
rect 56480 211122 56508 211874
rect 58216 211660 58268 211666
rect 58216 211602 58268 211608
rect 93544 211660 93596 211666
rect 93544 211602 93596 211608
rect 58228 211569 58256 211602
rect 58308 211592 58360 211598
rect 58214 211560 58270 211569
rect 92808 211592 92860 211598
rect 58308 211534 58360 211540
rect 92714 211560 92770 211569
rect 58214 211495 58270 211504
rect 56468 211116 56520 211122
rect 56468 211058 56520 211064
rect 58320 211025 58348 211534
rect 92808 211534 92860 211540
rect 92714 211495 92716 211504
rect 92768 211495 92770 211504
rect 92716 211466 92768 211472
rect 58400 211116 58452 211122
rect 58400 211058 58452 211064
rect 58306 211016 58362 211025
rect 58306 210951 58362 210960
rect 56284 210708 56336 210714
rect 56284 210650 56336 210656
rect 52696 210300 52748 210306
rect 52696 210242 52748 210248
rect 56296 209966 56324 210650
rect 58412 210345 58440 211058
rect 92820 211025 92848 211534
rect 92806 211016 92862 211025
rect 92806 210951 92862 210960
rect 92624 210368 92676 210374
rect 58398 210336 58454 210345
rect 58216 210300 58268 210306
rect 93556 210345 93584 211602
rect 97972 211530 98000 213166
rect 98064 213026 98092 214458
rect 98156 214386 98184 215818
rect 100994 215096 101050 215105
rect 100994 215031 101050 215040
rect 101008 214454 101036 215031
rect 100996 214448 101048 214454
rect 100996 214390 101048 214396
rect 98144 214380 98196 214386
rect 98144 214322 98196 214328
rect 100994 214008 101050 214017
rect 100994 213943 101050 213952
rect 98144 213156 98196 213162
rect 98144 213098 98196 213104
rect 98052 213020 98104 213026
rect 98052 212962 98104 212968
rect 98052 211796 98104 211802
rect 98052 211738 98104 211744
rect 97960 211524 98012 211530
rect 97960 211466 98012 211472
rect 94096 210504 94148 210510
rect 94096 210446 94148 210452
rect 94004 210436 94056 210442
rect 94004 210378 94056 210384
rect 92624 210310 92676 210316
rect 93542 210336 93598 210345
rect 58398 210271 58454 210280
rect 58216 210242 58268 210248
rect 56284 209960 56336 209966
rect 56284 209902 56336 209908
rect 58228 209801 58256 210242
rect 58308 209960 58360 209966
rect 58308 209902 58360 209908
rect 58214 209792 58270 209801
rect 58214 209727 58270 209736
rect 50946 209384 51002 209393
rect 50946 209319 51002 209328
rect 50960 196026 50988 209319
rect 58320 209257 58348 209902
rect 58306 209248 58362 209257
rect 58306 209183 58362 209192
rect 91244 209076 91296 209082
rect 91244 209018 91296 209024
rect 83056 209008 83108 209014
rect 61264 208934 61600 208962
rect 62980 208934 63316 208962
rect 64452 208934 64788 208962
rect 65832 208934 66168 208962
rect 67304 208934 67824 208962
rect 68684 208934 69204 208962
rect 70156 208934 70584 208962
rect 71536 208934 71964 208962
rect 51130 208840 51186 208849
rect 51130 208775 51186 208784
rect 51038 208296 51094 208305
rect 51038 208231 51094 208240
rect 51052 196094 51080 208231
rect 51144 207330 51172 208775
rect 51222 207752 51278 207761
rect 51222 207687 51224 207696
rect 51276 207687 51278 207696
rect 56100 207716 56152 207722
rect 51224 207658 51276 207664
rect 56100 207658 56152 207664
rect 51144 207302 51264 207330
rect 51130 207208 51186 207217
rect 51130 207143 51186 207152
rect 51040 196088 51092 196094
rect 51040 196030 51092 196036
rect 50948 196020 51000 196026
rect 50948 195962 51000 195968
rect 50856 195884 50908 195890
rect 50856 195826 50908 195832
rect 50672 195816 50724 195822
rect 50672 195758 50724 195764
rect 43772 195612 43824 195618
rect 43772 195554 43824 195560
rect 51144 195482 51172 207143
rect 51236 196162 51264 207302
rect 56112 196366 56140 207658
rect 61264 207518 61292 208934
rect 61252 207512 61304 207518
rect 61252 207454 61304 207460
rect 63288 206294 63316 208934
rect 63276 206288 63328 206294
rect 63276 206230 63328 206236
rect 64760 206226 64788 208934
rect 65116 206288 65168 206294
rect 65116 206230 65168 206236
rect 64748 206220 64800 206226
rect 64748 206162 64800 206168
rect 56100 196360 56152 196366
rect 56100 196302 56152 196308
rect 57572 196360 57624 196366
rect 57572 196302 57624 196308
rect 51224 196156 51276 196162
rect 51224 196098 51276 196104
rect 51132 195476 51184 195482
rect 51132 195418 51184 195424
rect 56468 195476 56520 195482
rect 56468 195418 56520 195424
rect 56480 193716 56508 195418
rect 57584 193716 57612 196302
rect 59780 196156 59832 196162
rect 59780 196098 59832 196104
rect 58676 196088 58728 196094
rect 58676 196030 58728 196036
rect 58688 193716 58716 196030
rect 59792 193716 59820 196098
rect 60884 196020 60936 196026
rect 60884 195962 60936 195968
rect 60896 193716 60924 195962
rect 61988 195952 62040 195958
rect 61988 195894 62040 195900
rect 62000 193716 62028 195894
rect 63092 195884 63144 195890
rect 63092 195826 63144 195832
rect 63104 193716 63132 195826
rect 64196 195816 64248 195822
rect 64196 195758 64248 195764
rect 64208 193716 64236 195758
rect 65128 193730 65156 206230
rect 66140 206226 66168 208934
rect 65208 206220 65260 206226
rect 65208 206162 65260 206168
rect 66128 206220 66180 206226
rect 66128 206162 66180 206168
rect 66588 206220 66640 206226
rect 66588 206162 66640 206168
rect 65220 194410 65248 206162
rect 65220 194382 65892 194410
rect 65128 193702 65326 193730
rect 65864 193594 65892 194382
rect 66600 193866 66628 206162
rect 67796 196366 67824 208934
rect 69176 206242 69204 208934
rect 69176 206214 69388 206242
rect 67784 196360 67836 196366
rect 67784 196302 67836 196308
rect 68612 196360 68664 196366
rect 68612 196302 68664 196308
rect 66600 193838 66996 193866
rect 66968 193594 66996 193838
rect 68624 193716 68652 196302
rect 69360 193866 69388 206214
rect 70556 195226 70584 208934
rect 71936 196314 71964 208934
rect 72672 208934 73008 208962
rect 74052 208934 74388 208962
rect 75524 208934 75860 208962
rect 76904 208934 77240 208962
rect 78376 208934 78712 208962
rect 78928 208934 80092 208962
rect 80308 208934 81564 208962
rect 81688 208934 82944 208962
rect 83056 208950 83108 208956
rect 84252 209008 84304 209014
rect 90600 209008 90652 209014
rect 84304 208956 84416 208962
rect 84252 208950 84416 208956
rect 72672 206226 72700 208934
rect 74052 206226 74080 208934
rect 75524 206226 75552 208934
rect 76904 206226 76932 208934
rect 78376 206226 78404 208934
rect 72108 206220 72160 206226
rect 72108 206162 72160 206168
rect 72660 206220 72712 206226
rect 72660 206162 72712 206168
rect 73396 206220 73448 206226
rect 73396 206162 73448 206168
rect 74040 206220 74092 206226
rect 74040 206162 74092 206168
rect 74776 206220 74828 206226
rect 74776 206162 74828 206168
rect 75512 206220 75564 206226
rect 75512 206162 75564 206168
rect 76156 206220 76208 206226
rect 76156 206162 76208 206168
rect 76892 206220 76944 206226
rect 76892 206162 76944 206168
rect 77536 206220 77588 206226
rect 77536 206162 77588 206168
rect 78364 206220 78416 206226
rect 78364 206162 78416 206168
rect 71936 196286 72056 196314
rect 70556 195198 70676 195226
rect 69360 193838 69572 193866
rect 69544 193730 69572 193838
rect 70648 193730 70676 195198
rect 69544 193702 69834 193730
rect 70648 193702 70938 193730
rect 72028 193716 72056 196286
rect 72120 193594 72148 206162
rect 73408 193594 73436 206162
rect 74788 193594 74816 206162
rect 76168 193730 76196 206162
rect 76168 193702 76458 193730
rect 77548 193716 77576 206162
rect 78928 195226 78956 208934
rect 80308 195226 80336 208934
rect 81688 196366 81716 208934
rect 83068 196366 83096 208950
rect 84264 208934 84416 208950
rect 85736 208934 85796 208962
rect 87268 208934 87604 208962
rect 90120 208934 90456 208962
rect 90600 208950 90652 208956
rect 85736 207489 85764 208934
rect 87576 207518 87604 208934
rect 87564 207512 87616 207518
rect 85722 207480 85778 207489
rect 87564 207454 87616 207460
rect 85722 207415 85778 207424
rect 90428 206566 90456 208934
rect 90416 206560 90468 206566
rect 90416 206502 90468 206508
rect 85724 206220 85776 206226
rect 85724 206162 85776 206168
rect 80848 196360 80900 196366
rect 80848 196302 80900 196308
rect 81676 196360 81728 196366
rect 81676 196302 81728 196308
rect 81952 196360 82004 196366
rect 81952 196302 82004 196308
rect 83056 196360 83108 196366
rect 83056 196302 83108 196308
rect 78836 195198 78956 195226
rect 80216 195198 80336 195226
rect 78836 193730 78864 195198
rect 80216 193730 80244 195198
rect 78666 193702 78864 193730
rect 79770 193702 80244 193730
rect 80860 193716 80888 196302
rect 81964 193716 81992 196302
rect 85736 193730 85764 206162
rect 90612 196366 90640 208950
rect 91152 206560 91204 206566
rect 91152 206502 91204 206508
rect 89772 196360 89824 196366
rect 89772 196302 89824 196308
rect 90600 196360 90652 196366
rect 90600 196302 90652 196308
rect 88668 195952 88720 195958
rect 88668 195894 88720 195900
rect 86460 195816 86512 195822
rect 86460 195758 86512 195764
rect 85382 193702 85764 193730
rect 86472 193716 86500 195758
rect 87564 195748 87616 195754
rect 87564 195690 87616 195696
rect 87576 193716 87604 195690
rect 88680 193716 88708 195894
rect 89784 193716 89812 196302
rect 91164 195890 91192 206502
rect 91152 195884 91204 195890
rect 91152 195826 91204 195832
rect 91256 193730 91284 209018
rect 92636 193866 92664 210310
rect 92716 210300 92768 210306
rect 93542 210271 93598 210280
rect 92716 210242 92768 210248
rect 92728 209801 92756 210242
rect 92714 209792 92770 209801
rect 92714 209727 92770 209736
rect 94016 196366 94044 210378
rect 94108 209257 94136 210446
rect 98064 210306 98092 211738
rect 98156 211598 98184 213098
rect 101008 213094 101036 213943
rect 101178 213464 101234 213473
rect 101178 213399 101234 213408
rect 101192 213230 101220 213399
rect 101180 213224 101232 213230
rect 101086 213192 101142 213201
rect 101180 213166 101232 213172
rect 101086 213127 101088 213136
rect 101140 213127 101142 213136
rect 101088 213098 101140 213104
rect 100996 213088 101048 213094
rect 100996 213030 101048 213036
rect 100994 212376 101050 212385
rect 100994 212311 101050 212320
rect 101008 211734 101036 212311
rect 101086 211968 101142 211977
rect 101086 211903 101142 211912
rect 101100 211802 101128 211903
rect 101088 211796 101140 211802
rect 101088 211738 101140 211744
rect 100996 211728 101048 211734
rect 100996 211670 101048 211676
rect 98144 211592 98196 211598
rect 98144 211534 98196 211540
rect 101178 211152 101234 211161
rect 101178 211087 101234 211096
rect 101086 210744 101142 210753
rect 101086 210679 101142 210688
rect 100994 210472 101050 210481
rect 101100 210442 101128 210679
rect 101192 210510 101220 211087
rect 101180 210504 101232 210510
rect 101180 210446 101232 210452
rect 100994 210407 101050 210416
rect 101088 210436 101140 210442
rect 101008 210374 101036 210407
rect 101088 210378 101140 210384
rect 100996 210368 101048 210374
rect 100996 210310 101048 210316
rect 98052 210300 98104 210306
rect 98052 210242 98104 210248
rect 101086 209520 101142 209529
rect 101086 209455 101142 209464
rect 94094 209248 94150 209257
rect 94094 209183 94150 209192
rect 100994 209112 101050 209121
rect 101100 209082 101128 209455
rect 100994 209047 101050 209056
rect 101088 209076 101140 209082
rect 101008 209014 101036 209047
rect 101088 209018 101140 209024
rect 100996 209008 101048 209014
rect 100996 208950 101048 208956
rect 101652 207518 101680 234071
rect 134298 233456 134354 233465
rect 134298 233391 134354 233400
rect 134312 232678 134340 233391
rect 134300 232672 134352 232678
rect 134300 232614 134352 232620
rect 134574 225976 134630 225985
rect 134574 225911 134630 225920
rect 134588 225606 134616 225911
rect 134576 225600 134628 225606
rect 134576 225542 134628 225548
rect 134482 222032 134538 222041
rect 134482 221967 134538 221976
rect 134496 221866 134524 221967
rect 134484 221860 134536 221866
rect 134484 221802 134536 221808
rect 101730 221488 101786 221497
rect 101730 221423 101786 221432
rect 101744 221322 101772 221423
rect 101732 221316 101784 221322
rect 101732 221258 101784 221264
rect 101730 220672 101786 220681
rect 101730 220607 101786 220616
rect 101744 219894 101772 220607
rect 101822 220264 101878 220273
rect 101822 220199 101878 220208
rect 101836 219962 101864 220199
rect 101914 219992 101970 220001
rect 101824 219956 101876 219962
rect 101914 219927 101970 219936
rect 101824 219898 101876 219904
rect 101732 219888 101784 219894
rect 101732 219830 101784 219836
rect 101730 219040 101786 219049
rect 101730 218975 101786 218984
rect 101744 218534 101772 218975
rect 101928 218602 101956 219927
rect 102006 218632 102062 218641
rect 101916 218596 101968 218602
rect 102006 218567 102062 218576
rect 101916 218538 101968 218544
rect 101732 218528 101784 218534
rect 101732 218470 101784 218476
rect 101914 217952 101970 217961
rect 101914 217887 101970 217896
rect 101822 217544 101878 217553
rect 101822 217479 101878 217488
rect 101836 217310 101864 217479
rect 101824 217304 101876 217310
rect 101730 217272 101786 217281
rect 101824 217246 101876 217252
rect 101730 217207 101732 217216
rect 101784 217207 101786 217216
rect 101732 217178 101784 217184
rect 101928 217174 101956 217887
rect 101916 217168 101968 217174
rect 101916 217110 101968 217116
rect 102020 217106 102048 218567
rect 102008 217100 102060 217106
rect 102008 217042 102060 217048
rect 101822 216184 101878 216193
rect 101822 216119 101878 216128
rect 101730 216048 101786 216057
rect 101730 215983 101786 215992
rect 101744 215882 101772 215983
rect 101732 215876 101784 215882
rect 101732 215818 101784 215824
rect 101836 215814 101864 216119
rect 101824 215808 101876 215814
rect 101824 215750 101876 215756
rect 101822 214960 101878 214969
rect 101822 214895 101878 214904
rect 101836 214522 101864 214895
rect 101824 214516 101876 214522
rect 101824 214458 101876 214464
rect 134666 214008 134722 214017
rect 134666 213943 134722 213952
rect 134680 213162 134708 213943
rect 134668 213156 134720 213162
rect 134668 213098 134720 213104
rect 102098 208432 102154 208441
rect 102098 208367 102154 208376
rect 101914 207888 101970 207897
rect 101914 207823 101970 207832
rect 101730 207616 101786 207625
rect 101730 207551 101786 207560
rect 101640 207512 101692 207518
rect 101640 207454 101692 207460
rect 100994 206528 101050 206537
rect 100994 206463 101050 206472
rect 101008 206226 101036 206463
rect 100996 206220 101048 206226
rect 100996 206162 101048 206168
rect 98972 204452 99024 204458
rect 98972 204394 99024 204400
rect 98880 203500 98932 203506
rect 98880 203442 98932 203448
rect 93084 196360 93136 196366
rect 93084 196302 93136 196308
rect 94004 196360 94056 196366
rect 94004 196302 94056 196308
rect 92268 193838 92664 193866
rect 92268 193730 92296 193838
rect 90902 193702 91284 193730
rect 92006 193702 92296 193730
rect 93096 193716 93124 196302
rect 94188 195884 94240 195890
rect 94188 195826 94240 195832
rect 94200 193716 94228 195826
rect 65864 193566 66430 193594
rect 66968 193566 67534 193594
rect 72120 193566 73146 193594
rect 73408 193566 74250 193594
rect 74788 193566 75354 193594
rect 41838 189256 41894 189265
rect 41760 189214 41838 189242
rect 41838 189191 41894 189200
rect 13410 185720 13466 185729
rect 13410 185655 13466 185664
rect 13424 185554 13452 185655
rect 13412 185548 13464 185554
rect 13412 185490 13464 185496
rect 16080 185548 16132 185554
rect 16080 185490 16132 185496
rect 13320 184052 13372 184058
rect 13320 183994 13372 184000
rect 16092 177190 16120 185490
rect 98892 185321 98920 203442
rect 98984 186545 99012 204394
rect 99432 204316 99484 204322
rect 99432 204258 99484 204264
rect 99248 204180 99300 204186
rect 99248 204122 99300 204128
rect 99156 203840 99208 203846
rect 99156 203782 99208 203788
rect 99064 203568 99116 203574
rect 99064 203510 99116 203516
rect 99076 187769 99104 203510
rect 99168 189537 99196 203782
rect 99260 190761 99288 204122
rect 99340 203636 99392 203642
rect 99340 203578 99392 203584
rect 99246 190752 99302 190761
rect 99246 190687 99302 190696
rect 99154 189528 99210 189537
rect 99154 189463 99210 189472
rect 99352 188993 99380 203578
rect 99444 192393 99472 204258
rect 99524 204112 99576 204118
rect 99524 204054 99576 204060
rect 99536 193753 99564 204054
rect 101744 195822 101772 207551
rect 101732 195816 101784 195822
rect 101732 195758 101784 195764
rect 101928 195754 101956 207823
rect 102112 195958 102140 208367
rect 134772 207518 134800 234479
rect 135402 234000 135458 234009
rect 135402 233935 135404 233944
rect 135456 233935 135458 233944
rect 142304 233964 142356 233970
rect 135404 233906 135456 233912
rect 142304 233906 142356 233912
rect 142316 233057 142344 233906
rect 142302 233048 142358 233057
rect 142302 232983 142358 232992
rect 135402 232912 135458 232921
rect 135402 232847 135458 232856
rect 135416 232746 135444 232847
rect 146548 232762 146576 235130
rect 156852 232762 156880 235198
rect 135404 232740 135456 232746
rect 135404 232682 135456 232688
rect 142212 232740 142264 232746
rect 146548 232734 146608 232762
rect 156544 232734 156880 232762
rect 159520 232762 159548 235266
rect 166236 232762 166264 235810
rect 169548 232762 169576 235878
rect 174056 235330 174084 241318
rect 208912 236616 208964 236622
rect 194926 236584 194982 236593
rect 208912 236558 208964 236564
rect 218296 236616 218348 236622
rect 218296 236558 218348 236564
rect 194926 236519 194982 236528
rect 173492 235324 173544 235330
rect 173492 235266 173544 235272
rect 174044 235324 174096 235330
rect 174044 235266 174096 235272
rect 173504 232762 173532 235266
rect 194940 234788 194968 236519
rect 208924 234788 208952 236558
rect 215720 235256 215772 235262
rect 215720 235198 215772 235204
rect 186002 234544 186058 234553
rect 186002 234479 186058 234488
rect 185082 234000 185138 234009
rect 185082 233935 185138 233944
rect 185096 233766 185124 233935
rect 177172 233760 177224 233766
rect 177172 233702 177224 233708
rect 185084 233760 185136 233766
rect 185084 233702 185136 233708
rect 177184 233057 177212 233702
rect 185174 233456 185230 233465
rect 185174 233391 185230 233400
rect 177170 233048 177226 233057
rect 177170 232983 177226 232992
rect 159520 232734 159856 232762
rect 166236 232734 166572 232762
rect 169548 232734 169884 232762
rect 173196 232734 173532 232762
rect 142212 232682 142264 232688
rect 135402 232232 135458 232241
rect 135402 232167 135458 232176
rect 134850 231688 134906 231697
rect 134850 231623 134906 231632
rect 134864 231522 134892 231623
rect 134852 231516 134904 231522
rect 134852 231458 134904 231464
rect 135310 231144 135366 231153
rect 135310 231079 135312 231088
rect 135364 231079 135366 231088
rect 135312 231050 135364 231056
rect 135416 231046 135444 232167
rect 139636 231516 139688 231522
rect 139636 231458 139688 231464
rect 136876 231108 136928 231114
rect 136876 231050 136928 231056
rect 135404 231040 135456 231046
rect 135404 230982 135456 230988
rect 135402 230600 135458 230609
rect 135402 230535 135458 230544
rect 135310 230056 135366 230065
rect 135310 229991 135312 230000
rect 135364 229991 135366 230000
rect 135312 229962 135364 229968
rect 135416 229686 135444 230535
rect 135404 229680 135456 229686
rect 135404 229622 135456 229628
rect 136888 229550 136916 231050
rect 139648 230638 139676 231458
rect 142224 231289 142252 232682
rect 142304 232672 142356 232678
rect 163554 232640 163610 232649
rect 142304 232614 142356 232620
rect 142316 231969 142344 232614
rect 163260 232598 163554 232626
rect 163554 232575 163610 232584
rect 182324 232536 182376 232542
rect 182324 232478 182376 232484
rect 177724 232400 177776 232406
rect 177724 232342 177776 232348
rect 177736 232241 177764 232342
rect 177722 232232 177778 232241
rect 177722 232167 177778 232176
rect 142302 231960 142358 231969
rect 142302 231895 142358 231904
rect 182336 231862 182364 232478
rect 185188 232474 185216 233391
rect 185266 232912 185322 232921
rect 185266 232847 185322 232856
rect 185280 232542 185308 232847
rect 185268 232536 185320 232542
rect 185268 232478 185320 232484
rect 185176 232468 185228 232474
rect 185176 232410 185228 232416
rect 185266 232232 185322 232241
rect 185266 232167 185322 232176
rect 177724 231856 177776 231862
rect 177724 231798 177776 231804
rect 182324 231856 182376 231862
rect 182324 231798 182376 231804
rect 177736 231561 177764 231798
rect 185174 231688 185230 231697
rect 185174 231623 185230 231632
rect 177722 231552 177778 231561
rect 177722 231487 177778 231496
rect 142210 231280 142266 231289
rect 142210 231215 142266 231224
rect 178276 231108 178328 231114
rect 178276 231050 178328 231056
rect 177724 230972 177776 230978
rect 177724 230914 177776 230920
rect 143684 230904 143736 230910
rect 143684 230846 143736 230852
rect 143696 230745 143724 230846
rect 143682 230736 143738 230745
rect 143682 230671 143738 230680
rect 139636 230632 139688 230638
rect 139636 230574 139688 230580
rect 142948 230632 143000 230638
rect 142948 230574 143000 230580
rect 142960 230201 142988 230574
rect 177736 230473 177764 230914
rect 178182 230872 178238 230881
rect 178288 230858 178316 231050
rect 185188 231046 185216 231623
rect 185280 231114 185308 232167
rect 185358 231144 185414 231153
rect 185268 231108 185320 231114
rect 185358 231079 185414 231088
rect 185268 231050 185320 231056
rect 185176 231040 185228 231046
rect 185176 230982 185228 230988
rect 178238 230830 178316 230858
rect 178182 230807 178238 230816
rect 185266 230600 185322 230609
rect 185266 230535 185322 230544
rect 177722 230464 177778 230473
rect 177722 230399 177778 230408
rect 142946 230192 143002 230201
rect 142946 230127 143002 230136
rect 185174 230056 185230 230065
rect 139636 230020 139688 230026
rect 185174 229991 185230 230000
rect 139636 229962 139688 229968
rect 136876 229544 136928 229550
rect 136876 229486 136928 229492
rect 139648 229482 139676 229962
rect 143592 229612 143644 229618
rect 143592 229554 143644 229560
rect 177632 229612 177684 229618
rect 177632 229554 177684 229560
rect 139636 229476 139688 229482
rect 139636 229418 139688 229424
rect 143500 229476 143552 229482
rect 143500 229418 143552 229424
rect 135402 229376 135458 229385
rect 135402 229311 135458 229320
rect 135310 228832 135366 228841
rect 135310 228767 135366 228776
rect 135324 228394 135352 228767
rect 135416 228462 135444 229311
rect 135404 228456 135456 228462
rect 135404 228398 135456 228404
rect 135312 228388 135364 228394
rect 135312 228330 135364 228336
rect 135404 228320 135456 228326
rect 135402 228288 135404 228297
rect 138164 228320 138216 228326
rect 135456 228288 135458 228297
rect 143512 228297 143540 229418
rect 143604 228977 143632 229554
rect 143684 229544 143736 229550
rect 143682 229512 143684 229521
rect 143736 229512 143738 229521
rect 143682 229447 143738 229456
rect 177644 229249 177672 229554
rect 185188 229550 185216 229991
rect 185280 229618 185308 230535
rect 185268 229612 185320 229618
rect 185268 229554 185320 229560
rect 177816 229544 177868 229550
rect 177816 229486 177868 229492
rect 185176 229544 185228 229550
rect 185176 229486 185228 229492
rect 177724 229476 177776 229482
rect 177724 229418 177776 229424
rect 177736 229385 177764 229418
rect 177722 229376 177778 229385
rect 177722 229311 177778 229320
rect 177630 229240 177686 229249
rect 177630 229175 177686 229184
rect 143590 228968 143646 228977
rect 143590 228903 143646 228912
rect 177828 228705 177856 229486
rect 185372 229482 185400 231079
rect 185360 229476 185412 229482
rect 185360 229418 185412 229424
rect 185634 229376 185690 229385
rect 185634 229311 185690 229320
rect 177814 228696 177870 228705
rect 177814 228631 177870 228640
rect 181128 228320 181180 228326
rect 138164 228262 138216 228268
rect 143498 228288 143554 228297
rect 135402 228223 135458 228232
rect 135402 227744 135458 227753
rect 135402 227679 135458 227688
rect 135310 227200 135366 227209
rect 135310 227135 135366 227144
rect 135324 226778 135352 227135
rect 135416 226898 135444 227679
rect 135404 226892 135456 226898
rect 135404 226834 135456 226840
rect 135324 226750 135536 226778
rect 138176 226762 138204 228262
rect 185176 228320 185228 228326
rect 181128 228262 181180 228268
rect 185174 228288 185176 228297
rect 185228 228288 185230 228297
rect 143498 228223 143554 228232
rect 143684 228252 143736 228258
rect 143684 228194 143736 228200
rect 177724 228252 177776 228258
rect 177724 228194 177776 228200
rect 143316 228184 143368 228190
rect 143316 228126 143368 228132
rect 143328 227209 143356 228126
rect 143696 227753 143724 228194
rect 177632 228184 177684 228190
rect 177632 228126 177684 228132
rect 143682 227744 143738 227753
rect 143682 227679 143738 227688
rect 177644 227481 177672 228126
rect 177736 228025 177764 228194
rect 177722 228016 177778 228025
rect 177722 227951 177778 227960
rect 177630 227472 177686 227481
rect 177630 227407 177686 227416
rect 143314 227200 143370 227209
rect 143314 227135 143370 227144
rect 143316 226824 143368 226830
rect 143316 226766 143368 226772
rect 177632 226824 177684 226830
rect 177632 226766 177684 226772
rect 135218 226520 135274 226529
rect 135218 226455 135274 226464
rect 135232 225538 135260 226455
rect 135220 225532 135272 225538
rect 135220 225474 135272 225480
rect 135508 225470 135536 226750
rect 138164 226756 138216 226762
rect 138164 226698 138216 226704
rect 143328 225985 143356 226766
rect 143684 226756 143736 226762
rect 143684 226698 143736 226704
rect 143696 226529 143724 226698
rect 143682 226520 143738 226529
rect 143682 226455 143738 226464
rect 177644 226257 177672 226766
rect 181140 226694 181168 228262
rect 185648 228258 185676 229311
rect 185910 228832 185966 228841
rect 185910 228767 185966 228776
rect 185174 228223 185230 228232
rect 185636 228252 185688 228258
rect 185636 228194 185688 228200
rect 185924 228190 185952 228767
rect 185912 228184 185964 228190
rect 185912 228126 185964 228132
rect 185174 227744 185230 227753
rect 185174 227679 185230 227688
rect 182324 226892 182376 226898
rect 182324 226834 182376 226840
rect 177724 226688 177776 226694
rect 177722 226656 177724 226665
rect 181128 226688 181180 226694
rect 177776 226656 177778 226665
rect 181128 226630 181180 226636
rect 177722 226591 177778 226600
rect 177630 226248 177686 226257
rect 177630 226183 177686 226192
rect 143314 225976 143370 225985
rect 143314 225911 143370 225920
rect 143500 225600 143552 225606
rect 143500 225542 143552 225548
rect 135496 225464 135548 225470
rect 135310 225432 135366 225441
rect 135496 225406 135548 225412
rect 135310 225367 135366 225376
rect 135218 224344 135274 224353
rect 135218 224279 135220 224288
rect 135272 224279 135274 224288
rect 135220 224250 135272 224256
rect 135324 224246 135352 225367
rect 135402 224888 135458 224897
rect 135402 224823 135458 224832
rect 135312 224240 135364 224246
rect 135312 224182 135364 224188
rect 135416 224178 135444 224823
rect 136876 224308 136928 224314
rect 136876 224250 136928 224256
rect 135404 224172 135456 224178
rect 135404 224114 135456 224120
rect 135402 223664 135458 223673
rect 135402 223599 135458 223608
rect 135310 223120 135366 223129
rect 135310 223055 135312 223064
rect 135364 223055 135366 223064
rect 135312 223026 135364 223032
rect 135416 222818 135444 223599
rect 135404 222812 135456 222818
rect 135404 222754 135456 222760
rect 136888 222682 136916 224250
rect 143512 224217 143540 225542
rect 143592 225532 143644 225538
rect 143592 225474 143644 225480
rect 143604 224761 143632 225474
rect 143684 225464 143736 225470
rect 143684 225406 143736 225412
rect 177632 225464 177684 225470
rect 177632 225406 177684 225412
rect 177722 225432 177778 225441
rect 143696 225305 143724 225406
rect 143682 225296 143738 225305
rect 143682 225231 143738 225240
rect 177644 225033 177672 225406
rect 177722 225367 177778 225376
rect 177816 225396 177868 225402
rect 177736 225334 177764 225367
rect 177816 225338 177868 225344
rect 177724 225328 177776 225334
rect 177724 225270 177776 225276
rect 177630 225024 177686 225033
rect 177630 224959 177686 224968
rect 143590 224752 143646 224761
rect 143590 224687 143646 224696
rect 177828 224489 177856 225338
rect 182336 225334 182364 226834
rect 185188 226830 185216 227679
rect 185266 227200 185322 227209
rect 185266 227135 185322 227144
rect 185280 226898 185308 227135
rect 185268 226892 185320 226898
rect 185268 226834 185320 226840
rect 185176 226824 185228 226830
rect 185176 226766 185228 226772
rect 185174 226520 185230 226529
rect 185174 226455 185230 226464
rect 185188 225470 185216 226455
rect 185266 225976 185322 225985
rect 185266 225911 185322 225920
rect 185176 225464 185228 225470
rect 185176 225406 185228 225412
rect 185280 225402 185308 225911
rect 185358 225432 185414 225441
rect 185268 225396 185320 225402
rect 185358 225367 185414 225376
rect 185268 225338 185320 225344
rect 182324 225328 182376 225334
rect 182324 225270 182376 225276
rect 185174 224888 185230 224897
rect 185174 224823 185230 224832
rect 177814 224480 177870 224489
rect 177814 224415 177870 224424
rect 143498 224208 143554 224217
rect 143498 224143 143554 224152
rect 143684 224104 143736 224110
rect 143684 224046 143736 224052
rect 177724 224104 177776 224110
rect 177724 224046 177776 224052
rect 143316 224036 143368 224042
rect 143316 223978 143368 223984
rect 137612 223084 137664 223090
rect 137612 223026 137664 223032
rect 136876 222676 136928 222682
rect 136876 222618 136928 222624
rect 134850 222576 134906 222585
rect 134850 222511 134906 222520
rect 134864 222410 134892 222511
rect 134852 222404 134904 222410
rect 134852 222346 134904 222352
rect 135310 221488 135366 221497
rect 135310 221423 135312 221432
rect 135364 221423 135366 221432
rect 136876 221452 136928 221458
rect 135312 221394 135364 221400
rect 136876 221394 136928 221400
rect 135402 220808 135458 220817
rect 135402 220743 135458 220752
rect 135310 220264 135366 220273
rect 135310 220199 135366 220208
rect 135324 220166 135352 220199
rect 135312 220160 135364 220166
rect 135312 220102 135364 220108
rect 135416 220030 135444 220743
rect 135404 220024 135456 220030
rect 135404 219966 135456 219972
rect 136888 219894 136916 221394
rect 137624 221322 137652 223026
rect 143328 222993 143356 223978
rect 143696 223537 143724 224046
rect 177356 224036 177408 224042
rect 177356 223978 177408 223984
rect 143682 223528 143738 223537
rect 143682 223463 143738 223472
rect 177368 223265 177396 223978
rect 177736 223809 177764 224046
rect 185188 224042 185216 224823
rect 185266 224344 185322 224353
rect 185266 224279 185322 224288
rect 185176 224036 185228 224042
rect 185176 223978 185228 223984
rect 177722 223800 177778 223809
rect 177722 223735 177778 223744
rect 185174 223664 185230 223673
rect 185174 223599 185230 223608
rect 177354 223256 177410 223265
rect 177354 223191 177410 223200
rect 143314 222984 143370 222993
rect 143314 222919 143370 222928
rect 185188 222750 185216 223599
rect 143316 222744 143368 222750
rect 143316 222686 143368 222692
rect 177632 222744 177684 222750
rect 177632 222686 177684 222692
rect 185176 222744 185228 222750
rect 185176 222686 185228 222692
rect 139728 222404 139780 222410
rect 139728 222346 139780 222352
rect 139636 221860 139688 221866
rect 139636 221802 139688 221808
rect 137612 221316 137664 221322
rect 137612 221258 137664 221264
rect 139648 220642 139676 221802
rect 139740 221186 139768 222346
rect 143328 221769 143356 222686
rect 143684 222676 143736 222682
rect 143684 222618 143736 222624
rect 143696 222313 143724 222618
rect 143682 222304 143738 222313
rect 143682 222239 143738 222248
rect 177644 222041 177672 222686
rect 185280 222682 185308 224279
rect 185372 224110 185400 225367
rect 185360 224104 185412 224110
rect 185360 224046 185412 224052
rect 185450 223120 185506 223129
rect 185450 223055 185506 223064
rect 177724 222676 177776 222682
rect 177724 222618 177776 222624
rect 185268 222676 185320 222682
rect 185268 222618 185320 222624
rect 177736 222449 177764 222618
rect 185266 222576 185322 222585
rect 185266 222511 185322 222520
rect 177722 222440 177778 222449
rect 177722 222375 177778 222384
rect 177630 222032 177686 222041
rect 177630 221967 177686 221976
rect 185174 222032 185230 222041
rect 185174 221967 185230 221976
rect 143314 221760 143370 221769
rect 143314 221695 143370 221704
rect 143684 221316 143736 221322
rect 143684 221258 143736 221264
rect 177632 221316 177684 221322
rect 177632 221258 177684 221264
rect 143696 221225 143724 221258
rect 143682 221216 143738 221225
rect 139728 221180 139780 221186
rect 139728 221122 139780 221128
rect 143592 221180 143644 221186
rect 143682 221151 143738 221160
rect 143592 221122 143644 221128
rect 139636 220636 139688 220642
rect 139636 220578 139688 220584
rect 143604 220545 143632 221122
rect 177644 220953 177672 221258
rect 185188 221254 185216 221967
rect 185280 221322 185308 222511
rect 185358 221488 185414 221497
rect 185358 221423 185414 221432
rect 185268 221316 185320 221322
rect 185268 221258 185320 221264
rect 177816 221248 177868 221254
rect 177816 221190 177868 221196
rect 185176 221248 185228 221254
rect 185176 221190 185228 221196
rect 177724 221180 177776 221186
rect 177724 221122 177776 221128
rect 177736 221089 177764 221122
rect 177722 221080 177778 221089
rect 177722 221015 177778 221024
rect 177630 220944 177686 220953
rect 177630 220879 177686 220888
rect 143684 220636 143736 220642
rect 143684 220578 143736 220584
rect 143590 220536 143646 220545
rect 143590 220471 143646 220480
rect 138164 220160 138216 220166
rect 138164 220102 138216 220108
rect 136876 219888 136928 219894
rect 136876 219830 136928 219836
rect 135402 219720 135458 219729
rect 135402 219655 135458 219664
rect 135034 219176 135090 219185
rect 135034 219111 135090 219120
rect 135048 218874 135076 219111
rect 135036 218868 135088 218874
rect 135036 218810 135088 218816
rect 135416 218738 135444 219655
rect 137520 218868 137572 218874
rect 137520 218810 137572 218816
rect 135404 218732 135456 218738
rect 135404 218674 135456 218680
rect 135312 218664 135364 218670
rect 135310 218632 135312 218641
rect 135364 218632 135366 218641
rect 135310 218567 135366 218576
rect 135402 217952 135458 217961
rect 135402 217887 135458 217896
rect 135416 217514 135444 217887
rect 135404 217508 135456 217514
rect 135404 217450 135456 217456
rect 135402 217408 135458 217417
rect 135402 217343 135404 217352
rect 135456 217343 135458 217352
rect 135404 217314 135456 217320
rect 137532 217174 137560 218810
rect 137980 218664 138032 218670
rect 137980 218606 138032 218612
rect 137704 217508 137756 217514
rect 137704 217450 137756 217456
rect 137612 217372 137664 217378
rect 137612 217314 137664 217320
rect 137520 217168 137572 217174
rect 137520 217110 137572 217116
rect 135402 216864 135458 216873
rect 135402 216799 135458 216808
rect 135416 215882 135444 216799
rect 135494 216320 135550 216329
rect 135494 216255 135550 216264
rect 135404 215876 135456 215882
rect 135404 215818 135456 215824
rect 135402 215776 135458 215785
rect 135402 215711 135458 215720
rect 134850 215096 134906 215105
rect 134850 215031 134906 215040
rect 134864 214930 134892 215031
rect 134852 214924 134904 214930
rect 134852 214866 134904 214872
rect 135312 214584 135364 214590
rect 135310 214552 135312 214561
rect 135364 214552 135366 214561
rect 135416 214522 135444 215711
rect 135310 214487 135366 214496
rect 135404 214516 135456 214522
rect 135404 214458 135456 214464
rect 135508 214454 135536 216255
rect 137624 215678 137652 217314
rect 137716 215746 137744 217450
rect 137992 217106 138020 218606
rect 138176 218534 138204 220102
rect 143696 220001 143724 220578
rect 177828 220273 177856 221190
rect 185174 220808 185230 220817
rect 185174 220743 185230 220752
rect 177814 220264 177870 220273
rect 177814 220199 177870 220208
rect 143682 219992 143738 220001
rect 143132 219956 143184 219962
rect 185188 219962 185216 220743
rect 143682 219927 143738 219936
rect 177632 219956 177684 219962
rect 143132 219898 143184 219904
rect 177632 219898 177684 219904
rect 185176 219956 185228 219962
rect 185176 219898 185228 219904
rect 143144 218777 143172 219898
rect 143684 219888 143736 219894
rect 143684 219830 143736 219836
rect 143696 219321 143724 219830
rect 143682 219312 143738 219321
rect 143682 219247 143738 219256
rect 177644 219049 177672 219898
rect 185372 219894 185400 221423
rect 185464 221186 185492 223055
rect 185452 221180 185504 221186
rect 185452 221122 185504 221128
rect 185542 220264 185598 220273
rect 185542 220199 185598 220208
rect 177724 219888 177776 219894
rect 177724 219830 177776 219836
rect 185360 219888 185412 219894
rect 185360 219830 185412 219836
rect 177736 219593 177764 219830
rect 177722 219584 177778 219593
rect 177722 219519 177778 219528
rect 177630 219040 177686 219049
rect 177630 218975 177686 218984
rect 143130 218768 143186 218777
rect 143130 218703 143186 218712
rect 185556 218602 185584 220199
rect 185726 219720 185782 219729
rect 185726 219655 185782 219664
rect 185634 219176 185690 219185
rect 185634 219111 185690 219120
rect 143500 218596 143552 218602
rect 143500 218538 143552 218544
rect 177724 218596 177776 218602
rect 177724 218538 177776 218544
rect 185544 218596 185596 218602
rect 185544 218538 185596 218544
rect 138164 218528 138216 218534
rect 138164 218470 138216 218476
rect 143512 217553 143540 218538
rect 143684 218528 143736 218534
rect 143684 218470 143736 218476
rect 177632 218528 177684 218534
rect 177632 218470 177684 218476
rect 143696 218233 143724 218470
rect 143682 218224 143738 218233
rect 143682 218159 143738 218168
rect 177644 217961 177672 218470
rect 177736 218369 177764 218538
rect 177722 218360 177778 218369
rect 177722 218295 177778 218304
rect 177630 217952 177686 217961
rect 177630 217887 177686 217896
rect 143498 217544 143554 217553
rect 143498 217479 143554 217488
rect 185542 217408 185598 217417
rect 185542 217343 185598 217352
rect 181036 217304 181088 217310
rect 181036 217246 181088 217252
rect 143684 217168 143736 217174
rect 177724 217168 177776 217174
rect 143684 217110 143736 217116
rect 177722 217136 177724 217145
rect 177776 217136 177778 217145
rect 137980 217100 138032 217106
rect 137980 217042 138032 217048
rect 143132 217100 143184 217106
rect 143132 217042 143184 217048
rect 143144 216329 143172 217042
rect 143696 217009 143724 217110
rect 177632 217100 177684 217106
rect 177722 217071 177778 217080
rect 177632 217042 177684 217048
rect 143682 217000 143738 217009
rect 143682 216935 143738 216944
rect 177644 216737 177672 217042
rect 177630 216728 177686 216737
rect 177630 216663 177686 216672
rect 143130 216320 143186 216329
rect 143130 216255 143186 216264
rect 143500 215808 143552 215814
rect 143130 215776 143186 215785
rect 137704 215740 137756 215746
rect 143500 215750 143552 215756
rect 177632 215808 177684 215814
rect 177632 215750 177684 215756
rect 143130 215711 143132 215720
rect 137704 215682 137756 215688
rect 143184 215711 143186 215720
rect 143132 215682 143184 215688
rect 137612 215672 137664 215678
rect 137612 215614 137664 215620
rect 142948 215672 143000 215678
rect 142948 215614 143000 215620
rect 142960 215241 142988 215614
rect 142946 215232 143002 215241
rect 142946 215167 143002 215176
rect 137612 214924 137664 214930
rect 137612 214866 137664 214872
rect 136876 214584 136928 214590
rect 136876 214526 136928 214532
rect 135496 214448 135548 214454
rect 135496 214390 135548 214396
rect 135402 213464 135458 213473
rect 135402 213399 135404 213408
rect 135456 213399 135458 213408
rect 135404 213370 135456 213376
rect 136888 213026 136916 214526
rect 137520 213428 137572 213434
rect 137520 213370 137572 213376
rect 136968 213156 137020 213162
rect 136968 213098 137020 213104
rect 136876 213020 136928 213026
rect 136876 212962 136928 212968
rect 134850 212920 134906 212929
rect 134850 212855 134906 212864
rect 134864 211938 134892 212855
rect 135402 212240 135458 212249
rect 135402 212175 135458 212184
rect 135416 212074 135444 212175
rect 135404 212068 135456 212074
rect 135404 212010 135456 212016
rect 134852 211932 134904 211938
rect 134852 211874 134904 211880
rect 135402 211696 135458 211705
rect 136980 211666 137008 213098
rect 135402 211631 135458 211640
rect 136968 211660 137020 211666
rect 135034 211152 135090 211161
rect 135034 211087 135090 211096
rect 134850 210608 134906 210617
rect 134850 210543 134906 210552
rect 134760 207512 134812 207518
rect 134760 207454 134812 207460
rect 104228 203506 104256 206908
rect 104780 204458 104808 206908
rect 104768 204452 104820 204458
rect 104768 204394 104820 204400
rect 105332 203574 105360 206908
rect 105884 203642 105912 206908
rect 106436 203846 106464 206908
rect 106988 204186 107016 206908
rect 107540 204322 107568 206908
rect 107528 204316 107580 204322
rect 107528 204258 107580 204264
rect 106976 204180 107028 204186
rect 106976 204122 107028 204128
rect 108092 204118 108120 206908
rect 108080 204112 108132 204118
rect 108080 204054 108132 204060
rect 106424 203840 106476 203846
rect 106424 203782 106476 203788
rect 105872 203636 105924 203642
rect 105872 203578 105924 203584
rect 105320 203568 105372 203574
rect 105320 203510 105372 203516
rect 104216 203500 104268 203506
rect 104216 203442 104268 203448
rect 108644 203438 108672 206908
rect 109196 203522 109224 206908
rect 109196 203494 109408 203522
rect 108632 203432 108684 203438
rect 108632 203374 108684 203380
rect 109276 203432 109328 203438
rect 109276 203374 109328 203380
rect 102100 195952 102152 195958
rect 102100 195894 102152 195900
rect 101916 195748 101968 195754
rect 101916 195690 101968 195696
rect 109288 193866 109316 203374
rect 109380 196366 109408 203494
rect 109748 203438 109776 206908
rect 110300 203506 110328 206908
rect 110288 203500 110340 203506
rect 110288 203442 110340 203448
rect 109736 203432 109788 203438
rect 109736 203374 109788 203380
rect 110852 203114 110880 206908
rect 111024 203500 111076 203506
rect 111024 203442 111076 203448
rect 110932 203432 110984 203438
rect 110932 203374 110984 203380
rect 110668 203086 110880 203114
rect 109368 196360 109420 196366
rect 109368 196302 109420 196308
rect 110288 196360 110340 196366
rect 110288 196302 110340 196308
rect 109288 193838 109776 193866
rect 99522 193744 99578 193753
rect 109748 193730 109776 193838
rect 110300 193730 110328 196302
rect 110668 195754 110696 203086
rect 110944 202978 110972 203374
rect 110760 202950 110972 202978
rect 110656 195748 110708 195754
rect 110656 195690 110708 195696
rect 110760 193730 110788 202950
rect 111036 202842 111064 203442
rect 111496 203438 111524 206908
rect 111484 203432 111536 203438
rect 111484 203374 111536 203380
rect 110852 202814 111064 202842
rect 110852 194138 110880 202814
rect 111668 195748 111720 195754
rect 111668 195690 111720 195696
rect 110852 194110 110972 194138
rect 109748 193702 110130 193730
rect 110300 193702 110498 193730
rect 110760 193702 110866 193730
rect 99522 193679 99578 193688
rect 110944 193594 110972 194110
rect 111680 193716 111708 195690
rect 112048 195482 112076 206908
rect 112312 203432 112364 203438
rect 112312 203374 112364 203380
rect 112036 195476 112088 195482
rect 112036 195418 112088 195424
rect 112324 193730 112352 203374
rect 112496 195476 112548 195482
rect 112496 195418 112548 195424
rect 112062 193702 112352 193730
rect 112508 193716 112536 195418
rect 112600 193730 112628 206908
rect 113152 193730 113180 206908
rect 112600 193702 112890 193730
rect 113152 193702 113258 193730
rect 113704 193716 113732 206908
rect 114256 193730 114284 206908
rect 114808 203522 114836 206908
rect 114716 203494 114836 203522
rect 114716 193730 114744 203494
rect 115256 196428 115308 196434
rect 115256 196370 115308 196376
rect 114888 196360 114940 196366
rect 114888 196302 114940 196308
rect 114086 193702 114284 193730
rect 114454 193702 114744 193730
rect 114900 193716 114928 196302
rect 115268 193716 115296 196370
rect 115360 196366 115388 206908
rect 115912 196434 115940 206908
rect 116084 203500 116136 203506
rect 116084 203442 116136 203448
rect 115992 203432 116044 203438
rect 115992 203374 116044 203380
rect 115900 196428 115952 196434
rect 115900 196370 115952 196376
rect 115348 196360 115400 196366
rect 115348 196302 115400 196308
rect 116004 193730 116032 203374
rect 115650 193702 116032 193730
rect 116096 193716 116124 203442
rect 116464 203438 116492 206908
rect 117016 203506 117044 206908
rect 117568 203522 117596 206908
rect 117004 203500 117056 203506
rect 117004 203442 117056 203448
rect 117384 203494 117596 203522
rect 117648 203500 117700 203506
rect 116452 203432 116504 203438
rect 116452 203374 116504 203380
rect 117280 203432 117332 203438
rect 117280 203374 117332 203380
rect 117292 196366 117320 203374
rect 116820 196360 116872 196366
rect 116820 196302 116872 196308
rect 117280 196360 117332 196366
rect 117280 196302 117332 196308
rect 116452 195612 116504 195618
rect 116452 195554 116504 195560
rect 116464 193716 116492 195554
rect 116832 193716 116860 196302
rect 117384 195618 117412 203494
rect 117648 203442 117700 203448
rect 117660 203386 117688 203442
rect 118212 203438 118240 206908
rect 118568 203568 118620 203574
rect 118568 203510 118620 203516
rect 117476 203358 117688 203386
rect 118200 203432 118252 203438
rect 118200 203374 118252 203380
rect 117372 195612 117424 195618
rect 117372 195554 117424 195560
rect 117476 193730 117504 203358
rect 117648 196020 117700 196026
rect 117648 195962 117700 195968
rect 117306 193702 117504 193730
rect 117660 193716 117688 195962
rect 118580 195754 118608 203510
rect 118764 203506 118792 206908
rect 118752 203500 118804 203506
rect 118752 203442 118804 203448
rect 118844 203500 118896 203506
rect 118844 203442 118896 203448
rect 118660 203432 118712 203438
rect 118660 203374 118712 203380
rect 118672 196026 118700 203374
rect 118752 203364 118804 203370
rect 118752 203306 118804 203312
rect 118660 196020 118712 196026
rect 118660 195962 118712 195968
rect 118108 195748 118160 195754
rect 118108 195690 118160 195696
rect 118568 195748 118620 195754
rect 118568 195690 118620 195696
rect 118120 193716 118148 195690
rect 118764 193730 118792 203306
rect 118502 193702 118792 193730
rect 118856 193716 118884 203442
rect 119316 203438 119344 206908
rect 119868 203574 119896 206908
rect 120224 204452 120276 204458
rect 120224 204394 120276 204400
rect 120132 203636 120184 203642
rect 120132 203578 120184 203584
rect 119856 203568 119908 203574
rect 119856 203510 119908 203516
rect 120040 203568 120092 203574
rect 120040 203510 120092 203516
rect 119304 203432 119356 203438
rect 119304 203374 119356 203380
rect 120052 196434 120080 203510
rect 119672 196428 119724 196434
rect 119672 196370 119724 196376
rect 120040 196428 120092 196434
rect 120040 196370 120092 196376
rect 119304 196360 119356 196366
rect 119304 196302 119356 196308
rect 119316 193716 119344 196302
rect 119684 193716 119712 196370
rect 120144 193730 120172 203578
rect 120236 196366 120264 204394
rect 120420 203438 120448 206908
rect 120972 203506 121000 206908
rect 121420 204656 121472 204662
rect 121420 204598 121472 204604
rect 120960 203500 121012 203506
rect 120960 203442 121012 203448
rect 120408 203432 120460 203438
rect 120408 203374 120460 203380
rect 120224 196360 120276 196366
rect 120224 196302 120276 196308
rect 120868 196360 120920 196366
rect 120868 196302 120920 196308
rect 120500 195544 120552 195550
rect 120500 195486 120552 195492
rect 120066 193702 120172 193730
rect 120512 193716 120540 195486
rect 120880 193716 120908 196302
rect 121432 193730 121460 204598
rect 121524 204458 121552 206908
rect 121512 204452 121564 204458
rect 121512 204394 121564 204400
rect 121512 204316 121564 204322
rect 121512 204258 121564 204264
rect 121524 195550 121552 204258
rect 121604 204248 121656 204254
rect 121604 204190 121656 204196
rect 121616 196366 121644 204190
rect 122076 203574 122104 206908
rect 122628 203642 122656 206908
rect 123180 204322 123208 206908
rect 123168 204316 123220 204322
rect 123168 204258 123220 204264
rect 123732 204254 123760 206908
rect 124284 204662 124312 206908
rect 124272 204656 124324 204662
rect 124272 204598 124324 204604
rect 123720 204248 123772 204254
rect 123720 204190 123772 204196
rect 124272 203840 124324 203846
rect 124272 203782 124324 203788
rect 123720 203772 123772 203778
rect 123720 203714 123772 203720
rect 122616 203636 122668 203642
rect 122616 203578 122668 203584
rect 122064 203568 122116 203574
rect 122064 203510 122116 203516
rect 122892 196496 122944 196502
rect 122892 196438 122944 196444
rect 121604 196360 121656 196366
rect 121604 196302 121656 196308
rect 122432 196224 122484 196230
rect 122432 196166 122484 196172
rect 122064 196088 122116 196094
rect 122064 196030 122116 196036
rect 121696 196020 121748 196026
rect 121696 195962 121748 195968
rect 121512 195544 121564 195550
rect 121512 195486 121564 195492
rect 121262 193702 121460 193730
rect 121708 193716 121736 195962
rect 122076 193716 122104 196030
rect 122444 193716 122472 196166
rect 122904 193716 122932 196438
rect 123628 196428 123680 196434
rect 123628 196370 123680 196376
rect 123260 196360 123312 196366
rect 123260 196302 123312 196308
rect 123272 193716 123300 196302
rect 123640 193716 123668 196370
rect 123732 196094 123760 203714
rect 124180 203704 124232 203710
rect 124180 203646 124232 203652
rect 123996 203636 124048 203642
rect 123996 203578 124048 203584
rect 123904 203568 123956 203574
rect 123904 203510 123956 203516
rect 123812 203500 123864 203506
rect 123812 203442 123864 203448
rect 123720 196088 123772 196094
rect 123720 196030 123772 196036
rect 123824 196026 123852 203442
rect 123916 196230 123944 203510
rect 124008 196502 124036 203578
rect 123996 196496 124048 196502
rect 123996 196438 124048 196444
rect 124192 196366 124220 203646
rect 124180 196360 124232 196366
rect 124180 196302 124232 196308
rect 123904 196224 123956 196230
rect 123904 196166 123956 196172
rect 123812 196020 123864 196026
rect 123812 195962 123864 195968
rect 124284 193730 124312 203782
rect 124836 203506 124864 206908
rect 125480 203778 125508 206908
rect 125468 203772 125520 203778
rect 125468 203714 125520 203720
rect 126032 203574 126060 206908
rect 126584 203642 126612 206908
rect 127136 203710 127164 206908
rect 127124 203704 127176 203710
rect 127124 203646 127176 203652
rect 126572 203636 126624 203642
rect 126572 203578 126624 203584
rect 126020 203568 126072 203574
rect 126020 203510 126072 203516
rect 124824 203500 124876 203506
rect 124824 203442 124876 203448
rect 127688 203438 127716 206908
rect 128240 203846 128268 206908
rect 128228 203840 128280 203846
rect 128228 203782 128280 203788
rect 127860 203636 127912 203642
rect 127860 203578 127912 203584
rect 124364 203432 124416 203438
rect 124364 203374 124416 203380
rect 127676 203432 127728 203438
rect 127676 203374 127728 203380
rect 124376 196434 124404 203374
rect 124364 196428 124416 196434
rect 124364 196370 124416 196376
rect 125652 196428 125704 196434
rect 125652 196370 125704 196376
rect 125284 196360 125336 196366
rect 125284 196302 125336 196308
rect 124456 195816 124508 195822
rect 124456 195758 124508 195764
rect 124114 193702 124312 193730
rect 124468 193716 124496 195758
rect 124824 195612 124876 195618
rect 124824 195554 124876 195560
rect 124836 193716 124864 195554
rect 125296 193716 125324 196302
rect 125664 193716 125692 196370
rect 127872 196366 127900 203578
rect 128044 203568 128096 203574
rect 128044 203510 128096 203516
rect 127952 203500 128004 203506
rect 127952 203442 128004 203448
rect 127860 196360 127912 196366
rect 127860 196302 127912 196308
rect 127964 195618 127992 203442
rect 128056 196434 128084 203510
rect 128792 203438 128820 206908
rect 129344 203506 129372 206908
rect 129896 203642 129924 206908
rect 129884 203636 129936 203642
rect 129884 203578 129936 203584
rect 130448 203574 130476 206908
rect 130436 203568 130488 203574
rect 130436 203510 130488 203516
rect 129332 203500 129384 203506
rect 129332 203442 129384 203448
rect 128136 203432 128188 203438
rect 128136 203374 128188 203380
rect 128780 203432 128832 203438
rect 128780 203374 128832 203380
rect 128044 196428 128096 196434
rect 128044 196370 128096 196376
rect 128148 195822 128176 203374
rect 134864 195890 134892 210543
rect 134942 209384 134998 209393
rect 134942 209319 134998 209328
rect 134956 196026 134984 209319
rect 134944 196020 134996 196026
rect 134944 195962 134996 195968
rect 134852 195884 134904 195890
rect 134852 195826 134904 195832
rect 135048 195822 135076 211087
rect 135416 210374 135444 211631
rect 136968 211602 137020 211608
rect 137532 211394 137560 213370
rect 137624 213094 137652 214866
rect 143512 214561 143540 215750
rect 177644 214969 177672 215750
rect 181048 215678 181076 217246
rect 185556 217242 185584 217343
rect 181220 217236 181272 217242
rect 181220 217178 181272 217184
rect 185544 217236 185596 217242
rect 185544 217178 185596 217184
rect 181128 215876 181180 215882
rect 181128 215818 181180 215824
rect 177724 215672 177776 215678
rect 177722 215640 177724 215649
rect 181036 215672 181088 215678
rect 177776 215640 177778 215649
rect 181036 215614 181088 215620
rect 177722 215575 177778 215584
rect 177724 215536 177776 215542
rect 177724 215478 177776 215484
rect 177736 215377 177764 215478
rect 177722 215368 177778 215377
rect 177722 215303 177778 215312
rect 177630 214960 177686 214969
rect 177630 214895 177686 214904
rect 143498 214552 143554 214561
rect 143498 214487 143554 214496
rect 143684 214516 143736 214522
rect 143684 214458 143736 214464
rect 181036 214516 181088 214522
rect 181036 214458 181088 214464
rect 142948 214448 143000 214454
rect 142948 214390 143000 214396
rect 142960 214017 142988 214390
rect 142946 214008 143002 214017
rect 142946 213943 143002 213952
rect 143696 213337 143724 214458
rect 177632 214448 177684 214454
rect 177632 214390 177684 214396
rect 177644 213745 177672 214390
rect 177724 214312 177776 214318
rect 177724 214254 177776 214260
rect 177736 214153 177764 214254
rect 177722 214144 177778 214153
rect 177722 214079 177778 214088
rect 177630 213736 177686 213745
rect 177630 213671 177686 213680
rect 143682 213328 143738 213337
rect 143682 213263 143738 213272
rect 181048 213094 181076 214458
rect 181140 214318 181168 215818
rect 181232 215542 181260 217178
rect 185648 217174 185676 219111
rect 185740 218534 185768 219655
rect 186016 218670 186044 234479
rect 215732 230745 215760 235198
rect 216916 235188 216968 235194
rect 216916 235130 216968 235136
rect 215718 230736 215774 230745
rect 215718 230671 215774 230680
rect 185820 218664 185872 218670
rect 186004 218664 186056 218670
rect 185820 218606 185872 218612
rect 185910 218632 185966 218641
rect 185728 218528 185780 218534
rect 185728 218470 185780 218476
rect 185726 217952 185782 217961
rect 185726 217887 185782 217896
rect 185740 217310 185768 217887
rect 185728 217304 185780 217310
rect 185728 217246 185780 217252
rect 185636 217168 185688 217174
rect 185636 217110 185688 217116
rect 185726 216320 185782 216329
rect 185726 216255 185782 216264
rect 185740 215882 185768 216255
rect 185728 215876 185780 215882
rect 185728 215818 185780 215824
rect 185634 215776 185690 215785
rect 185634 215711 185690 215720
rect 181220 215536 181272 215542
rect 181220 215478 181272 215484
rect 181220 214584 181272 214590
rect 185268 214584 185320 214590
rect 181220 214526 181272 214532
rect 185266 214552 185268 214561
rect 185320 214552 185322 214561
rect 181128 214312 181180 214318
rect 181128 214254 181180 214260
rect 137612 213088 137664 213094
rect 137612 213030 137664 213036
rect 143684 213088 143736 213094
rect 143684 213030 143736 213036
rect 177724 213088 177776 213094
rect 177724 213030 177776 213036
rect 181036 213088 181088 213094
rect 181036 213030 181088 213036
rect 143500 213020 143552 213026
rect 143500 212962 143552 212968
rect 143512 212249 143540 212962
rect 143696 212793 143724 213030
rect 177736 212929 177764 213030
rect 177722 212920 177778 212929
rect 177722 212855 177778 212864
rect 143682 212784 143738 212793
rect 143682 212719 143738 212728
rect 181232 212550 181260 214526
rect 185266 214487 185322 214496
rect 185648 214454 185676 215711
rect 185726 215096 185782 215105
rect 185726 215031 185782 215040
rect 185740 214522 185768 215031
rect 185728 214516 185780 214522
rect 185728 214458 185780 214464
rect 185636 214448 185688 214454
rect 185636 214390 185688 214396
rect 185726 214008 185782 214017
rect 185726 213943 185782 213952
rect 185174 213464 185230 213473
rect 185174 213399 185230 213408
rect 185188 213230 185216 213399
rect 181956 213224 182008 213230
rect 181956 213166 182008 213172
rect 185176 213224 185228 213230
rect 185176 213166 185228 213172
rect 181864 213156 181916 213162
rect 181864 213098 181916 213104
rect 177724 212544 177776 212550
rect 177724 212486 177776 212492
rect 181220 212544 181272 212550
rect 181220 212486 181272 212492
rect 177736 212385 177764 212486
rect 177722 212376 177778 212385
rect 177722 212311 177778 212320
rect 143498 212240 143554 212249
rect 143498 212175 143554 212184
rect 137612 212068 137664 212074
rect 137612 212010 137664 212016
rect 137520 211388 137572 211394
rect 137520 211330 137572 211336
rect 135404 210368 135456 210374
rect 135404 210310 135456 210316
rect 137624 210238 137652 212010
rect 139636 211932 139688 211938
rect 139636 211874 139688 211880
rect 139648 210986 139676 211874
rect 181680 211728 181732 211734
rect 177722 211696 177778 211705
rect 143684 211660 143736 211666
rect 181680 211670 181732 211676
rect 177722 211631 177724 211640
rect 143684 211602 143736 211608
rect 177776 211631 177778 211640
rect 177724 211602 177776 211608
rect 143696 211569 143724 211602
rect 143682 211560 143738 211569
rect 143682 211495 143738 211504
rect 143684 211388 143736 211394
rect 143684 211330 143736 211336
rect 143696 211025 143724 211330
rect 177724 211320 177776 211326
rect 177724 211262 177776 211268
rect 177736 211161 177764 211262
rect 177722 211152 177778 211161
rect 177722 211087 177778 211096
rect 177724 211048 177776 211054
rect 143682 211016 143738 211025
rect 139636 210980 139688 210986
rect 139636 210922 139688 210928
rect 143592 210980 143644 210986
rect 177724 210990 177776 210996
rect 143682 210951 143738 210960
rect 143592 210922 143644 210928
rect 143604 210345 143632 210922
rect 177736 210753 177764 210990
rect 177722 210744 177778 210753
rect 177722 210679 177778 210688
rect 178276 210504 178328 210510
rect 178276 210446 178328 210452
rect 178092 210436 178144 210442
rect 178092 210378 178144 210384
rect 176804 210368 176856 210374
rect 143590 210336 143646 210345
rect 176804 210310 176856 210316
rect 143590 210271 143646 210280
rect 143684 210300 143736 210306
rect 143684 210242 143736 210248
rect 137612 210232 137664 210238
rect 137612 210174 137664 210180
rect 142948 210232 143000 210238
rect 142948 210174 143000 210180
rect 135126 210064 135182 210073
rect 135126 209999 135182 210008
rect 135140 195958 135168 209999
rect 142960 209801 142988 210174
rect 142946 209792 143002 209801
rect 142946 209727 143002 209736
rect 143696 209257 143724 210242
rect 143682 209248 143738 209257
rect 143682 209183 143738 209192
rect 175424 209076 175476 209082
rect 175424 209018 175476 209024
rect 174780 209008 174832 209014
rect 169902 208976 169958 208985
rect 145352 208934 145596 208962
rect 146976 208934 147312 208962
rect 148448 208934 148784 208962
rect 149828 208934 150164 208962
rect 151300 208934 152004 208962
rect 152680 208934 153016 208962
rect 154152 208934 154764 208962
rect 135310 208840 135366 208849
rect 135310 208775 135366 208784
rect 135218 208296 135274 208305
rect 135218 208231 135274 208240
rect 135232 196094 135260 208231
rect 135324 207466 135352 208775
rect 135402 207752 135458 207761
rect 135402 207687 135458 207696
rect 135416 207654 135444 207687
rect 135404 207648 135456 207654
rect 135404 207590 135456 207596
rect 140280 207648 140332 207654
rect 140280 207590 140332 207596
rect 135324 207438 135444 207466
rect 135310 207208 135366 207217
rect 135310 207143 135366 207152
rect 135220 196088 135272 196094
rect 135220 196030 135272 196036
rect 135128 195952 135180 195958
rect 135128 195894 135180 195900
rect 128136 195816 128188 195822
rect 128136 195758 128188 195764
rect 135036 195816 135088 195822
rect 135036 195758 135088 195764
rect 135324 195618 135352 207143
rect 135416 195754 135444 207438
rect 140292 196366 140320 207590
rect 145352 207518 145380 208934
rect 145340 207512 145392 207518
rect 145340 207454 145392 207460
rect 147284 206226 147312 208934
rect 148756 206838 148784 208934
rect 148744 206832 148796 206838
rect 148744 206774 148796 206780
rect 149388 206832 149440 206838
rect 149388 206774 149440 206780
rect 147272 206220 147324 206226
rect 147272 206162 147324 206168
rect 149296 206220 149348 206226
rect 149296 206162 149348 206168
rect 140280 196360 140332 196366
rect 140280 196302 140332 196308
rect 141568 196360 141620 196366
rect 141568 196302 141620 196308
rect 135404 195748 135456 195754
rect 135404 195690 135456 195696
rect 127952 195612 128004 195618
rect 127952 195554 128004 195560
rect 135312 195612 135364 195618
rect 135312 195554 135364 195560
rect 140464 195612 140516 195618
rect 140464 195554 140516 195560
rect 140476 193716 140504 195554
rect 141580 193716 141608 196302
rect 142672 196088 142724 196094
rect 142672 196030 142724 196036
rect 142684 193716 142712 196030
rect 144880 196020 144932 196026
rect 144880 195962 144932 195968
rect 143776 195748 143828 195754
rect 143776 195690 143828 195696
rect 143788 193716 143816 195690
rect 144892 193716 144920 195962
rect 145984 195952 146036 195958
rect 145984 195894 146036 195900
rect 145996 193716 146024 195894
rect 147088 195884 147140 195890
rect 147088 195826 147140 195832
rect 147100 193716 147128 195826
rect 148192 195816 148244 195822
rect 148192 195758 148244 195764
rect 148204 193716 148232 195758
rect 149308 193716 149336 206162
rect 149400 194818 149428 206774
rect 150136 206226 150164 208934
rect 150124 206220 150176 206226
rect 150124 206162 150176 206168
rect 150768 206220 150820 206226
rect 150768 206162 150820 206168
rect 149400 194790 150164 194818
rect 150136 193730 150164 194790
rect 150780 193866 150808 206162
rect 151976 196178 152004 208934
rect 152988 206226 153016 208934
rect 152976 206220 153028 206226
rect 152976 206162 153028 206168
rect 153528 206220 153580 206226
rect 153528 206162 153580 206168
rect 151976 196150 152096 196178
rect 150780 193838 151268 193866
rect 151240 193730 151268 193838
rect 152068 193730 152096 196150
rect 153540 193730 153568 206162
rect 154736 195226 154764 208934
rect 154920 208934 155532 208962
rect 156668 208934 157004 208962
rect 158048 208934 158384 208962
rect 159520 208934 159856 208962
rect 160900 208934 161236 208962
rect 161728 208934 162708 208962
rect 163108 208934 164088 208962
rect 164488 208934 165560 208962
rect 165868 208934 166940 208962
rect 167248 208934 168412 208962
rect 169792 208934 169902 208962
rect 154736 195198 154856 195226
rect 154828 193730 154856 195198
rect 154920 194818 154948 208934
rect 156668 206226 156696 208934
rect 158048 206226 158076 208934
rect 159520 206226 159548 208934
rect 160900 206226 160928 208934
rect 156196 206220 156248 206226
rect 156196 206162 156248 206168
rect 156656 206220 156708 206226
rect 156656 206162 156708 206168
rect 157576 206220 157628 206226
rect 157576 206162 157628 206168
rect 158036 206220 158088 206226
rect 158036 206162 158088 206168
rect 158956 206220 159008 206226
rect 158956 206162 159008 206168
rect 159508 206220 159560 206226
rect 159508 206162 159560 206168
rect 160336 206220 160388 206226
rect 160336 206162 160388 206168
rect 160888 206220 160940 206226
rect 160888 206162 160940 206168
rect 154920 194790 155500 194818
rect 150136 193702 150426 193730
rect 151240 193702 151530 193730
rect 152068 193702 152634 193730
rect 153540 193702 153830 193730
rect 154828 193702 154934 193730
rect 155472 193594 155500 194790
rect 156208 193594 156236 206162
rect 157588 193594 157616 206162
rect 158968 193730 158996 206162
rect 160348 193730 160376 206162
rect 161728 195226 161756 208934
rect 163108 195226 163136 208934
rect 164488 196366 164516 208934
rect 165868 196366 165896 208934
rect 163740 196360 163792 196366
rect 163740 196302 163792 196308
rect 164476 196360 164528 196366
rect 164476 196302 164528 196308
rect 164844 196360 164896 196366
rect 164844 196302 164896 196308
rect 165856 196360 165908 196366
rect 165856 196302 165908 196308
rect 161636 195198 161756 195226
rect 163016 195198 163136 195226
rect 161636 193730 161664 195198
rect 163016 193730 163044 195198
rect 158968 193702 159350 193730
rect 160348 193702 160454 193730
rect 161558 193702 161664 193730
rect 162662 193702 163044 193730
rect 163752 193716 163780 196302
rect 164856 193716 164884 196302
rect 167248 196298 167276 208934
rect 169902 208911 169958 208920
rect 171204 208934 171264 208962
rect 172584 208934 172644 208962
rect 174056 208934 174116 208962
rect 174780 208950 174832 208956
rect 171204 207518 171232 208934
rect 171192 207512 171244 207518
rect 171192 207454 171244 207460
rect 172584 206974 172612 208934
rect 174056 207450 174084 208934
rect 174044 207444 174096 207450
rect 174044 207386 174096 207392
rect 172572 206968 172624 206974
rect 172572 206910 172624 206916
rect 169904 206220 169956 206226
rect 169904 206162 169956 206168
rect 165948 196292 166000 196298
rect 165948 196234 166000 196240
rect 167236 196292 167288 196298
rect 167236 196234 167288 196240
rect 165960 193716 165988 196234
rect 167142 195240 167198 195249
rect 167142 195175 167198 195184
rect 167156 193716 167184 195175
rect 169916 193594 169944 206162
rect 174792 196366 174820 208950
rect 173768 196360 173820 196366
rect 173768 196302 173820 196308
rect 174780 196360 174832 196366
rect 174780 196302 174832 196308
rect 172664 195952 172716 195958
rect 172664 195894 172716 195900
rect 171560 195884 171612 195890
rect 171560 195826 171612 195832
rect 170456 195816 170508 195822
rect 170456 195758 170508 195764
rect 170468 193716 170496 195758
rect 171572 193716 171600 195826
rect 172676 193716 172704 195894
rect 173780 193716 173808 196302
rect 175436 193866 175464 209018
rect 176816 196366 176844 210310
rect 177724 210096 177776 210102
rect 177724 210038 177776 210044
rect 177736 209937 177764 210038
rect 177722 209928 177778 209937
rect 177722 209863 177778 209872
rect 178104 208826 178132 210378
rect 178182 209520 178238 209529
rect 178288 209506 178316 210446
rect 181692 210102 181720 211670
rect 181876 211666 181904 213098
rect 181864 211660 181916 211666
rect 181864 211602 181916 211608
rect 181968 211326 181996 213166
rect 185740 213162 185768 213943
rect 185728 213156 185780 213162
rect 185728 213098 185780 213104
rect 185726 212920 185782 212929
rect 185726 212855 185782 212864
rect 185740 211802 185768 212855
rect 182140 211796 182192 211802
rect 182140 211738 182192 211744
rect 185728 211796 185780 211802
rect 185728 211738 185780 211744
rect 181956 211320 182008 211326
rect 181956 211262 182008 211268
rect 182152 211054 182180 211738
rect 185726 211696 185782 211705
rect 185726 211631 185782 211640
rect 182140 211048 182192 211054
rect 182140 210990 182192 210996
rect 185740 210510 185768 211631
rect 185832 211274 185860 218606
rect 186004 218606 186056 218612
rect 185910 218567 185966 218576
rect 185924 217106 185952 218567
rect 185912 217100 185964 217106
rect 185912 217042 185964 217048
rect 185910 216864 185966 216873
rect 185910 216799 185966 216808
rect 185924 215814 185952 216799
rect 185912 215808 185964 215814
rect 185912 215750 185964 215756
rect 185910 212240 185966 212249
rect 185910 212175 185966 212184
rect 185924 211734 185952 212175
rect 185912 211728 185964 211734
rect 185912 211670 185964 211676
rect 216928 211569 216956 235130
rect 218308 232406 218336 236558
rect 218296 232400 218348 232406
rect 218296 232342 218348 232348
rect 222344 232400 222396 232406
rect 222344 232342 222396 232348
rect 222356 231697 222384 232342
rect 222342 231688 222398 231697
rect 222342 231623 222398 231632
rect 220318 220808 220374 220817
rect 220318 220743 220374 220752
rect 216914 211560 216970 211569
rect 216914 211495 216970 211504
rect 185832 211246 185952 211274
rect 185818 211152 185874 211161
rect 185818 211087 185874 211096
rect 185728 210504 185780 210510
rect 185728 210446 185780 210452
rect 185832 210442 185860 211087
rect 185820 210436 185872 210442
rect 185820 210378 185872 210384
rect 181680 210096 181732 210102
rect 181680 210038 181732 210044
rect 185726 210064 185782 210073
rect 185726 209999 185782 210008
rect 178238 209478 178316 209506
rect 178182 209455 178238 209464
rect 185740 209082 185768 209999
rect 185818 209384 185874 209393
rect 185818 209319 185874 209328
rect 185728 209076 185780 209082
rect 185728 209018 185780 209024
rect 185832 209014 185860 209319
rect 185820 209008 185872 209014
rect 185820 208950 185872 208956
rect 178104 208798 178224 208826
rect 177540 206968 177592 206974
rect 177540 206910 177592 206916
rect 175976 196360 176028 196366
rect 175976 196302 176028 196308
rect 176804 196360 176856 196366
rect 176804 196302 176856 196308
rect 177080 196360 177132 196366
rect 177080 196302 177132 196308
rect 175252 193838 175464 193866
rect 175252 193730 175280 193838
rect 174898 193702 175280 193730
rect 175988 193716 176016 196302
rect 177092 193716 177120 196302
rect 177552 195346 177580 206910
rect 178196 196366 178224 208798
rect 185924 207518 185952 211246
rect 186002 210608 186058 210617
rect 186002 210543 186058 210552
rect 186016 210374 186044 210543
rect 186004 210368 186056 210374
rect 186004 210310 186056 210316
rect 186094 208840 186150 208849
rect 186094 208775 186150 208784
rect 186002 207752 186058 207761
rect 186002 207687 186058 207696
rect 185912 207512 185964 207518
rect 185912 207454 185964 207460
rect 185174 207208 185230 207217
rect 185174 207143 185230 207152
rect 185188 206226 185216 207143
rect 185176 206220 185228 206226
rect 185176 206162 185228 206168
rect 183612 204180 183664 204186
rect 183612 204122 183664 204128
rect 183428 204112 183480 204118
rect 183428 204054 183480 204060
rect 183336 203704 183388 203710
rect 183336 203646 183388 203652
rect 183244 203636 183296 203642
rect 183244 203578 183296 203584
rect 183152 203568 183204 203574
rect 183152 203510 183204 203516
rect 183060 203500 183112 203506
rect 183060 203442 183112 203448
rect 178184 196360 178236 196366
rect 178184 196302 178236 196308
rect 177540 195340 177592 195346
rect 177540 195282 177592 195288
rect 179288 195340 179340 195346
rect 179288 195282 179340 195288
rect 179300 193716 179328 195282
rect 110944 193566 111326 193594
rect 155472 193566 156038 193594
rect 156208 193566 157142 193594
rect 157588 193566 158246 193594
rect 169378 193566 169944 193594
rect 182876 193232 182928 193238
rect 182874 193200 182876 193209
rect 182928 193200 182930 193209
rect 182874 193135 182930 193144
rect 105778 192520 105834 192529
rect 105778 192455 105834 192464
rect 99430 192384 99486 192393
rect 99430 192319 99486 192328
rect 99338 188984 99394 188993
rect 99338 188919 99394 188928
rect 99062 187760 99118 187769
rect 99062 187695 99118 187704
rect 99432 186908 99484 186914
rect 99432 186850 99484 186856
rect 98970 186536 99026 186545
rect 98970 186471 99026 186480
rect 98878 185312 98934 185321
rect 98878 185247 98934 185256
rect 22336 184052 22388 184058
rect 22336 183994 22388 184000
rect 22348 183825 22376 183994
rect 22334 183816 22390 183825
rect 22334 183751 22390 183760
rect 98604 182692 98656 182698
rect 98604 182634 98656 182640
rect 98616 182465 98644 182634
rect 98602 182456 98658 182465
rect 98602 182391 98658 182400
rect 99444 181105 99472 186850
rect 104400 184120 104452 184126
rect 104400 184062 104452 184068
rect 99524 184052 99576 184058
rect 99524 183994 99576 184000
rect 99536 183689 99564 183994
rect 99522 183680 99578 183689
rect 99522 183615 99578 183624
rect 99430 181096 99486 181105
rect 99430 181031 99486 181040
rect 98420 179904 98472 179910
rect 98420 179846 98472 179852
rect 99522 179872 99578 179881
rect 98432 179337 98460 179846
rect 99522 179807 99578 179816
rect 99536 179570 99564 179807
rect 104412 179570 104440 184062
rect 105792 184058 105820 192455
rect 107158 190208 107214 190217
rect 107158 190143 107214 190152
rect 106790 187896 106846 187905
rect 106790 187831 106846 187840
rect 106804 186914 106832 187831
rect 106792 186908 106844 186914
rect 106792 186850 106844 186856
rect 106790 185448 106846 185457
rect 106790 185383 106846 185392
rect 106804 184126 106832 185383
rect 106792 184120 106844 184126
rect 106792 184062 106844 184068
rect 105780 184052 105832 184058
rect 105780 183994 105832 184000
rect 107172 183258 107200 190143
rect 183072 184641 183100 203442
rect 183164 185865 183192 203510
rect 183256 187089 183284 203578
rect 183348 189537 183376 203646
rect 183440 190761 183468 204054
rect 183520 203432 183572 203438
rect 183520 203374 183572 203380
rect 183426 190752 183482 190761
rect 183426 190687 183482 190696
rect 183334 189528 183390 189537
rect 183334 189463 183390 189472
rect 183532 188313 183560 203374
rect 183624 191985 183652 204122
rect 186016 203522 186044 207687
rect 185924 203494 186044 203522
rect 185924 195822 185952 203494
rect 186108 195958 186136 208775
rect 186278 208296 186334 208305
rect 186278 208231 186334 208240
rect 186096 195952 186148 195958
rect 186096 195894 186148 195900
rect 186292 195890 186320 208231
rect 187936 207444 187988 207450
rect 187936 207386 187988 207392
rect 187948 206945 187976 207386
rect 200828 207030 201302 207058
rect 187934 206936 187990 206945
rect 187934 206871 187990 206880
rect 187200 203772 187252 203778
rect 187200 203714 187252 203720
rect 186280 195884 186332 195890
rect 186280 195826 186332 195832
rect 185912 195816 185964 195822
rect 185912 195758 185964 195764
rect 187212 193238 187240 203714
rect 188132 203506 188160 206908
rect 188592 203574 188620 206908
rect 189144 203642 189172 206908
rect 189132 203636 189184 203642
rect 189132 203578 189184 203584
rect 188580 203568 188632 203574
rect 188580 203510 188632 203516
rect 188120 203500 188172 203506
rect 188120 203442 188172 203448
rect 189696 203438 189724 206908
rect 190248 203710 190276 206908
rect 190800 204118 190828 206908
rect 191352 204186 191380 206908
rect 191340 204180 191392 204186
rect 191340 204122 191392 204128
rect 190788 204112 190840 204118
rect 190788 204054 190840 204060
rect 191904 203778 191932 206908
rect 191984 204112 192036 204118
rect 191984 204054 192036 204060
rect 191892 203772 191944 203778
rect 191892 203714 191944 203720
rect 190236 203704 190288 203710
rect 190236 203646 190288 203652
rect 189684 203432 189736 203438
rect 189684 203374 189736 203380
rect 187200 193232 187252 193238
rect 187200 193174 187252 193180
rect 191996 192801 192024 204054
rect 192456 203438 192484 206908
rect 193022 206894 193312 206922
rect 192444 203432 192496 203438
rect 192444 203374 192496 203380
rect 193284 196026 193312 206894
rect 193560 203438 193588 206908
rect 194126 206894 194600 206922
rect 194678 206894 194784 206922
rect 193364 203432 193416 203438
rect 193364 203374 193416 203380
rect 193548 203432 193600 203438
rect 193548 203374 193600 203380
rect 193272 196020 193324 196026
rect 193272 195962 193324 195968
rect 193376 195226 193404 203374
rect 194572 196366 194600 206894
rect 194652 203432 194704 203438
rect 194652 203374 194704 203380
rect 194560 196360 194612 196366
rect 194560 196302 194612 196308
rect 194664 196314 194692 203374
rect 194756 196434 194784 206894
rect 194848 206894 195230 206922
rect 195782 206894 196164 206922
rect 194848 196502 194876 206894
rect 194836 196496 194888 196502
rect 194836 196438 194888 196444
rect 196032 196496 196084 196502
rect 196032 196438 196084 196444
rect 194744 196428 194796 196434
rect 194744 196370 194796 196376
rect 195664 196428 195716 196434
rect 195664 196370 195716 196376
rect 195296 196360 195348 196366
rect 194664 196286 194876 196314
rect 195296 196302 195348 196308
rect 194468 196020 194520 196026
rect 194468 195962 194520 195968
rect 193376 195198 193680 195226
rect 193652 193730 193680 195198
rect 193652 193702 194126 193730
rect 194480 193716 194508 195962
rect 194848 193716 194876 196286
rect 195308 193716 195336 196302
rect 195676 193716 195704 196370
rect 196044 193716 196072 196438
rect 196136 195226 196164 206894
rect 196136 195198 196256 195226
rect 196228 193730 196256 195198
rect 196320 194002 196348 206908
rect 196412 206894 196886 206922
rect 197438 206894 197544 206922
rect 196412 196366 196440 206894
rect 196400 196360 196452 196366
rect 196400 196302 196452 196308
rect 197228 196360 197280 196366
rect 197228 196302 197280 196308
rect 196320 193974 196624 194002
rect 196596 193730 196624 193974
rect 196228 193702 196518 193730
rect 196596 193702 196886 193730
rect 197240 193716 197268 196302
rect 197516 195226 197544 206894
rect 197700 206894 197990 206922
rect 198160 206894 198542 206922
rect 198988 206894 199094 206922
rect 199264 206894 199646 206922
rect 199816 206894 200198 206922
rect 200368 206894 200750 206922
rect 197596 199556 197648 199562
rect 197596 199498 197648 199504
rect 197608 196366 197636 199498
rect 197596 196360 197648 196366
rect 197596 196302 197648 196308
rect 197516 195198 197636 195226
rect 197608 193730 197636 195198
rect 197700 194138 197728 206894
rect 198160 199562 198188 206894
rect 198988 203522 199016 206894
rect 198896 203494 199016 203522
rect 198148 199556 198200 199562
rect 198148 199498 198200 199504
rect 198424 196360 198476 196366
rect 198424 196302 198476 196308
rect 197700 194110 197820 194138
rect 197792 193730 197820 194110
rect 197608 193702 197714 193730
rect 197792 193702 198082 193730
rect 198436 193716 198464 196302
rect 198896 193716 198924 203494
rect 199160 203092 199212 203098
rect 199160 203034 199212 203040
rect 199172 196366 199200 203034
rect 199160 196360 199212 196366
rect 199160 196302 199212 196308
rect 199264 193716 199292 206894
rect 199816 203098 199844 206894
rect 200368 204474 200396 206894
rect 200276 204446 200396 204474
rect 199804 203092 199856 203098
rect 199804 203034 199856 203040
rect 199620 196360 199672 196366
rect 199620 196302 199672 196308
rect 199632 193716 199660 196302
rect 200276 193730 200304 204446
rect 200828 199306 200856 207030
rect 201748 206894 201854 206922
rect 201552 203636 201604 203642
rect 201552 203578 201604 203584
rect 201460 203432 201512 203438
rect 201460 203374 201512 203380
rect 200552 199278 200856 199306
rect 200552 193730 200580 199278
rect 200816 196020 200868 196026
rect 200816 195962 200868 195968
rect 200106 193702 200304 193730
rect 200474 193702 200580 193730
rect 200828 193716 200856 195962
rect 201472 193730 201500 203374
rect 201302 193702 201500 193730
rect 201564 193730 201592 203578
rect 201748 203488 201776 206894
rect 201656 203460 201776 203488
rect 201656 196026 201684 203460
rect 202300 203438 202328 206908
rect 202852 203642 202880 206908
rect 203128 206894 203418 206922
rect 202840 203636 202892 203642
rect 202840 203578 202892 203584
rect 203128 203522 203156 206894
rect 202852 203494 203156 203522
rect 202288 203432 202340 203438
rect 202288 203374 202340 203380
rect 202472 196360 202524 196366
rect 202472 196302 202524 196308
rect 202104 196156 202156 196162
rect 202104 196098 202156 196104
rect 201644 196020 201696 196026
rect 201644 195962 201696 195968
rect 201564 193702 201670 193730
rect 202116 193716 202144 196098
rect 202484 193716 202512 196302
rect 202852 196162 202880 203494
rect 203956 203438 203984 206908
rect 204312 203636 204364 203642
rect 204312 203578 204364 203584
rect 202932 203432 202984 203438
rect 202932 203374 202984 203380
rect 203024 203432 203076 203438
rect 203024 203374 203076 203380
rect 203944 203432 203996 203438
rect 203944 203374 203996 203380
rect 204220 203432 204272 203438
rect 204220 203374 204272 203380
rect 202840 196156 202892 196162
rect 202840 196098 202892 196104
rect 202944 193730 202972 203374
rect 203036 196366 203064 203374
rect 203668 196428 203720 196434
rect 203668 196370 203720 196376
rect 203024 196360 203076 196366
rect 203024 196302 203076 196308
rect 203300 196360 203352 196366
rect 203300 196302 203352 196308
rect 202866 193702 202972 193730
rect 203312 193716 203340 196302
rect 203680 193716 203708 196370
rect 204232 196366 204260 203374
rect 204220 196360 204272 196366
rect 204220 196302 204272 196308
rect 204324 193730 204352 203578
rect 204508 203574 204536 206908
rect 204496 203568 204548 203574
rect 204496 203510 204548 203516
rect 204404 203500 204456 203506
rect 204404 203442 204456 203448
rect 204416 196434 204444 203442
rect 205060 203438 205088 206908
rect 205416 204724 205468 204730
rect 205416 204666 205468 204672
rect 205428 203438 205456 204666
rect 205508 203568 205560 203574
rect 205508 203510 205560 203516
rect 205048 203432 205100 203438
rect 205048 203374 205100 203380
rect 205416 203432 205468 203438
rect 205416 203374 205468 203380
rect 204404 196428 204456 196434
rect 204404 196370 204456 196376
rect 204864 196360 204916 196366
rect 204864 196302 204916 196308
rect 204496 195952 204548 195958
rect 204496 195894 204548 195900
rect 204062 193702 204352 193730
rect 204508 193716 204536 195894
rect 204876 193716 204904 196302
rect 205520 193730 205548 203510
rect 205612 203506 205640 206908
rect 206164 203642 206192 206908
rect 206152 203636 206204 203642
rect 206152 203578 206204 203584
rect 205600 203500 205652 203506
rect 205600 203442 205652 203448
rect 205692 203500 205744 203506
rect 205692 203442 205744 203448
rect 205600 203364 205652 203370
rect 205600 203306 205652 203312
rect 205258 193702 205548 193730
rect 205612 193730 205640 203306
rect 205704 196366 205732 203442
rect 206716 203438 206744 206908
rect 207268 203506 207296 206908
rect 207820 203574 207848 206908
rect 208372 204730 208400 206908
rect 208360 204724 208412 204730
rect 208360 204666 208412 204672
rect 208360 204588 208412 204594
rect 208360 204530 208412 204536
rect 208268 204452 208320 204458
rect 208268 204394 208320 204400
rect 207808 203568 207860 203574
rect 207808 203510 207860 203516
rect 207900 203568 207952 203574
rect 207900 203510 207952 203516
rect 207256 203500 207308 203506
rect 207256 203442 207308 203448
rect 205784 203432 205836 203438
rect 205784 203374 205836 203380
rect 206704 203432 206756 203438
rect 206704 203374 206756 203380
rect 205692 196360 205744 196366
rect 205692 196302 205744 196308
rect 205796 195958 205824 203374
rect 206888 196360 206940 196366
rect 206888 196302 206940 196308
rect 205784 195952 205836 195958
rect 205784 195894 205836 195900
rect 206060 195952 206112 195958
rect 206060 195894 206112 195900
rect 205612 193702 205718 193730
rect 206072 193716 206100 195894
rect 206428 195340 206480 195346
rect 206428 195282 206480 195288
rect 206440 193716 206468 195282
rect 206900 193716 206928 196302
rect 207256 196156 207308 196162
rect 207256 196098 207308 196104
rect 207268 193716 207296 196098
rect 207912 195346 207940 203510
rect 208084 203500 208136 203506
rect 208084 203442 208136 203448
rect 207992 203432 208044 203438
rect 207992 203374 208044 203380
rect 208004 195958 208032 203374
rect 208096 196366 208124 203442
rect 208084 196360 208136 196366
rect 208084 196302 208136 196308
rect 208280 196162 208308 204394
rect 208268 196156 208320 196162
rect 208268 196098 208320 196104
rect 207992 195952 208044 195958
rect 207992 195894 208044 195900
rect 207900 195340 207952 195346
rect 207900 195282 207952 195288
rect 208372 194274 208400 204530
rect 208544 204520 208596 204526
rect 208544 204462 208596 204468
rect 208452 204248 208504 204254
rect 208452 204190 208504 204196
rect 208004 194246 208400 194274
rect 208004 193730 208032 194246
rect 208464 194138 208492 204190
rect 208372 194110 208492 194138
rect 208372 193730 208400 194110
rect 208556 193730 208584 204462
rect 208924 203438 208952 206908
rect 209476 203574 209504 206908
rect 209464 203568 209516 203574
rect 209464 203510 209516 203516
rect 210028 203506 210056 206908
rect 210580 204458 210608 206908
rect 211132 204594 211160 206908
rect 211120 204588 211172 204594
rect 211120 204530 211172 204536
rect 210568 204452 210620 204458
rect 210568 204394 210620 204400
rect 211684 204254 211712 206908
rect 212236 204526 212264 206908
rect 212802 206894 213000 206922
rect 212224 204520 212276 204526
rect 212224 204462 212276 204468
rect 211672 204248 211724 204254
rect 211672 204190 211724 204196
rect 210016 203500 210068 203506
rect 210016 203442 210068 203448
rect 208912 203432 208964 203438
rect 208912 203374 208964 203380
rect 212868 203092 212920 203098
rect 212868 203034 212920 203040
rect 209280 195952 209332 195958
rect 209280 195894 209332 195900
rect 208820 195884 208872 195890
rect 208820 195826 208872 195832
rect 207650 193702 208032 193730
rect 208110 193702 208400 193730
rect 208478 193702 208584 193730
rect 208832 193716 208860 195826
rect 209292 193716 209320 195894
rect 212880 195822 212908 203034
rect 212972 195890 213000 206894
rect 213064 206894 213354 206922
rect 213616 206894 213906 206922
rect 213064 195958 213092 206894
rect 213616 203098 213644 206894
rect 214444 204118 214472 206908
rect 214432 204112 214484 204118
rect 214432 204054 214484 204060
rect 213604 203092 213656 203098
rect 213604 203034 213656 203040
rect 213052 195952 213104 195958
rect 213052 195894 213104 195900
rect 212960 195884 213012 195890
rect 212960 195826 213012 195832
rect 209648 195816 209700 195822
rect 209648 195758 209700 195764
rect 212868 195816 212920 195822
rect 212868 195758 212920 195764
rect 209660 193716 209688 195758
rect 191982 192792 192038 192801
rect 191982 192727 192038 192736
rect 183610 191976 183666 191985
rect 183610 191911 183666 191920
rect 209752 190846 209964 190874
rect 191982 188712 192038 188721
rect 191982 188647 192038 188656
rect 183518 188304 183574 188313
rect 191996 188274 192024 188647
rect 183518 188239 183574 188248
rect 187936 188268 187988 188274
rect 187936 188210 187988 188216
rect 191984 188268 192036 188274
rect 191984 188210 192036 188216
rect 183242 187080 183298 187089
rect 183242 187015 183298 187024
rect 183150 185856 183206 185865
rect 183150 185791 183206 185800
rect 183058 184632 183114 184641
rect 183058 184567 183114 184576
rect 187948 184058 187976 188210
rect 191154 186808 191210 186817
rect 191154 186743 191210 186752
rect 182876 184052 182928 184058
rect 182876 183994 182928 184000
rect 187936 184052 187988 184058
rect 187936 183994 187988 184000
rect 128502 183816 128558 183825
rect 128502 183751 128558 183760
rect 106988 183230 107200 183258
rect 104492 182760 104544 182766
rect 104492 182702 104544 182708
rect 104504 179910 104532 182702
rect 106988 182698 107016 183230
rect 107158 183136 107214 183145
rect 107158 183071 107214 183080
rect 107172 182766 107200 183071
rect 128516 182766 128544 183751
rect 182888 183417 182916 183994
rect 182874 183408 182930 183417
rect 182874 183343 182930 183352
rect 107160 182760 107212 182766
rect 107160 182702 107212 182708
rect 128504 182760 128556 182766
rect 128504 182702 128556 182708
rect 137520 182760 137572 182766
rect 137520 182702 137572 182708
rect 190602 182728 190658 182737
rect 106976 182692 107028 182698
rect 106976 182634 107028 182640
rect 106974 180824 107030 180833
rect 106974 180759 107030 180768
rect 106988 180386 107016 180759
rect 105136 180380 105188 180386
rect 105136 180322 105188 180328
rect 106976 180380 107028 180386
rect 106976 180322 107028 180328
rect 104492 179904 104544 179910
rect 104492 179846 104544 179852
rect 99524 179564 99576 179570
rect 99524 179506 99576 179512
rect 104400 179564 104452 179570
rect 104400 179506 104452 179512
rect 98418 179328 98474 179337
rect 98418 179263 98474 179272
rect 44414 178784 44470 178793
rect 44414 178719 44470 178728
rect 44428 178618 44456 178719
rect 44416 178612 44468 178618
rect 44416 178554 44468 178560
rect 49292 178612 49344 178618
rect 49292 178554 49344 178560
rect 16080 177184 16132 177190
rect 22336 177184 22388 177190
rect 16080 177126 16132 177132
rect 22334 177152 22336 177161
rect 22388 177152 22390 177161
rect 22334 177087 22390 177096
rect 49304 174402 49332 178554
rect 99522 177424 99578 177433
rect 105148 177394 105176 180322
rect 106790 178376 106846 178385
rect 106790 178311 106846 178320
rect 99522 177359 99524 177368
rect 99576 177359 99578 177368
rect 105136 177388 105188 177394
rect 99524 177330 99576 177336
rect 105136 177330 105188 177336
rect 106804 177190 106832 178311
rect 98604 177184 98656 177190
rect 98604 177126 98656 177132
rect 106792 177184 106844 177190
rect 106792 177126 106844 177132
rect 98616 176753 98644 177126
rect 98602 176744 98658 176753
rect 98602 176679 98658 176688
rect 106606 176064 106662 176073
rect 106606 175999 106662 176008
rect 106620 175830 106648 175999
rect 98236 175824 98288 175830
rect 98236 175766 98288 175772
rect 106608 175824 106660 175830
rect 106608 175766 106660 175772
rect 98248 175393 98276 175766
rect 98234 175384 98290 175393
rect 98234 175319 98290 175328
rect 137532 174441 137560 182702
rect 183152 182692 183204 182698
rect 191168 182698 191196 186743
rect 191982 184768 192038 184777
rect 191982 184703 192038 184712
rect 190602 182663 190658 182672
rect 191156 182692 191208 182698
rect 183152 182634 183204 182640
rect 183164 182193 183192 182634
rect 183150 182184 183206 182193
rect 183150 182119 183206 182128
rect 183704 181332 183756 181338
rect 183704 181274 183756 181280
rect 183716 181105 183744 181274
rect 183702 181096 183758 181105
rect 183702 181031 183758 181040
rect 182508 179904 182560 179910
rect 182508 179846 182560 179852
rect 183702 179872 183758 179881
rect 182520 178657 182548 179846
rect 190616 179842 190644 182663
rect 191156 182634 191208 182640
rect 191996 181338 192024 184703
rect 191984 181332 192036 181338
rect 191984 181274 192036 181280
rect 190694 180824 190750 180833
rect 190694 180759 190750 180768
rect 190708 179910 190736 180759
rect 190696 179904 190748 179910
rect 190696 179846 190748 179852
rect 183702 179807 183704 179816
rect 183756 179807 183758 179816
rect 190604 179836 190656 179842
rect 183704 179778 183756 179784
rect 190604 179778 190656 179784
rect 191982 178784 192038 178793
rect 191982 178719 192038 178728
rect 182506 178648 182562 178657
rect 182506 178583 182562 178592
rect 191996 178550 192024 178719
rect 182508 178544 182560 178550
rect 182508 178486 182560 178492
rect 191984 178544 192036 178550
rect 191984 178486 192036 178492
rect 182520 177433 182548 178486
rect 182506 177424 182562 177433
rect 182506 177359 182562 177368
rect 191982 176744 192038 176753
rect 191982 176679 192038 176688
rect 191996 176510 192024 176679
rect 183244 176504 183296 176510
rect 183244 176446 183296 176452
rect 191984 176504 192036 176510
rect 191984 176446 192036 176452
rect 183256 176209 183284 176446
rect 183242 176200 183298 176209
rect 183242 176135 183298 176144
rect 183704 175144 183756 175150
rect 183704 175086 183756 175092
rect 191524 175144 191576 175150
rect 191524 175086 191576 175092
rect 183716 174985 183744 175086
rect 183702 174976 183758 174985
rect 183702 174911 183758 174920
rect 191536 174849 191564 175086
rect 191522 174840 191578 174849
rect 191522 174775 191578 174784
rect 137518 174432 137574 174441
rect 49292 174396 49344 174402
rect 49292 174338 49344 174344
rect 52696 174396 52748 174402
rect 137518 174367 137574 174376
rect 52696 174338 52748 174344
rect 52708 173897 52736 174338
rect 52694 173888 52750 173897
rect 52694 173823 52750 173832
rect 99522 173752 99578 173761
rect 99522 173687 99524 173696
rect 99576 173687 99578 173696
rect 106790 173752 106846 173761
rect 106790 173687 106792 173696
rect 99524 173658 99576 173664
rect 106844 173687 106846 173696
rect 183334 173752 183390 173761
rect 183334 173687 183390 173696
rect 106792 173658 106844 173664
rect 183348 173110 183376 173687
rect 183336 173104 183388 173110
rect 183336 173046 183388 173052
rect 191984 173104 192036 173110
rect 191984 173046 192036 173052
rect 191996 172809 192024 173046
rect 191982 172800 192038 172809
rect 191982 172735 192038 172744
rect 99522 172528 99578 172537
rect 99522 172463 99578 172472
rect 183518 172528 183574 172537
rect 183518 172463 183574 172472
rect 99536 171750 99564 172463
rect 183532 171750 183560 172463
rect 99524 171744 99576 171750
rect 99524 171686 99576 171692
rect 106792 171744 106844 171750
rect 106792 171686 106844 171692
rect 183520 171744 183572 171750
rect 183520 171686 183572 171692
rect 191156 171744 191208 171750
rect 191156 171686 191208 171692
rect 106804 171449 106832 171686
rect 106790 171440 106846 171449
rect 106790 171375 106846 171384
rect 99246 171304 99302 171313
rect 99246 171239 99302 171248
rect 182690 171304 182746 171313
rect 182690 171239 182692 171248
rect 22978 170488 23034 170497
rect 22978 170423 23034 170432
rect 22992 163386 23020 170423
rect 99260 170322 99288 171239
rect 182744 171239 182746 171248
rect 185084 171268 185136 171274
rect 182692 171210 182744 171216
rect 185084 171210 185136 171216
rect 99248 170316 99300 170322
rect 99248 170258 99300 170264
rect 106792 170248 106844 170254
rect 106792 170190 106844 170196
rect 99522 170080 99578 170089
rect 99522 170015 99578 170024
rect 99536 168962 99564 170015
rect 106804 169001 106832 170190
rect 182506 170080 182562 170089
rect 182506 170015 182562 170024
rect 106790 168992 106846 169001
rect 99524 168956 99576 168962
rect 99524 168898 99576 168904
rect 106700 168956 106752 168962
rect 182520 168962 182548 170015
rect 106790 168927 106846 168936
rect 182508 168956 182560 168962
rect 106700 168898 106752 168904
rect 182508 168898 182560 168904
rect 99430 168856 99486 168865
rect 99430 168791 99486 168800
rect 44414 168720 44470 168729
rect 44414 168655 44470 168664
rect 44428 167602 44456 168655
rect 99444 167602 99472 168791
rect 99522 167768 99578 167777
rect 99522 167703 99578 167712
rect 99536 167670 99564 167703
rect 99524 167664 99576 167670
rect 99524 167606 99576 167612
rect 44416 167596 44468 167602
rect 44416 167538 44468 167544
rect 53340 167596 53392 167602
rect 53340 167538 53392 167544
rect 99432 167596 99484 167602
rect 99432 167538 99484 167544
rect 23622 163824 23678 163833
rect 23622 163759 23678 163768
rect 13136 163380 13188 163386
rect 13136 163322 13188 163328
rect 22980 163380 23032 163386
rect 22980 163322 23032 163328
rect 13148 162201 13176 163322
rect 13134 162192 13190 162201
rect 13134 162127 13190 162136
rect 23636 157169 23664 163759
rect 53352 160569 53380 167538
rect 106712 166689 106740 168898
rect 185096 168894 185124 171210
rect 191168 170769 191196 171686
rect 209752 171018 209780 190846
rect 209936 190761 209964 190846
rect 209922 190752 209978 190761
rect 209922 190687 209978 190696
rect 212130 190480 212186 190489
rect 212130 190415 212186 190424
rect 212038 183816 212094 183825
rect 212038 183751 212094 183760
rect 211578 177152 211634 177161
rect 211578 177087 211634 177096
rect 211592 175898 211620 177087
rect 211580 175892 211632 175898
rect 211580 175834 211632 175840
rect 209830 171032 209886 171041
rect 209752 170990 209830 171018
rect 209830 170967 209886 170976
rect 191154 170760 191210 170769
rect 191154 170695 191210 170704
rect 191892 168956 191944 168962
rect 191892 168898 191944 168904
rect 185084 168888 185136 168894
rect 183702 168856 183758 168865
rect 185084 168830 185136 168836
rect 183702 168791 183758 168800
rect 106884 167664 106936 167670
rect 106884 167606 106936 167612
rect 106792 167596 106844 167602
rect 106792 167538 106844 167544
rect 106698 166680 106754 166689
rect 106698 166615 106754 166624
rect 99522 166544 99578 166553
rect 99522 166479 99578 166488
rect 99536 166242 99564 166479
rect 99524 166236 99576 166242
rect 99524 166178 99576 166184
rect 99522 165320 99578 165329
rect 99522 165255 99578 165264
rect 99536 164814 99564 165255
rect 99524 164808 99576 164814
rect 99524 164750 99576 164756
rect 106804 164377 106832 167538
rect 106790 164368 106846 164377
rect 106790 164303 106846 164312
rect 99522 164096 99578 164105
rect 99522 164031 99578 164040
rect 99536 163454 99564 164031
rect 99524 163448 99576 163454
rect 99524 163390 99576 163396
rect 104400 163448 104452 163454
rect 104400 163390 104452 163396
rect 98970 162872 99026 162881
rect 98970 162807 99026 162816
rect 53338 160560 53394 160569
rect 53338 160495 53394 160504
rect 44506 158792 44562 158801
rect 44506 158727 44562 158736
rect 23622 157160 23678 157169
rect 23622 157095 23678 157104
rect 25108 153854 26134 153882
rect 25004 151480 25056 151486
rect 25004 151422 25056 151428
rect 24912 151412 24964 151418
rect 24912 151354 24964 151360
rect 21784 144000 21836 144006
rect 21784 143942 21836 143948
rect 20772 143592 20824 143598
rect 20772 143534 20824 143540
rect 20496 143320 20548 143326
rect 20496 143262 20548 143268
rect 20508 140690 20536 143262
rect 20784 140826 20812 143534
rect 20784 140798 20890 140826
rect 21796 140690 21824 143942
rect 24924 143734 24952 151354
rect 24452 143728 24504 143734
rect 24452 143670 24504 143676
rect 24912 143728 24964 143734
rect 24912 143670 24964 143676
rect 23532 143660 23584 143666
rect 23532 143602 23584 143608
rect 22152 143388 22204 143394
rect 22152 143330 22204 143336
rect 22164 140826 22192 143330
rect 23256 142844 23308 142850
rect 23256 142786 23308 142792
rect 22164 140798 22270 140826
rect 23268 140690 23296 142786
rect 23544 140826 23572 143602
rect 23544 140798 23650 140826
rect 24464 140690 24492 143670
rect 25016 140690 25044 151422
rect 25108 143598 25136 153854
rect 26384 151344 26436 151350
rect 26384 151286 26436 151292
rect 25740 151276 25792 151282
rect 25740 151218 25792 151224
rect 25752 143666 25780 151218
rect 26292 151208 26344 151214
rect 26292 151150 26344 151156
rect 25924 151140 25976 151146
rect 25924 151082 25976 151088
rect 25832 151072 25884 151078
rect 25832 151014 25884 151020
rect 25740 143660 25792 143666
rect 25740 143602 25792 143608
rect 25096 143592 25148 143598
rect 25096 143534 25148 143540
rect 25844 143394 25872 151014
rect 25832 143388 25884 143394
rect 25832 143330 25884 143336
rect 25936 142850 25964 151082
rect 26016 151004 26068 151010
rect 26016 150946 26068 150952
rect 26028 144006 26056 150946
rect 26016 144000 26068 144006
rect 26016 143942 26068 143948
rect 26304 143666 26332 151150
rect 26016 143660 26068 143666
rect 26016 143602 26068 143608
rect 26292 143660 26344 143666
rect 26292 143602 26344 143608
rect 25924 142844 25976 142850
rect 25924 142786 25976 142792
rect 26028 140690 26056 143602
rect 26396 140690 26424 151286
rect 26488 151010 26516 153868
rect 26856 151078 26884 153868
rect 27316 151146 27344 153868
rect 27684 151282 27712 153868
rect 28052 151418 28080 153868
rect 28512 151486 28540 153868
rect 28500 151480 28552 151486
rect 28500 151422 28552 151428
rect 28040 151412 28092 151418
rect 28040 151354 28092 151360
rect 27672 151276 27724 151282
rect 27672 151218 27724 151224
rect 28880 151214 28908 153868
rect 29248 151350 29276 153868
rect 29236 151344 29288 151350
rect 29236 151286 29288 151292
rect 28868 151208 28920 151214
rect 28868 151150 28920 151156
rect 29144 151208 29196 151214
rect 29144 151150 29196 151156
rect 27304 151140 27356 151146
rect 27304 151082 27356 151088
rect 29052 151140 29104 151146
rect 29052 151082 29104 151088
rect 26844 151072 26896 151078
rect 26844 151014 26896 151020
rect 27672 151072 27724 151078
rect 27672 151014 27724 151020
rect 26476 151004 26528 151010
rect 26476 150946 26528 150952
rect 27304 143660 27356 143666
rect 27304 143602 27356 143608
rect 27316 140690 27344 143602
rect 27684 140962 27712 151014
rect 27764 151004 27816 151010
rect 27764 150946 27816 150952
rect 27776 143666 27804 150946
rect 27764 143660 27816 143666
rect 27764 143602 27816 143608
rect 28592 143660 28644 143666
rect 28592 143602 28644 143608
rect 27684 140934 27804 140962
rect 27776 140690 27804 140934
rect 28604 140690 28632 143602
rect 29064 140962 29092 151082
rect 29156 143666 29184 151150
rect 29708 151010 29736 153868
rect 30076 151078 30104 153868
rect 30444 151214 30472 153868
rect 30432 151208 30484 151214
rect 30432 151150 30484 151156
rect 30904 151146 30932 153868
rect 30892 151140 30944 151146
rect 30892 151082 30944 151088
rect 30064 151072 30116 151078
rect 30064 151014 30116 151020
rect 30432 151072 30484 151078
rect 30432 151014 30484 151020
rect 29696 151004 29748 151010
rect 29696 150946 29748 150952
rect 29144 143660 29196 143666
rect 29144 143602 29196 143608
rect 30064 143660 30116 143666
rect 30064 143602 30116 143608
rect 29064 140934 29184 140962
rect 29156 140690 29184 140934
rect 30076 140690 30104 143602
rect 30444 140962 30472 151014
rect 31272 151010 31300 153868
rect 31640 151078 31668 153868
rect 32008 153854 32114 153882
rect 32008 152250 32036 153854
rect 32088 152364 32140 152370
rect 32088 152306 32140 152312
rect 31916 152222 32036 152250
rect 31812 151888 31864 151894
rect 31812 151830 31864 151836
rect 31628 151072 31680 151078
rect 31628 151014 31680 151020
rect 30524 151004 30576 151010
rect 30524 150946 30576 150952
rect 31260 151004 31312 151010
rect 31260 150946 31312 150952
rect 30536 143666 30564 150946
rect 30524 143660 30576 143666
rect 30524 143602 30576 143608
rect 31352 142980 31404 142986
rect 31352 142922 31404 142928
rect 30444 140934 30564 140962
rect 30536 140690 30564 140934
rect 31364 140690 31392 142922
rect 31824 140962 31852 151830
rect 31916 142986 31944 152222
rect 31996 151820 32048 151826
rect 31996 151762 32048 151768
rect 32008 143666 32036 151762
rect 31996 143660 32048 143666
rect 31996 143602 32048 143608
rect 31904 142980 31956 142986
rect 31904 142922 31956 142928
rect 31824 140934 31944 140962
rect 31916 140690 31944 140934
rect 32100 140826 32128 152306
rect 32468 151894 32496 153868
rect 32836 152370 32864 153868
rect 32824 152364 32876 152370
rect 32824 152306 32876 152312
rect 32456 151888 32508 151894
rect 32456 151830 32508 151836
rect 33296 151826 33324 153868
rect 33480 153854 33678 153882
rect 33376 152364 33428 152370
rect 33376 152306 33428 152312
rect 33284 151820 33336 151826
rect 33284 151762 33336 151768
rect 33388 147406 33416 152306
rect 33376 147400 33428 147406
rect 33376 147342 33428 147348
rect 32732 143660 32784 143666
rect 32732 143602 32784 143608
rect 32744 140826 32772 143602
rect 33480 140826 33508 153854
rect 34124 152370 34152 153868
rect 34112 152364 34164 152370
rect 34112 152306 34164 152312
rect 34204 147400 34256 147406
rect 34204 147342 34256 147348
rect 34216 140826 34244 147342
rect 34492 143666 34520 153868
rect 34480 143660 34532 143666
rect 34480 143602 34532 143608
rect 34860 143598 34888 153868
rect 35320 152302 35348 153868
rect 35308 152296 35360 152302
rect 35308 152238 35360 152244
rect 34940 143660 34992 143666
rect 34940 143602 34992 143608
rect 34848 143592 34900 143598
rect 34848 143534 34900 143540
rect 34952 140826 34980 143602
rect 35492 143592 35544 143598
rect 35492 143534 35544 143540
rect 35504 140826 35532 143534
rect 35688 143122 35716 153868
rect 35872 153854 36070 153882
rect 35872 143598 35900 153854
rect 36516 152302 36544 153868
rect 36884 152370 36912 153868
rect 36872 152364 36924 152370
rect 36872 152306 36924 152312
rect 35952 152296 36004 152302
rect 35952 152238 36004 152244
rect 36504 152296 36556 152302
rect 36504 152238 36556 152244
rect 35964 143666 35992 152238
rect 35952 143660 36004 143666
rect 35952 143602 36004 143608
rect 36228 143660 36280 143666
rect 36228 143602 36280 143608
rect 35860 143592 35912 143598
rect 35860 143534 35912 143540
rect 35676 143116 35728 143122
rect 35676 143058 35728 143064
rect 36240 140826 36268 143602
rect 37252 143258 37280 153868
rect 37712 152370 37740 153868
rect 37424 152364 37476 152370
rect 37424 152306 37476 152312
rect 37700 152364 37752 152370
rect 37700 152306 37752 152312
rect 37332 152296 37384 152302
rect 37332 152238 37384 152244
rect 37240 143252 37292 143258
rect 37240 143194 37292 143200
rect 36964 143116 37016 143122
rect 36964 143058 37016 143064
rect 36976 140826 37004 143058
rect 37344 142850 37372 152238
rect 37436 143666 37464 152306
rect 38080 152302 38108 153868
rect 38462 153854 38752 153882
rect 38068 152296 38120 152302
rect 38068 152238 38120 152244
rect 38620 152296 38672 152302
rect 38620 152238 38672 152244
rect 37424 143660 37476 143666
rect 37424 143602 37476 143608
rect 37516 143592 37568 143598
rect 37516 143534 37568 143540
rect 37332 142844 37384 142850
rect 37332 142786 37384 142792
rect 37528 140826 37556 143534
rect 38632 142986 38660 152238
rect 38724 143870 38752 153854
rect 38804 152364 38856 152370
rect 38804 152306 38856 152312
rect 38712 143864 38764 143870
rect 38712 143806 38764 143812
rect 38816 143462 38844 152306
rect 38908 151010 38936 153868
rect 39276 152166 39304 153868
rect 39644 152234 39672 153868
rect 39632 152228 39684 152234
rect 39632 152170 39684 152176
rect 39264 152160 39316 152166
rect 39264 152102 39316 152108
rect 40104 151622 40132 153868
rect 40472 151826 40500 153868
rect 40840 152030 40868 153868
rect 41300 152098 41328 153868
rect 41668 152370 41696 153868
rect 41656 152364 41708 152370
rect 41656 152306 41708 152312
rect 43680 152364 43732 152370
rect 43680 152306 43732 152312
rect 43128 152228 43180 152234
rect 43128 152170 43180 152176
rect 43036 152160 43088 152166
rect 43036 152102 43088 152108
rect 41288 152092 41340 152098
rect 41288 152034 41340 152040
rect 40828 152024 40880 152030
rect 40828 151966 40880 151972
rect 40460 151820 40512 151826
rect 40460 151762 40512 151768
rect 40092 151616 40144 151622
rect 40092 151558 40144 151564
rect 38896 151004 38948 151010
rect 38896 150946 38948 150952
rect 41840 151004 41892 151010
rect 41840 150946 41892 150952
rect 41852 144006 41880 150946
rect 41840 144000 41892 144006
rect 41840 143942 41892 143948
rect 42300 144000 42352 144006
rect 42300 143942 42352 143948
rect 41840 143864 41892 143870
rect 41840 143806 41892 143812
rect 38988 143660 39040 143666
rect 38988 143602 39040 143608
rect 38804 143456 38856 143462
rect 38804 143398 38856 143404
rect 38620 142980 38672 142986
rect 38620 142922 38672 142928
rect 38252 142844 38304 142850
rect 38252 142786 38304 142792
rect 38264 140826 38292 142786
rect 39000 140826 39028 143602
rect 40276 143456 40328 143462
rect 40276 143398 40328 143404
rect 39724 143252 39776 143258
rect 39724 143194 39776 143200
rect 39736 140826 39764 143194
rect 40288 140826 40316 143398
rect 41012 142980 41064 142986
rect 41012 142922 41064 142928
rect 41024 140826 41052 142922
rect 41852 140826 41880 143806
rect 42312 140826 42340 143942
rect 43048 140826 43076 152102
rect 43140 140962 43168 152170
rect 43692 143598 43720 152306
rect 43772 151616 43824 151622
rect 43772 151558 43824 151564
rect 43784 143666 43812 151558
rect 43772 143660 43824 143666
rect 43772 143602 43824 143608
rect 44416 143660 44468 143666
rect 44416 143602 44468 143608
rect 43680 143592 43732 143598
rect 43680 143534 43732 143540
rect 43140 140934 43536 140962
rect 43508 140826 43536 140934
rect 44428 140826 44456 143602
rect 44520 143394 44548 158727
rect 45152 152092 45204 152098
rect 45152 152034 45204 152040
rect 45060 152024 45112 152030
rect 45060 151966 45112 151972
rect 44784 151820 44836 151826
rect 44784 151762 44836 151768
rect 44508 143388 44560 143394
rect 44508 143330 44560 143336
rect 44796 140962 44824 151762
rect 45072 142986 45100 151966
rect 45164 143258 45192 152034
rect 47176 143592 47228 143598
rect 47176 143534 47228 143540
rect 45152 143252 45204 143258
rect 45152 143194 45204 143200
rect 46532 143252 46584 143258
rect 46532 143194 46584 143200
rect 45060 142980 45112 142986
rect 45060 142922 45112 142928
rect 45796 142980 45848 142986
rect 45796 142922 45848 142928
rect 44796 140934 45100 140962
rect 45072 140826 45100 140934
rect 45808 140826 45836 142922
rect 46544 140826 46572 143194
rect 47188 140826 47216 143534
rect 32100 140798 32482 140826
rect 32744 140798 33126 140826
rect 33480 140798 33862 140826
rect 34216 140798 34506 140826
rect 34952 140798 35242 140826
rect 35504 140798 35886 140826
rect 36240 140798 36530 140826
rect 36976 140798 37266 140826
rect 37528 140798 37910 140826
rect 38264 140798 38646 140826
rect 39000 140798 39290 140826
rect 39736 140798 40026 140826
rect 40288 140798 40670 140826
rect 41024 140798 41314 140826
rect 41852 140798 42050 140826
rect 42312 140798 42694 140826
rect 43048 140798 43430 140826
rect 43508 140798 44074 140826
rect 44428 140798 44718 140826
rect 45072 140798 45454 140826
rect 45808 140798 46098 140826
rect 46544 140798 46834 140826
rect 47188 140798 47478 140826
rect 20246 140662 20536 140690
rect 21534 140662 21824 140690
rect 22914 140662 23296 140690
rect 24294 140662 24492 140690
rect 24938 140662 25044 140690
rect 25674 140662 26056 140690
rect 26318 140662 26424 140690
rect 27054 140662 27344 140690
rect 27698 140662 27804 140690
rect 28342 140662 28632 140690
rect 29078 140662 29184 140690
rect 29722 140662 30104 140690
rect 30458 140662 30564 140690
rect 31102 140662 31392 140690
rect 31838 140662 31944 140690
rect 53352 140470 53380 160495
rect 98786 154440 98842 154449
rect 98786 154375 98842 154384
rect 59240 146862 59268 153868
rect 72580 151758 72608 153868
rect 79204 151826 79232 153868
rect 79192 151820 79244 151826
rect 79192 151762 79244 151768
rect 72568 151752 72620 151758
rect 72568 151694 72620 151700
rect 92544 151690 92572 153868
rect 96120 151820 96172 151826
rect 96120 151762 96172 151768
rect 96132 151690 96160 151762
rect 69164 151684 69216 151690
rect 69164 151626 69216 151632
rect 92532 151684 92584 151690
rect 92532 151626 92584 151632
rect 96120 151684 96172 151690
rect 96120 151626 96172 151632
rect 59228 146856 59280 146862
rect 59228 146798 59280 146804
rect 59412 146788 59464 146794
rect 59412 146730 59464 146736
rect 59424 144074 59452 146730
rect 59412 144068 59464 144074
rect 59412 144010 59464 144016
rect 69176 142714 69204 151626
rect 68704 142708 68756 142714
rect 68704 142650 68756 142656
rect 69164 142708 69216 142714
rect 69164 142650 69216 142656
rect 49936 140464 49988 140470
rect 49934 140432 49936 140441
rect 53340 140464 53392 140470
rect 49988 140432 49990 140441
rect 53340 140406 53392 140412
rect 49934 140367 49990 140376
rect 49934 140160 49990 140169
rect 49934 140095 49990 140104
rect 49948 139994 49976 140095
rect 49936 139988 49988 139994
rect 49936 139930 49988 139936
rect 49658 139072 49714 139081
rect 49658 139007 49714 139016
rect 13318 138528 13374 138537
rect 49672 138498 49700 139007
rect 49934 138800 49990 138809
rect 49934 138735 49990 138744
rect 49948 138634 49976 138735
rect 49936 138628 49988 138634
rect 49936 138570 49988 138576
rect 13318 138463 13374 138472
rect 49660 138492 49712 138498
rect 13332 90218 13360 138463
rect 49660 138434 49712 138440
rect 50026 137848 50082 137857
rect 50026 137783 50082 137792
rect 49934 137440 49990 137449
rect 49934 137375 49990 137384
rect 49948 137274 49976 137375
rect 49936 137268 49988 137274
rect 49936 137210 49988 137216
rect 50040 137206 50068 137783
rect 50028 137200 50080 137206
rect 50028 137142 50080 137148
rect 51038 136760 51094 136769
rect 51038 136695 51094 136704
rect 51052 135846 51080 136695
rect 51130 136216 51186 136225
rect 51130 136151 51186 136160
rect 51144 135914 51172 136151
rect 51224 135976 51276 135982
rect 51222 135944 51224 135953
rect 51276 135944 51278 135953
rect 51132 135908 51184 135914
rect 51222 135879 51278 135888
rect 51132 135850 51184 135856
rect 51040 135840 51092 135846
rect 51040 135782 51092 135788
rect 51130 134992 51186 135001
rect 51130 134927 51186 134936
rect 51144 134554 51172 134927
rect 51222 134720 51278 134729
rect 51222 134655 51278 134664
rect 51132 134548 51184 134554
rect 51132 134490 51184 134496
rect 51236 134486 51264 134655
rect 51224 134480 51276 134486
rect 51224 134422 51276 134428
rect 50394 133904 50450 133913
rect 50394 133839 50450 133848
rect 18102 133360 18158 133369
rect 50408 133330 50436 133839
rect 51130 133360 51186 133369
rect 18102 133295 18158 133304
rect 50396 133324 50448 133330
rect 18010 119352 18066 119361
rect 18010 119287 18066 119296
rect 13410 115000 13466 115009
rect 13410 114935 13466 114944
rect 13320 90212 13372 90218
rect 13320 90154 13372 90160
rect 13424 83350 13452 114935
rect 18024 113338 18052 119287
rect 18012 113332 18064 113338
rect 18012 113274 18064 113280
rect 18116 97154 18144 133295
rect 51130 133295 51186 133304
rect 50396 133266 50448 133272
rect 51144 133058 51172 133295
rect 51224 133120 51276 133126
rect 51222 133088 51224 133097
rect 51276 133088 51278 133097
rect 51132 133052 51184 133058
rect 51222 133023 51278 133032
rect 51132 132994 51184 133000
rect 51130 132136 51186 132145
rect 51130 132071 51186 132080
rect 51144 131766 51172 132071
rect 51222 131864 51278 131873
rect 51222 131799 51278 131808
rect 51132 131760 51184 131766
rect 51132 131702 51184 131708
rect 51236 131698 51264 131799
rect 51224 131692 51276 131698
rect 51224 131634 51276 131640
rect 50210 131048 50266 131057
rect 50210 130983 50266 130992
rect 50224 130338 50252 130983
rect 51130 130640 51186 130649
rect 51130 130575 51186 130584
rect 51144 130474 51172 130575
rect 51222 130504 51278 130513
rect 51132 130468 51184 130474
rect 51222 130439 51278 130448
rect 51132 130410 51184 130416
rect 51236 130406 51264 130439
rect 51224 130400 51276 130406
rect 51224 130342 51276 130348
rect 50212 130332 50264 130338
rect 50212 130274 50264 130280
rect 51130 129280 51186 129289
rect 51130 129215 51186 129224
rect 51144 128978 51172 129215
rect 51224 129040 51276 129046
rect 51222 129008 51224 129017
rect 51276 129008 51278 129017
rect 51132 128972 51184 128978
rect 51222 128943 51278 128952
rect 51132 128914 51184 128920
rect 50762 128192 50818 128201
rect 50762 128127 50818 128136
rect 50776 127618 50804 128127
rect 51222 127784 51278 127793
rect 51222 127719 51278 127728
rect 50764 127612 50816 127618
rect 50764 127554 50816 127560
rect 51236 127550 51264 127719
rect 51224 127544 51276 127550
rect 51224 127486 51276 127492
rect 50210 126968 50266 126977
rect 50210 126903 50266 126912
rect 50224 126190 50252 126903
rect 50394 126560 50450 126569
rect 50394 126495 50450 126504
rect 50408 126394 50436 126495
rect 50396 126388 50448 126394
rect 50396 126330 50448 126336
rect 51224 126252 51276 126258
rect 51224 126194 51276 126200
rect 50212 126184 50264 126190
rect 51236 126161 51264 126194
rect 50212 126126 50264 126132
rect 51222 126152 51278 126161
rect 51222 126087 51278 126096
rect 51130 125336 51186 125345
rect 51130 125271 51186 125280
rect 51144 124898 51172 125271
rect 51222 125064 51278 125073
rect 51222 124999 51278 125008
rect 51132 124892 51184 124898
rect 51132 124834 51184 124840
rect 51236 124830 51264 124999
rect 51224 124824 51276 124830
rect 51224 124766 51276 124772
rect 50210 124112 50266 124121
rect 50210 124047 50266 124056
rect 50224 123402 50252 124047
rect 51222 123840 51278 123849
rect 51222 123775 51278 123784
rect 51236 123674 51264 123775
rect 51224 123668 51276 123674
rect 51224 123610 51276 123616
rect 51222 123568 51278 123577
rect 51222 123503 51224 123512
rect 51276 123503 51278 123512
rect 51224 123474 51276 123480
rect 50212 123396 50264 123402
rect 50212 123338 50264 123344
rect 51130 122480 51186 122489
rect 51130 122415 51186 122424
rect 51144 122042 51172 122415
rect 51222 122208 51278 122217
rect 51222 122143 51224 122152
rect 51276 122143 51278 122152
rect 51224 122114 51276 122120
rect 51132 122036 51184 122042
rect 51132 121978 51184 121984
rect 51130 121256 51186 121265
rect 51130 121191 51186 121200
rect 51144 120682 51172 121191
rect 51222 120984 51278 120993
rect 51222 120919 51278 120928
rect 51236 120750 51264 120919
rect 51224 120744 51276 120750
rect 51224 120686 51276 120692
rect 51132 120676 51184 120682
rect 51132 120618 51184 120624
rect 50210 120168 50266 120177
rect 50210 120103 50266 120112
rect 50224 119322 50252 120103
rect 51222 119760 51278 119769
rect 51222 119695 51278 119704
rect 51236 119594 51264 119695
rect 51224 119588 51276 119594
rect 51224 119530 51276 119536
rect 51224 119452 51276 119458
rect 51224 119394 51276 119400
rect 51236 119361 51264 119394
rect 51222 119352 51278 119361
rect 50212 119316 50264 119322
rect 51222 119287 51278 119296
rect 50212 119258 50264 119264
rect 50578 118400 50634 118409
rect 50578 118335 50634 118344
rect 50592 117962 50620 118335
rect 51222 118128 51278 118137
rect 51222 118063 51224 118072
rect 51276 118063 51278 118072
rect 51224 118034 51276 118040
rect 50580 117956 50632 117962
rect 50580 117898 50632 117904
rect 50026 117312 50082 117321
rect 50026 117247 50082 117256
rect 50040 116534 50068 117247
rect 50578 116768 50634 116777
rect 50578 116703 50634 116712
rect 50028 116528 50080 116534
rect 50028 116470 50080 116476
rect 50486 113912 50542 113921
rect 50486 113847 50542 113856
rect 29722 113054 30288 113082
rect 20232 110278 20260 112932
rect 20220 110272 20272 110278
rect 20220 110214 20272 110220
rect 20876 109598 20904 112932
rect 21520 109734 21548 112932
rect 21508 109728 21560 109734
rect 21508 109670 21560 109676
rect 22256 109666 22284 112932
rect 22900 109870 22928 112932
rect 22888 109864 22940 109870
rect 22888 109806 22940 109812
rect 23636 109802 23664 112932
rect 23624 109796 23676 109802
rect 23624 109738 23676 109744
rect 22244 109660 22296 109666
rect 22244 109602 22296 109608
rect 24280 109598 24308 112932
rect 24924 109938 24952 112932
rect 25674 112918 25964 112946
rect 26318 112918 26424 112946
rect 25936 110006 25964 112918
rect 25924 110000 25976 110006
rect 25924 109942 25976 109948
rect 26292 110000 26344 110006
rect 26292 109942 26344 109948
rect 24912 109932 24964 109938
rect 24912 109874 24964 109880
rect 20864 109592 20916 109598
rect 20864 109534 20916 109540
rect 22980 109592 23032 109598
rect 22980 109534 23032 109540
rect 24268 109592 24320 109598
rect 24268 109534 24320 109540
rect 22992 102458 23020 109534
rect 22980 102452 23032 102458
rect 22980 102394 23032 102400
rect 26108 102452 26160 102458
rect 26108 102394 26160 102400
rect 26120 99740 26148 102394
rect 26304 102050 26332 109942
rect 26292 102044 26344 102050
rect 26292 101986 26344 101992
rect 26396 101778 26424 112918
rect 26476 109728 26528 109734
rect 26476 109670 26528 109676
rect 26384 101772 26436 101778
rect 26384 101714 26436 101720
rect 26488 99740 26516 109670
rect 27040 109666 27068 112932
rect 27684 109938 27712 112932
rect 27672 109932 27724 109938
rect 27672 109874 27724 109880
rect 27304 109864 27356 109870
rect 27304 109806 27356 109812
rect 26568 109660 26620 109666
rect 26568 109602 26620 109608
rect 27028 109660 27080 109666
rect 27028 109602 27080 109608
rect 26580 99754 26608 109602
rect 26580 99726 26870 99754
rect 27316 99740 27344 109806
rect 27672 109796 27724 109802
rect 27672 109738 27724 109744
rect 27684 99740 27712 109738
rect 28328 109598 28356 112932
rect 29064 110006 29092 112932
rect 29052 110000 29104 110006
rect 29052 109942 29104 109948
rect 30064 109932 30116 109938
rect 30064 109874 30116 109880
rect 28500 109864 28552 109870
rect 28500 109806 28552 109812
rect 28132 109592 28184 109598
rect 28132 109534 28184 109540
rect 28316 109592 28368 109598
rect 28316 109534 28368 109540
rect 28144 99754 28172 109534
rect 28066 99726 28172 99754
rect 28512 99740 28540 109806
rect 29696 109660 29748 109666
rect 29696 109602 29748 109608
rect 29144 109592 29196 109598
rect 29144 109534 29196 109540
rect 29156 102050 29184 109534
rect 28868 102044 28920 102050
rect 28868 101986 28920 101992
rect 29144 102044 29196 102050
rect 29144 101986 29196 101992
rect 28880 99740 28908 101986
rect 29236 101772 29288 101778
rect 29236 101714 29288 101720
rect 29248 99740 29276 101714
rect 29708 99740 29736 109602
rect 30076 99740 30104 109874
rect 30260 102662 30288 113054
rect 32560 113054 33126 113082
rect 33940 113054 34506 113082
rect 36608 113054 37266 113082
rect 38080 113054 38646 113082
rect 40840 113054 41314 113082
rect 43600 113054 44074 113082
rect 44888 113054 45454 113082
rect 30458 112918 30564 112946
rect 30248 102656 30300 102662
rect 30248 102598 30300 102604
rect 30432 102044 30484 102050
rect 30432 101986 30484 101992
rect 30444 99740 30472 101986
rect 30536 101846 30564 112918
rect 30892 110000 30944 110006
rect 30892 109942 30944 109948
rect 30524 101840 30576 101846
rect 30524 101782 30576 101788
rect 30904 99740 30932 109942
rect 31088 109598 31116 112932
rect 31838 112918 31944 112946
rect 31076 109592 31128 109598
rect 31076 109534 31128 109540
rect 31812 109592 31864 109598
rect 31812 109534 31864 109540
rect 31260 102656 31312 102662
rect 31260 102598 31312 102604
rect 31272 99740 31300 102598
rect 31628 101840 31680 101846
rect 31628 101782 31680 101788
rect 31640 99740 31668 101782
rect 31824 101386 31852 109534
rect 31916 101522 31944 112918
rect 32008 112918 32482 112946
rect 32008 102662 32036 112918
rect 32560 112674 32588 113054
rect 32100 112646 32588 112674
rect 33388 112918 33862 112946
rect 31996 102656 32048 102662
rect 31996 102598 32048 102604
rect 32100 102594 32128 112646
rect 32824 102656 32876 102662
rect 32824 102598 32876 102604
rect 32088 102588 32140 102594
rect 32088 102530 32140 102536
rect 31916 101494 32128 101522
rect 32100 101386 32128 101494
rect 31824 101358 32036 101386
rect 32100 101358 32220 101386
rect 32008 99754 32036 101358
rect 32192 99754 32220 101358
rect 32008 99726 32114 99754
rect 32192 99726 32482 99754
rect 32836 99740 32864 102598
rect 33284 102588 33336 102594
rect 33284 102530 33336 102536
rect 33296 99740 33324 102530
rect 33388 99754 33416 112918
rect 33940 112674 33968 113054
rect 33480 112646 33968 112674
rect 34860 112918 35242 112946
rect 35504 112918 35886 112946
rect 36148 112918 36530 112946
rect 33480 102662 33508 112646
rect 33468 102656 33520 102662
rect 33468 102598 33520 102604
rect 34112 102656 34164 102662
rect 34112 102598 34164 102604
rect 33388 99726 33678 99754
rect 34124 99740 34152 102598
rect 34860 101250 34888 112918
rect 35504 102662 35532 112918
rect 35124 102656 35176 102662
rect 35124 102598 35176 102604
rect 35492 102656 35544 102662
rect 35492 102598 35544 102604
rect 35676 102656 35728 102662
rect 35676 102598 35728 102604
rect 34676 101222 34888 101250
rect 34676 99754 34704 101222
rect 35136 99754 35164 102598
rect 35308 101704 35360 101710
rect 35308 101646 35360 101652
rect 34506 99726 34704 99754
rect 34874 99726 35164 99754
rect 35320 99740 35348 101646
rect 35688 99740 35716 102598
rect 36148 101710 36176 112918
rect 36608 102662 36636 113054
rect 37528 112918 37910 112946
rect 36596 102656 36648 102662
rect 36596 102598 36648 102604
rect 36504 102588 36556 102594
rect 36504 102530 36556 102536
rect 36136 101704 36188 101710
rect 36136 101646 36188 101652
rect 36044 101636 36096 101642
rect 36044 101578 36096 101584
rect 36056 99740 36084 101578
rect 36516 99740 36544 102530
rect 36872 102452 36924 102458
rect 36872 102394 36924 102400
rect 36884 99740 36912 102394
rect 37240 102044 37292 102050
rect 37240 101986 37292 101992
rect 37252 99740 37280 101986
rect 37528 101642 37556 112918
rect 37700 102656 37752 102662
rect 37700 102598 37752 102604
rect 37516 101636 37568 101642
rect 37516 101578 37568 101584
rect 37712 99740 37740 102598
rect 38080 102594 38108 113054
rect 38252 109660 38304 109666
rect 38252 109602 38304 109608
rect 38160 109592 38212 109598
rect 38160 109534 38212 109540
rect 38068 102588 38120 102594
rect 38068 102530 38120 102536
rect 38172 102458 38200 109534
rect 38160 102452 38212 102458
rect 38160 102394 38212 102400
rect 38068 102384 38120 102390
rect 38068 102326 38120 102332
rect 38080 99740 38108 102326
rect 38264 102050 38292 109602
rect 39276 109598 39304 112932
rect 40012 109666 40040 112932
rect 40288 112918 40670 112946
rect 40000 109660 40052 109666
rect 40000 109602 40052 109608
rect 39264 109592 39316 109598
rect 39264 109534 39316 109540
rect 40288 102662 40316 112918
rect 40276 102656 40328 102662
rect 40276 102598 40328 102604
rect 40840 102390 40868 113054
rect 41852 112918 42050 112946
rect 42312 112918 42694 112946
rect 43048 112918 43430 112946
rect 41748 110272 41800 110278
rect 41748 110214 41800 110220
rect 40828 102384 40880 102390
rect 40828 102326 40880 102332
rect 38252 102044 38304 102050
rect 38252 101986 38304 101992
rect 41656 102044 41708 102050
rect 41656 101986 41708 101992
rect 40092 101908 40144 101914
rect 40092 101850 40144 101856
rect 39632 101772 39684 101778
rect 39632 101714 39684 101720
rect 39264 101704 39316 101710
rect 39264 101646 39316 101652
rect 38436 101636 38488 101642
rect 38436 101578 38488 101584
rect 38448 99740 38476 101578
rect 38896 101500 38948 101506
rect 38896 101442 38948 101448
rect 38908 99740 38936 101442
rect 39276 99740 39304 101646
rect 39644 99740 39672 101714
rect 40104 99740 40132 101850
rect 40828 101840 40880 101846
rect 40828 101782 40880 101788
rect 40460 101568 40512 101574
rect 40460 101510 40512 101516
rect 40472 99740 40500 101510
rect 40840 99740 40868 101782
rect 41288 101432 41340 101438
rect 41288 101374 41340 101380
rect 41300 99740 41328 101374
rect 41668 99740 41696 101986
rect 18104 97148 18156 97154
rect 18104 97090 18156 97096
rect 22336 97148 22388 97154
rect 22336 97090 22388 97096
rect 22348 96513 22376 97090
rect 22334 96504 22390 96513
rect 22334 96439 22390 96448
rect 41760 95266 41788 110214
rect 41852 101642 41880 112918
rect 41840 101636 41892 101642
rect 41840 101578 41892 101584
rect 42312 101506 42340 112918
rect 42944 109728 42996 109734
rect 42944 109670 42996 109676
rect 42956 102050 42984 109670
rect 42944 102044 42996 102050
rect 42944 101986 42996 101992
rect 43048 101710 43076 112918
rect 43600 101778 43628 113054
rect 44428 112918 44718 112946
rect 44428 101914 44456 112918
rect 44416 101908 44468 101914
rect 44416 101850 44468 101856
rect 43588 101772 43640 101778
rect 43588 101714 43640 101720
rect 43036 101704 43088 101710
rect 43036 101646 43088 101652
rect 44888 101574 44916 113054
rect 45060 109660 45112 109666
rect 45060 109602 45112 109608
rect 44876 101568 44928 101574
rect 44876 101510 44928 101516
rect 42300 101500 42352 101506
rect 42300 101442 42352 101448
rect 45072 101438 45100 109602
rect 46084 109598 46112 112932
rect 46820 109666 46848 112932
rect 47464 109734 47492 112932
rect 47452 109728 47504 109734
rect 47452 109670 47504 109676
rect 46808 109660 46860 109666
rect 46808 109602 46860 109608
rect 45152 109592 45204 109598
rect 45152 109534 45204 109540
rect 46072 109592 46124 109598
rect 46072 109534 46124 109540
rect 45164 101846 45192 109534
rect 50500 101982 50528 113847
rect 50592 102050 50620 116703
rect 50762 116496 50818 116505
rect 50762 116431 50818 116440
rect 50670 115544 50726 115553
rect 50670 115479 50726 115488
rect 50684 102186 50712 115479
rect 50672 102180 50724 102186
rect 50672 102122 50724 102128
rect 50776 102118 50804 116431
rect 50854 115136 50910 115145
rect 50854 115071 50910 115080
rect 50868 102254 50896 115071
rect 51130 114456 51186 114465
rect 51130 114391 51186 114400
rect 50946 113776 51002 113785
rect 50946 113711 51002 113720
rect 50960 102458 50988 113711
rect 50948 102452 51000 102458
rect 50948 102394 51000 102400
rect 51144 102390 51172 114391
rect 51222 112824 51278 112833
rect 51222 112759 51224 112768
rect 51276 112759 51278 112768
rect 51224 112730 51276 112736
rect 53352 110278 53380 140406
rect 58492 139988 58544 139994
rect 58492 139930 58544 139936
rect 58504 138945 58532 139930
rect 58490 138936 58546 138945
rect 58490 138871 58546 138880
rect 68716 138786 68744 142650
rect 68408 138758 68744 138786
rect 58400 138628 58452 138634
rect 58400 138570 58452 138576
rect 58308 137268 58360 137274
rect 58308 137210 58360 137216
rect 58216 137200 58268 137206
rect 58216 137142 58268 137148
rect 58228 136633 58256 137142
rect 58214 136624 58270 136633
rect 58214 136559 58270 136568
rect 58320 136089 58348 137210
rect 58412 137177 58440 138570
rect 92716 138560 92768 138566
rect 92714 138528 92716 138537
rect 92768 138528 92770 138537
rect 58952 138492 59004 138498
rect 92714 138463 92770 138472
rect 92808 138492 92860 138498
rect 58952 138434 59004 138440
rect 92808 138434 92860 138440
rect 58964 138265 58992 138434
rect 58950 138256 59006 138265
rect 58950 138191 59006 138200
rect 92820 138129 92848 138434
rect 92806 138120 92862 138129
rect 92806 138055 92862 138064
rect 58398 137168 58454 137177
rect 58398 137103 58454 137112
rect 92714 137168 92770 137177
rect 92714 137103 92716 137112
rect 92768 137103 92770 137112
rect 92716 137074 92768 137080
rect 92808 137064 92860 137070
rect 92808 137006 92860 137012
rect 92716 136996 92768 137002
rect 92716 136938 92768 136944
rect 92728 136497 92756 136938
rect 92820 136905 92848 137006
rect 92806 136896 92862 136905
rect 92806 136831 92862 136840
rect 92714 136488 92770 136497
rect 92714 136423 92770 136432
rect 58306 136080 58362 136089
rect 58306 136015 58362 136024
rect 56652 135976 56704 135982
rect 56652 135918 56704 135924
rect 56560 135840 56612 135846
rect 56560 135782 56612 135788
rect 56572 135642 56600 135782
rect 56560 135636 56612 135642
rect 56560 135578 56612 135584
rect 56100 134480 56152 134486
rect 56100 134422 56152 134428
rect 56112 133738 56140 134422
rect 56664 134282 56692 135918
rect 56744 135908 56796 135914
rect 56744 135850 56796 135856
rect 56756 135370 56784 135850
rect 92808 135772 92860 135778
rect 92808 135714 92860 135720
rect 92716 135704 92768 135710
rect 92716 135646 92768 135652
rect 58216 135636 58268 135642
rect 58216 135578 58268 135584
rect 58228 135409 58256 135578
rect 92728 135545 92756 135646
rect 92714 135536 92770 135545
rect 92714 135471 92770 135480
rect 58214 135400 58270 135409
rect 56744 135364 56796 135370
rect 58214 135335 58270 135344
rect 58308 135364 58360 135370
rect 56744 135306 56796 135312
rect 58308 135306 58360 135312
rect 58320 134865 58348 135306
rect 92820 135273 92848 135714
rect 92806 135264 92862 135273
rect 92806 135199 92862 135208
rect 58306 134856 58362 134865
rect 58306 134791 58362 134800
rect 59412 134548 59464 134554
rect 59412 134490 59464 134496
rect 58216 134412 58268 134418
rect 58216 134354 58268 134360
rect 56652 134276 56704 134282
rect 56652 134218 56704 134224
rect 56100 133732 56152 133738
rect 56100 133674 56152 133680
rect 58228 133641 58256 134354
rect 58400 134276 58452 134282
rect 58400 134218 58452 134224
rect 58412 134185 58440 134218
rect 58398 134176 58454 134185
rect 58398 134111 58454 134120
rect 58308 133732 58360 133738
rect 58308 133674 58360 133680
rect 58214 133632 58270 133641
rect 58214 133567 58270 133576
rect 56744 133324 56796 133330
rect 56744 133266 56796 133272
rect 55548 133120 55600 133126
rect 55548 133062 55600 133068
rect 55456 131760 55508 131766
rect 55456 131702 55508 131708
rect 55468 131154 55496 131702
rect 55560 131426 55588 133062
rect 56756 132922 56784 133266
rect 58320 133097 58348 133674
rect 58306 133088 58362 133097
rect 58306 133023 58362 133032
rect 59424 132990 59452 134490
rect 92900 134412 92952 134418
rect 92900 134354 92952 134360
rect 92808 134344 92860 134350
rect 92808 134286 92860 134292
rect 92716 134276 92768 134282
rect 92716 134218 92768 134224
rect 92728 134185 92756 134218
rect 92714 134176 92770 134185
rect 92714 134111 92770 134120
rect 92820 134049 92848 134286
rect 92806 134040 92862 134049
rect 92806 133975 92862 133984
rect 92912 133505 92940 134354
rect 92898 133496 92954 133505
rect 92898 133431 92954 133440
rect 58216 132984 58268 132990
rect 58216 132926 58268 132932
rect 59412 132984 59464 132990
rect 59412 132926 59464 132932
rect 92808 132984 92860 132990
rect 92808 132926 92860 132932
rect 56744 132916 56796 132922
rect 56744 132858 56796 132864
rect 58228 131873 58256 132926
rect 58308 132916 58360 132922
rect 58308 132858 58360 132864
rect 92716 132916 92768 132922
rect 92716 132858 92768 132864
rect 58320 132417 58348 132858
rect 92728 132689 92756 132858
rect 92714 132680 92770 132689
rect 92714 132615 92770 132624
rect 58306 132408 58362 132417
rect 58306 132343 58362 132352
rect 92820 132281 92848 132926
rect 92806 132272 92862 132281
rect 92806 132207 92862 132216
rect 58214 131864 58270 131873
rect 58214 131799 58270 131808
rect 58492 131692 58544 131698
rect 58492 131634 58544 131640
rect 55548 131420 55600 131426
rect 55548 131362 55600 131368
rect 58216 131420 58268 131426
rect 58216 131362 58268 131368
rect 58228 131193 58256 131362
rect 58214 131184 58270 131193
rect 55456 131148 55508 131154
rect 58214 131119 58270 131128
rect 58308 131148 58360 131154
rect 55456 131090 55508 131096
rect 58308 131090 58360 131096
rect 58320 130649 58348 131090
rect 58306 130640 58362 130649
rect 58306 130575 58362 130584
rect 56744 130468 56796 130474
rect 56744 130410 56796 130416
rect 56560 130400 56612 130406
rect 56560 130342 56612 130348
rect 56376 128972 56428 128978
rect 56376 128914 56428 128920
rect 56388 128570 56416 128914
rect 56572 128774 56600 130342
rect 56652 129040 56704 129046
rect 56652 128982 56704 128988
rect 56560 128768 56612 128774
rect 56560 128710 56612 128716
rect 56376 128564 56428 128570
rect 56376 128506 56428 128512
rect 56664 127482 56692 128982
rect 56756 128842 56784 130410
rect 58216 130196 58268 130202
rect 58216 130138 58268 130144
rect 58228 129425 58256 130138
rect 58504 130105 58532 131634
rect 92808 131624 92860 131630
rect 92808 131566 92860 131572
rect 92716 131556 92768 131562
rect 92716 131498 92768 131504
rect 92728 131329 92756 131498
rect 92714 131320 92770 131329
rect 92714 131255 92770 131264
rect 92820 131057 92848 131566
rect 92806 131048 92862 131057
rect 92806 130983 92862 130992
rect 92808 130264 92860 130270
rect 92808 130206 92860 130212
rect 92716 130196 92768 130202
rect 92716 130138 92768 130144
rect 92728 130105 92756 130138
rect 58490 130096 58546 130105
rect 58490 130031 58546 130040
rect 92714 130096 92770 130105
rect 92714 130031 92770 130040
rect 92820 129833 92848 130206
rect 92806 129824 92862 129833
rect 92806 129759 92862 129768
rect 58214 129416 58270 129425
rect 58214 129351 58270 129360
rect 92900 128904 92952 128910
rect 58214 128872 58270 128881
rect 56744 128836 56796 128842
rect 58214 128807 58216 128816
rect 56744 128778 56796 128784
rect 58268 128807 58270 128816
rect 92714 128872 92770 128881
rect 92900 128846 92952 128852
rect 92714 128807 92770 128816
rect 92808 128836 92860 128842
rect 58216 128778 58268 128784
rect 92728 128774 92756 128807
rect 92808 128778 92860 128784
rect 58400 128768 58452 128774
rect 58400 128710 58452 128716
rect 92716 128768 92768 128774
rect 92716 128710 92768 128716
rect 58308 128564 58360 128570
rect 58308 128506 58360 128512
rect 58320 127657 58348 128506
rect 58412 128201 58440 128710
rect 92820 128473 92848 128778
rect 92806 128464 92862 128473
rect 92806 128399 92862 128408
rect 58398 128192 58454 128201
rect 58398 128127 58454 128136
rect 92912 128065 92940 128846
rect 92898 128056 92954 128065
rect 92898 127991 92954 128000
rect 58306 127648 58362 127657
rect 58216 127612 58268 127618
rect 58306 127583 58362 127592
rect 58216 127554 58268 127560
rect 56652 127476 56704 127482
rect 56652 127418 56704 127424
rect 58228 126433 58256 127554
rect 58308 127544 58360 127550
rect 58308 127486 58360 127492
rect 58214 126424 58270 126433
rect 56744 126388 56796 126394
rect 58214 126359 58270 126368
rect 56744 126330 56796 126336
rect 56100 126252 56152 126258
rect 56100 126194 56152 126200
rect 55456 124892 55508 124898
rect 55456 124834 55508 124840
rect 55468 124762 55496 124834
rect 55456 124756 55508 124762
rect 55456 124698 55508 124704
rect 56112 124626 56140 126194
rect 56756 124694 56784 126330
rect 58216 126184 58268 126190
rect 58216 126126 58268 126132
rect 58228 125209 58256 126126
rect 58320 125889 58348 127486
rect 58400 127476 58452 127482
rect 58400 127418 58452 127424
rect 92808 127476 92860 127482
rect 92808 127418 92860 127424
rect 58412 127113 58440 127418
rect 92716 127408 92768 127414
rect 92716 127350 92768 127356
rect 92728 127249 92756 127350
rect 92714 127240 92770 127249
rect 92714 127175 92770 127184
rect 58398 127104 58454 127113
rect 58398 127039 58454 127048
rect 92820 126977 92848 127418
rect 92806 126968 92862 126977
rect 92806 126903 92862 126912
rect 92716 126116 92768 126122
rect 92716 126058 92768 126064
rect 92728 126025 92756 126058
rect 92808 126048 92860 126054
rect 92714 126016 92770 126025
rect 92808 125990 92860 125996
rect 92714 125951 92770 125960
rect 58306 125880 58362 125889
rect 58306 125815 58362 125824
rect 92820 125617 92848 125990
rect 92806 125608 92862 125617
rect 92806 125543 92862 125552
rect 58214 125200 58270 125209
rect 58214 125135 58270 125144
rect 58400 124824 58452 124830
rect 58400 124766 58452 124772
rect 58216 124756 58268 124762
rect 58216 124698 58268 124704
rect 56744 124688 56796 124694
rect 56744 124630 56796 124636
rect 56100 124620 56152 124626
rect 56100 124562 56152 124568
rect 55548 123668 55600 123674
rect 55548 123610 55600 123616
rect 55456 123532 55508 123538
rect 55456 123474 55508 123480
rect 55468 121566 55496 123474
rect 55560 121838 55588 123610
rect 58228 123441 58256 124698
rect 58308 124688 58360 124694
rect 58306 124656 58308 124665
rect 58360 124656 58362 124665
rect 58306 124591 58362 124600
rect 58214 123432 58270 123441
rect 58214 123367 58270 123376
rect 58216 123260 58268 123266
rect 58216 123202 58268 123208
rect 58228 122217 58256 123202
rect 58412 122897 58440 124766
rect 92900 124756 92952 124762
rect 92900 124698 92952 124704
rect 92716 124688 92768 124694
rect 92714 124656 92716 124665
rect 92768 124656 92770 124665
rect 58492 124620 58544 124626
rect 92714 124591 92770 124600
rect 92808 124620 92860 124626
rect 58492 124562 58544 124568
rect 92808 124562 92860 124568
rect 58504 124121 58532 124562
rect 92820 124393 92848 124562
rect 92806 124384 92862 124393
rect 92806 124319 92862 124328
rect 58490 124112 58546 124121
rect 58490 124047 58546 124056
rect 92912 123985 92940 124698
rect 92898 123976 92954 123985
rect 92898 123911 92954 123920
rect 92808 123328 92860 123334
rect 92808 123270 92860 123276
rect 92716 123260 92768 123266
rect 92716 123202 92768 123208
rect 92728 123033 92756 123202
rect 92714 123024 92770 123033
rect 92714 122959 92770 122968
rect 58398 122888 58454 122897
rect 58398 122823 58454 122832
rect 92820 122761 92848 123270
rect 92806 122752 92862 122761
rect 92806 122687 92862 122696
rect 58214 122208 58270 122217
rect 55732 122172 55784 122178
rect 58214 122143 58270 122152
rect 55732 122114 55784 122120
rect 55640 122036 55692 122042
rect 55640 121978 55692 121984
rect 55548 121832 55600 121838
rect 55548 121774 55600 121780
rect 55456 121560 55508 121566
rect 55456 121502 55508 121508
rect 55652 120614 55680 121978
rect 55640 120608 55692 120614
rect 55640 120550 55692 120556
rect 55744 120546 55772 122114
rect 92808 121968 92860 121974
rect 92808 121910 92860 121916
rect 92716 121900 92768 121906
rect 92716 121842 92768 121848
rect 58216 121832 58268 121838
rect 92728 121809 92756 121842
rect 58216 121774 58268 121780
rect 92714 121800 92770 121809
rect 58228 121673 58256 121774
rect 92714 121735 92770 121744
rect 58214 121664 58270 121673
rect 58214 121599 58270 121608
rect 58216 121560 58268 121566
rect 92820 121537 92848 121910
rect 58216 121502 58268 121508
rect 92806 121528 92862 121537
rect 58228 121129 58256 121502
rect 92806 121463 92862 121472
rect 58214 121120 58270 121129
rect 58214 121055 58270 121064
rect 58492 120744 58544 120750
rect 58492 120686 58544 120692
rect 58308 120676 58360 120682
rect 58308 120618 58360 120624
rect 58216 120608 58268 120614
rect 58216 120550 58268 120556
rect 55732 120540 55784 120546
rect 55732 120482 55784 120488
rect 58228 120449 58256 120550
rect 58214 120440 58270 120449
rect 58214 120375 58270 120384
rect 56744 119588 56796 119594
rect 56744 119530 56796 119536
rect 56284 119452 56336 119458
rect 56284 119394 56336 119400
rect 55548 117956 55600 117962
rect 55548 117898 55600 117904
rect 55560 116466 55588 117898
rect 56296 117758 56324 119394
rect 56560 118092 56612 118098
rect 56560 118034 56612 118040
rect 56284 117752 56336 117758
rect 56284 117694 56336 117700
rect 55548 116460 55600 116466
rect 55548 116402 55600 116408
rect 56572 116398 56600 118034
rect 56756 117826 56784 119530
rect 58320 119225 58348 120618
rect 58400 120540 58452 120546
rect 58400 120482 58452 120488
rect 58412 119905 58440 120482
rect 58398 119896 58454 119905
rect 58398 119831 58454 119840
rect 58306 119216 58362 119225
rect 58216 119180 58268 119186
rect 58306 119151 58362 119160
rect 58216 119122 58268 119128
rect 58228 118137 58256 119122
rect 58504 118681 58532 120686
rect 92808 120608 92860 120614
rect 92808 120550 92860 120556
rect 92716 120540 92768 120546
rect 92716 120482 92768 120488
rect 92728 120449 92756 120482
rect 92714 120440 92770 120449
rect 92714 120375 92770 120384
rect 92820 120041 92848 120550
rect 92806 120032 92862 120041
rect 92806 119967 92862 119976
rect 92900 119248 92952 119254
rect 92714 119216 92770 119225
rect 92900 119190 92952 119196
rect 92714 119151 92770 119160
rect 92808 119180 92860 119186
rect 92728 119118 92756 119151
rect 92808 119122 92860 119128
rect 92716 119112 92768 119118
rect 92716 119054 92768 119060
rect 92820 118953 92848 119122
rect 92806 118944 92862 118953
rect 92806 118879 92862 118888
rect 58490 118672 58546 118681
rect 58490 118607 58546 118616
rect 92912 118545 92940 119190
rect 92898 118536 92954 118545
rect 92898 118471 92954 118480
rect 58214 118128 58270 118137
rect 58214 118063 58270 118072
rect 56744 117820 56796 117826
rect 56744 117762 56796 117768
rect 58216 117820 58268 117826
rect 58216 117762 58268 117768
rect 92808 117820 92860 117826
rect 92808 117762 92860 117768
rect 58228 117457 58256 117762
rect 58308 117752 58360 117758
rect 58308 117694 58360 117700
rect 92716 117752 92768 117758
rect 92716 117694 92768 117700
rect 58214 117448 58270 117457
rect 58214 117383 58270 117392
rect 58320 116913 58348 117694
rect 92728 117593 92756 117694
rect 92714 117584 92770 117593
rect 92714 117519 92770 117528
rect 92820 117185 92848 117762
rect 92806 117176 92862 117185
rect 92806 117111 92862 117120
rect 58306 116904 58362 116913
rect 58306 116839 58362 116848
rect 94004 116596 94056 116602
rect 94004 116538 94056 116544
rect 58216 116528 58268 116534
rect 58216 116470 58268 116476
rect 92624 116528 92676 116534
rect 92624 116470 92676 116476
rect 56560 116392 56612 116398
rect 56560 116334 56612 116340
rect 58228 115145 58256 116470
rect 58308 116460 58360 116466
rect 58308 116402 58360 116408
rect 58320 116233 58348 116402
rect 58400 116392 58452 116398
rect 58400 116334 58452 116340
rect 58306 116224 58362 116233
rect 58306 116159 58362 116168
rect 58412 115689 58440 116334
rect 58398 115680 58454 115689
rect 58398 115615 58454 115624
rect 91244 115236 91296 115242
rect 91244 115178 91296 115184
rect 59320 115168 59372 115174
rect 58214 115136 58270 115145
rect 59320 115110 59372 115116
rect 90600 115168 90652 115174
rect 90600 115110 90652 115116
rect 58214 115071 58270 115080
rect 54720 112788 54772 112794
rect 54720 112730 54772 112736
rect 53340 110272 53392 110278
rect 53340 110214 53392 110220
rect 51132 102384 51184 102390
rect 51132 102326 51184 102332
rect 50856 102248 50908 102254
rect 50856 102190 50908 102196
rect 50764 102112 50816 102118
rect 50764 102054 50816 102060
rect 50580 102044 50632 102050
rect 50580 101986 50632 101992
rect 50488 101976 50540 101982
rect 50488 101918 50540 101924
rect 45152 101840 45204 101846
rect 45152 101782 45204 101788
rect 45060 101432 45112 101438
rect 45060 101374 45112 101380
rect 41838 95280 41894 95289
rect 41760 95238 41838 95266
rect 41838 95215 41894 95224
rect 13502 91336 13558 91345
rect 13502 91271 13558 91280
rect 13412 83344 13464 83350
rect 13412 83286 13464 83292
rect 13516 77842 13544 91271
rect 22336 90212 22388 90218
rect 22336 90154 22388 90160
rect 22348 89849 22376 90154
rect 22334 89840 22390 89849
rect 22334 89775 22390 89784
rect 44414 84808 44470 84817
rect 44414 84743 44416 84752
rect 44468 84743 44470 84752
rect 52696 84772 52748 84778
rect 44416 84714 44468 84720
rect 52696 84714 52748 84720
rect 22336 83344 22388 83350
rect 22336 83286 22388 83292
rect 22348 83185 22376 83286
rect 22334 83176 22390 83185
rect 22334 83111 22390 83120
rect 52708 79921 52736 84714
rect 52694 79912 52750 79921
rect 52694 79847 52750 79856
rect 13504 77836 13556 77842
rect 13504 77778 13556 77784
rect 22336 77836 22388 77842
rect 22336 77778 22388 77784
rect 22348 76521 22376 77778
rect 22334 76512 22390 76521
rect 22334 76447 22390 76456
rect 44414 74744 44470 74753
rect 44414 74679 44470 74688
rect 44428 74374 44456 74679
rect 53352 74374 53380 110214
rect 54732 102662 54760 112730
rect 59332 108238 59360 115110
rect 61448 114822 61600 114850
rect 62980 114822 63316 114850
rect 61448 110958 61476 114822
rect 61436 110952 61488 110958
rect 61436 110894 61488 110900
rect 61448 110278 61476 110894
rect 63288 110890 63316 114822
rect 64116 114822 64452 114850
rect 65312 114822 65832 114850
rect 66508 114822 67304 114850
rect 67888 114822 68684 114850
rect 69268 114822 70156 114850
rect 70648 114822 71536 114850
rect 72028 114822 73008 114850
rect 73500 114822 74388 114850
rect 75524 114822 75860 114850
rect 76904 114822 77240 114850
rect 77548 114822 78712 114850
rect 79756 114822 80092 114850
rect 81228 114822 81564 114850
rect 82608 114822 82944 114850
rect 84080 114822 84416 114850
rect 85460 114822 85796 114850
rect 87208 114822 87268 114850
rect 90120 114822 90456 114850
rect 64116 113338 64144 114822
rect 64104 113332 64156 113338
rect 64104 113274 64156 113280
rect 63276 110884 63328 110890
rect 63276 110826 63328 110832
rect 61436 110272 61488 110278
rect 61436 110214 61488 110220
rect 59320 108232 59372 108238
rect 59320 108174 59372 108180
rect 59412 108164 59464 108170
rect 59412 108106 59464 108112
rect 54720 102656 54772 102662
rect 54720 102598 54772 102604
rect 56468 102656 56520 102662
rect 56468 102598 56520 102604
rect 56480 99740 56508 102598
rect 57572 102452 57624 102458
rect 57572 102394 57624 102400
rect 57584 99740 57612 102394
rect 59424 101982 59452 108106
rect 59780 102384 59832 102390
rect 59780 102326 59832 102332
rect 58676 101976 58728 101982
rect 58676 101918 58728 101924
rect 59412 101976 59464 101982
rect 59412 101918 59464 101924
rect 58688 99740 58716 101918
rect 59792 99740 59820 102326
rect 60884 102248 60936 102254
rect 60884 102190 60936 102196
rect 60896 99740 60924 102190
rect 61988 102180 62040 102186
rect 61988 102122 62040 102128
rect 62000 99740 62028 102122
rect 63092 102112 63144 102118
rect 63092 102054 63144 102060
rect 63104 99740 63132 102054
rect 64196 102044 64248 102050
rect 64196 101986 64248 101992
rect 64208 99740 64236 101986
rect 65312 99740 65340 114822
rect 66508 101386 66536 114822
rect 67888 101386 67916 114822
rect 66416 101358 66536 101386
rect 67704 101358 67916 101386
rect 69268 101370 69296 114822
rect 70648 101370 70676 114822
rect 72028 101370 72056 114822
rect 73500 101438 73528 114822
rect 75524 111094 75552 114822
rect 74040 111088 74092 111094
rect 74040 111030 74092 111036
rect 75512 111088 75564 111094
rect 75512 111030 75564 111036
rect 72384 101432 72436 101438
rect 72384 101374 72436 101380
rect 73488 101432 73540 101438
rect 73488 101374 73540 101380
rect 68612 101364 68664 101370
rect 66416 99740 66444 101358
rect 67704 99754 67732 101358
rect 68612 101306 68664 101312
rect 69256 101364 69308 101370
rect 69256 101306 69308 101312
rect 69808 101364 69860 101370
rect 69808 101306 69860 101312
rect 70636 101364 70688 101370
rect 70636 101306 70688 101312
rect 70912 101364 70964 101370
rect 70912 101306 70964 101312
rect 72016 101364 72068 101370
rect 72016 101306 72068 101312
rect 67534 99726 67732 99754
rect 68624 99740 68652 101306
rect 69820 99740 69848 101306
rect 70924 99740 70952 101306
rect 72396 99754 72424 101374
rect 74052 101370 74080 111030
rect 76904 111026 76932 114822
rect 77444 111088 77496 111094
rect 77444 111030 77496 111036
rect 74684 111020 74736 111026
rect 74684 110962 74736 110968
rect 76892 111020 76944 111026
rect 76892 110962 76944 110968
rect 73120 101364 73172 101370
rect 73120 101306 73172 101312
rect 74040 101364 74092 101370
rect 74040 101306 74092 101312
rect 72042 99726 72424 99754
rect 73132 99740 73160 101306
rect 74696 99754 74724 110962
rect 75328 101568 75380 101574
rect 75328 101510 75380 101516
rect 74250 99726 74724 99754
rect 75340 99740 75368 101510
rect 77456 101370 77484 111030
rect 77548 101574 77576 114822
rect 79560 111156 79612 111162
rect 79560 111098 79612 111104
rect 77536 101568 77588 101574
rect 77536 101510 77588 101516
rect 77536 101432 77588 101438
rect 77536 101374 77588 101380
rect 76432 101364 76484 101370
rect 76432 101306 76484 101312
rect 77444 101364 77496 101370
rect 77444 101306 77496 101312
rect 76444 99740 76472 101306
rect 77548 99740 77576 101374
rect 79572 101370 79600 111098
rect 79756 111094 79784 114822
rect 80940 111496 80992 111502
rect 80940 111438 80992 111444
rect 79744 111088 79796 111094
rect 79744 111030 79796 111036
rect 79652 111020 79704 111026
rect 79652 110962 79704 110968
rect 79664 101438 79692 110962
rect 79652 101432 79704 101438
rect 79652 101374 79704 101380
rect 80848 101432 80900 101438
rect 80848 101374 80900 101380
rect 78640 101364 78692 101370
rect 78640 101306 78692 101312
rect 79560 101364 79612 101370
rect 79560 101306 79612 101312
rect 79744 101364 79796 101370
rect 79744 101306 79796 101312
rect 78652 99740 78680 101306
rect 79756 99740 79784 101306
rect 80860 99740 80888 101374
rect 80952 101370 80980 111438
rect 81228 111026 81256 114822
rect 82320 111632 82372 111638
rect 82320 111574 82372 111580
rect 81216 111020 81268 111026
rect 81216 110962 81268 110968
rect 82332 101438 82360 111574
rect 82608 111162 82636 114822
rect 83700 111564 83752 111570
rect 83700 111506 83752 111512
rect 82596 111156 82648 111162
rect 82596 111098 82648 111104
rect 83148 101976 83200 101982
rect 83148 101918 83200 101924
rect 82320 101432 82372 101438
rect 82320 101374 82372 101380
rect 80940 101364 80992 101370
rect 80940 101306 80992 101312
rect 81952 101364 82004 101370
rect 81952 101306 82004 101312
rect 81964 99740 81992 101306
rect 83160 99740 83188 101918
rect 83712 101370 83740 111506
rect 84080 111502 84108 114822
rect 85460 111638 85488 114822
rect 85724 112380 85776 112386
rect 85724 112322 85776 112328
rect 85448 111632 85500 111638
rect 85448 111574 85500 111580
rect 84068 111496 84120 111502
rect 84068 111438 84120 111444
rect 83700 101364 83752 101370
rect 83700 101306 83752 101312
rect 85736 99754 85764 112322
rect 87208 111570 87236 114822
rect 90428 112250 90456 114822
rect 90416 112244 90468 112250
rect 90416 112186 90468 112192
rect 87196 111564 87248 111570
rect 87196 111506 87248 111512
rect 88668 102112 88720 102118
rect 88668 102054 88720 102060
rect 87564 102044 87616 102050
rect 87564 101986 87616 101992
rect 86460 101976 86512 101982
rect 86460 101918 86512 101924
rect 85382 99726 85764 99754
rect 86472 99740 86500 101918
rect 87576 99740 87604 101986
rect 88680 99740 88708 102054
rect 90612 101370 90640 115110
rect 89772 101364 89824 101370
rect 89772 101306 89824 101312
rect 90600 101364 90652 101370
rect 90600 101306 90652 101312
rect 89784 99740 89812 101306
rect 91256 99754 91284 115178
rect 92636 101370 92664 116470
rect 92900 116460 92952 116466
rect 92900 116402 92952 116408
rect 92808 116392 92860 116398
rect 92808 116334 92860 116340
rect 92716 116324 92768 116330
rect 92716 116266 92768 116272
rect 92728 116233 92756 116266
rect 92714 116224 92770 116233
rect 92714 116159 92770 116168
rect 92820 115825 92848 116334
rect 92806 115816 92862 115825
rect 92806 115751 92862 115760
rect 92912 115553 92940 116402
rect 92898 115544 92954 115553
rect 92898 115479 92954 115488
rect 93360 112244 93412 112250
rect 93360 112186 93412 112192
rect 93372 102458 93400 112186
rect 93360 102452 93412 102458
rect 93360 102394 93412 102400
rect 94016 101370 94044 116538
rect 94188 102452 94240 102458
rect 94188 102394 94240 102400
rect 91980 101364 92032 101370
rect 91980 101306 92032 101312
rect 92624 101364 92676 101370
rect 92624 101306 92676 101312
rect 93084 101364 93136 101370
rect 93084 101306 93136 101312
rect 94004 101364 94056 101370
rect 94004 101306 94056 101312
rect 90902 99726 91284 99754
rect 91992 99740 92020 101306
rect 93096 99740 93124 101306
rect 94200 99740 94228 102394
rect 44416 74368 44468 74374
rect 44416 74310 44468 74316
rect 53340 74368 53392 74374
rect 53340 74310 53392 74316
rect 23622 69848 23678 69857
rect 23622 69783 23678 69792
rect 23636 63193 23664 69783
rect 53352 66593 53380 74310
rect 53338 66584 53394 66593
rect 53338 66519 53394 66528
rect 44414 64816 44470 64825
rect 44414 64751 44470 64760
rect 23622 63184 23678 63193
rect 23622 63119 23678 63128
rect 26502 60026 26792 60042
rect 26502 60020 26804 60026
rect 26502 60014 26752 60020
rect 26752 59962 26804 59968
rect 26936 60020 26988 60026
rect 26936 59962 26988 59968
rect 25108 59878 26134 59906
rect 26672 59878 26870 59906
rect 13320 57844 13372 57850
rect 13320 57786 13372 57792
rect 13332 44153 13360 57786
rect 22244 50092 22296 50098
rect 22244 50034 22296 50040
rect 21508 50024 21560 50030
rect 21508 49966 21560 49972
rect 20864 49888 20916 49894
rect 20864 49830 20916 49836
rect 20220 49548 20272 49554
rect 20220 49490 20272 49496
rect 20232 46428 20260 49490
rect 20876 46428 20904 49830
rect 21520 46428 21548 49966
rect 22256 46428 22284 50034
rect 25108 49894 25136 59878
rect 26568 57164 26620 57170
rect 26568 57106 26620 57112
rect 26476 57096 26528 57102
rect 26476 57038 26528 57044
rect 25648 50228 25700 50234
rect 25648 50170 25700 50176
rect 25096 49888 25148 49894
rect 25096 49830 25148 49836
rect 23624 49752 23676 49758
rect 23624 49694 23676 49700
rect 22888 49276 22940 49282
rect 22888 49218 22940 49224
rect 22900 46428 22928 49218
rect 23636 46428 23664 49694
rect 24268 49684 24320 49690
rect 24268 49626 24320 49632
rect 24280 46428 24308 49626
rect 24912 49412 24964 49418
rect 24912 49354 24964 49360
rect 24924 46428 24952 49354
rect 25660 46428 25688 50170
rect 26488 49894 26516 57038
rect 26476 49888 26528 49894
rect 26476 49830 26528 49836
rect 26292 49752 26344 49758
rect 26292 49694 26344 49700
rect 26304 46428 26332 49694
rect 26580 49282 26608 57106
rect 26672 50098 26700 59878
rect 26660 50092 26712 50098
rect 26660 50034 26712 50040
rect 26948 50030 26976 59962
rect 27040 59878 27330 59906
rect 27408 59878 27698 59906
rect 27960 59878 28066 59906
rect 28236 59878 28526 59906
rect 28604 59878 28894 59906
rect 29262 59878 29552 59906
rect 27040 57170 27068 59878
rect 27028 57164 27080 57170
rect 27028 57106 27080 57112
rect 27408 57102 27436 59878
rect 27856 57164 27908 57170
rect 27856 57106 27908 57112
rect 27396 57096 27448 57102
rect 27396 57038 27448 57044
rect 27868 50234 27896 57106
rect 27856 50228 27908 50234
rect 27856 50170 27908 50176
rect 26936 50024 26988 50030
rect 26936 49966 26988 49972
rect 27960 49826 27988 59878
rect 28236 57186 28264 59878
rect 28052 57158 28264 57186
rect 28604 57170 28632 59878
rect 29144 57368 29196 57374
rect 29144 57310 29196 57316
rect 28592 57164 28644 57170
rect 27948 49820 28000 49826
rect 27948 49762 28000 49768
rect 28052 49418 28080 57158
rect 28592 57106 28644 57112
rect 29156 50234 29184 57310
rect 29328 57164 29380 57170
rect 29328 57106 29380 57112
rect 28316 50228 28368 50234
rect 28316 50170 28368 50176
rect 29144 50228 29196 50234
rect 29144 50170 29196 50176
rect 28040 49412 28092 49418
rect 28040 49354 28092 49360
rect 26568 49276 26620 49282
rect 26568 49218 26620 49224
rect 27672 49276 27724 49282
rect 27672 49218 27724 49224
rect 27028 49072 27080 49078
rect 27028 49014 27080 49020
rect 27040 46428 27068 49014
rect 27684 46428 27712 49218
rect 28328 46428 28356 50170
rect 29052 50160 29104 50166
rect 29052 50102 29104 50108
rect 29064 46428 29092 50102
rect 29340 49078 29368 57106
rect 29420 57096 29472 57102
rect 29420 57038 29472 57044
rect 29432 49282 29460 57038
rect 29524 49758 29552 59878
rect 29616 59878 29722 59906
rect 29800 59878 30090 59906
rect 29616 57170 29644 59878
rect 29604 57164 29656 57170
rect 29604 57106 29656 57112
rect 29800 57102 29828 59878
rect 30444 57374 30472 59892
rect 30720 59878 30918 59906
rect 30432 57368 30484 57374
rect 30432 57310 30484 57316
rect 30432 57232 30484 57238
rect 30432 57174 30484 57180
rect 29788 57096 29840 57102
rect 29788 57038 29840 57044
rect 30444 50234 30472 57174
rect 30524 57164 30576 57170
rect 30524 57106 30576 57112
rect 29696 50228 29748 50234
rect 29696 50170 29748 50176
rect 30432 50228 30484 50234
rect 30432 50170 30484 50176
rect 29512 49752 29564 49758
rect 29512 49694 29564 49700
rect 29420 49276 29472 49282
rect 29420 49218 29472 49224
rect 29328 49072 29380 49078
rect 29328 49014 29380 49020
rect 29708 46428 29736 50170
rect 30536 46442 30564 57106
rect 30720 50166 30748 59878
rect 31272 57238 31300 59892
rect 31260 57232 31312 57238
rect 31260 57174 31312 57180
rect 31640 57170 31668 59892
rect 32008 59878 32114 59906
rect 32192 59878 32482 59906
rect 32560 59878 32850 59906
rect 32008 57186 32036 59878
rect 32192 57186 32220 59878
rect 31628 57164 31680 57170
rect 31628 57106 31680 57112
rect 31824 57158 32036 57186
rect 32100 57158 32220 57186
rect 31824 50234 31852 57158
rect 32100 57050 32128 57158
rect 31916 57022 32128 57050
rect 31076 50228 31128 50234
rect 31076 50170 31128 50176
rect 31812 50228 31864 50234
rect 31812 50170 31864 50176
rect 30708 50160 30760 50166
rect 30708 50102 30760 50108
rect 30458 46414 30564 46442
rect 31088 46428 31116 50170
rect 31916 46442 31944 57022
rect 32560 56914 32588 59878
rect 33296 57170 33324 59892
rect 33388 59878 33678 59906
rect 33284 57164 33336 57170
rect 33284 57106 33336 57112
rect 31838 46414 31944 46442
rect 32008 56886 32588 56914
rect 32008 46442 32036 56886
rect 32088 56824 32140 56830
rect 32088 56766 32140 56772
rect 32100 46714 32128 56766
rect 32100 46686 32864 46714
rect 32836 46442 32864 46686
rect 33388 46442 33416 59878
rect 34124 57170 34152 59892
rect 34506 59878 34704 59906
rect 34874 59878 34980 59906
rect 33468 57164 33520 57170
rect 33468 57106 33520 57112
rect 34112 57164 34164 57170
rect 34112 57106 34164 57112
rect 33480 50302 33508 57106
rect 33468 50296 33520 50302
rect 33468 50238 33520 50244
rect 34296 50296 34348 50302
rect 34296 50238 34348 50244
rect 34308 46442 34336 50238
rect 34676 48890 34704 59878
rect 34676 48862 34888 48890
rect 34860 46442 34888 48862
rect 34952 46714 34980 59878
rect 35320 57170 35348 59892
rect 35702 59878 35992 59906
rect 35308 57164 35360 57170
rect 35308 57106 35360 57112
rect 35964 50114 35992 59878
rect 36056 58682 36084 59892
rect 36056 58654 36176 58682
rect 36148 58530 36176 58654
rect 36136 58524 36188 58530
rect 36136 58466 36188 58472
rect 36516 57170 36544 59892
rect 36884 57306 36912 59892
rect 36872 57300 36924 57306
rect 36872 57242 36924 57248
rect 37252 57238 37280 59892
rect 37608 58524 37660 58530
rect 37608 58466 37660 58472
rect 37240 57232 37292 57238
rect 37240 57174 37292 57180
rect 36044 57164 36096 57170
rect 36044 57106 36096 57112
rect 36504 57164 36556 57170
rect 36504 57106 36556 57112
rect 37516 57164 37568 57170
rect 37516 57106 37568 57112
rect 36056 50250 36084 57106
rect 36056 50222 36268 50250
rect 35964 50086 36176 50114
rect 36148 48942 36176 50086
rect 36136 48936 36188 48942
rect 36136 48878 36188 48884
rect 34952 46686 35624 46714
rect 35596 46442 35624 46686
rect 36240 46442 36268 50222
rect 37528 50098 37556 57106
rect 37516 50092 37568 50098
rect 37516 50034 37568 50040
rect 37240 48936 37292 48942
rect 37240 48878 37292 48884
rect 32008 46414 32482 46442
rect 32836 46414 33126 46442
rect 33388 46414 33862 46442
rect 34308 46414 34506 46442
rect 34860 46414 35242 46442
rect 35596 46414 35886 46442
rect 36240 46414 36530 46442
rect 37252 46428 37280 48878
rect 37620 46442 37648 58466
rect 37712 57374 37740 59892
rect 37700 57368 37752 57374
rect 37700 57310 37752 57316
rect 38080 57170 38108 59892
rect 38252 57300 38304 57306
rect 38252 57242 38304 57248
rect 38160 57232 38212 57238
rect 38160 57174 38212 57180
rect 38068 57164 38120 57170
rect 38068 57106 38120 57112
rect 38172 50166 38200 57174
rect 38264 50234 38292 57242
rect 38448 57238 38476 59892
rect 38908 57306 38936 59892
rect 39276 57510 39304 59892
rect 39264 57504 39316 57510
rect 39264 57446 39316 57452
rect 39644 57442 39672 59892
rect 40104 57578 40132 59892
rect 40092 57572 40144 57578
rect 40092 57514 40144 57520
rect 39632 57436 39684 57442
rect 39632 57378 39684 57384
rect 40276 57368 40328 57374
rect 40276 57310 40328 57316
rect 38896 57300 38948 57306
rect 38896 57242 38948 57248
rect 38436 57232 38488 57238
rect 38436 57174 38488 57180
rect 38252 50228 38304 50234
rect 38252 50170 38304 50176
rect 39264 50228 39316 50234
rect 39264 50170 39316 50176
rect 38160 50160 38212 50166
rect 38160 50102 38212 50108
rect 38252 50092 38304 50098
rect 38252 50034 38304 50040
rect 38264 46442 38292 50034
rect 37620 46414 37910 46442
rect 38264 46414 38646 46442
rect 39276 46428 39304 50170
rect 40000 50160 40052 50166
rect 40000 50102 40052 50108
rect 40012 46428 40040 50102
rect 40288 46442 40316 57310
rect 40472 57170 40500 59892
rect 40840 57782 40868 59892
rect 41300 58462 41328 59892
rect 41288 58456 41340 58462
rect 41288 58398 41340 58404
rect 41668 58394 41696 59892
rect 41656 58388 41708 58394
rect 41656 58330 41708 58336
rect 40828 57776 40880 57782
rect 40828 57718 40880 57724
rect 43772 57572 43824 57578
rect 43772 57514 43824 57520
rect 43036 57504 43088 57510
rect 43036 57446 43088 57452
rect 41840 57300 41892 57306
rect 41840 57242 41892 57248
rect 40920 57232 40972 57238
rect 40920 57174 40972 57180
rect 40368 57164 40420 57170
rect 40368 57106 40420 57112
rect 40460 57164 40512 57170
rect 40460 57106 40512 57112
rect 40380 46714 40408 57106
rect 40932 50234 40960 57174
rect 41852 50386 41880 57242
rect 41852 50358 42432 50386
rect 40920 50228 40972 50234
rect 40920 50170 40972 50176
rect 42024 50228 42076 50234
rect 42024 50170 42076 50176
rect 40380 46686 40960 46714
rect 40932 46442 40960 46686
rect 40288 46414 40670 46442
rect 40932 46414 41314 46442
rect 42036 46428 42064 50170
rect 42404 46442 42432 50358
rect 43048 46442 43076 57446
rect 43128 57436 43180 57442
rect 43128 57378 43180 57384
rect 43140 46714 43168 57378
rect 43680 57164 43732 57170
rect 43680 57106 43732 57112
rect 43692 49826 43720 57106
rect 43784 50234 43812 57514
rect 43772 50228 43824 50234
rect 43772 50170 43824 50176
rect 43680 49820 43732 49826
rect 43680 49762 43732 49768
rect 44428 49554 44456 64751
rect 45888 58456 45940 58462
rect 45888 58398 45940 58404
rect 45796 57776 45848 57782
rect 45796 57718 45848 57724
rect 44692 50228 44744 50234
rect 44692 50170 44744 50176
rect 44416 49548 44468 49554
rect 44416 49490 44468 49496
rect 43140 46686 43720 46714
rect 43692 46442 43720 46686
rect 42404 46414 42694 46442
rect 43048 46414 43430 46442
rect 43692 46414 44074 46442
rect 44704 46428 44732 50170
rect 45428 49820 45480 49826
rect 45428 49762 45480 49768
rect 45440 46428 45468 49762
rect 45808 46442 45836 57718
rect 45900 46714 45928 58398
rect 46440 58388 46492 58394
rect 46440 58330 46492 58336
rect 46452 50234 46480 58330
rect 46440 50228 46492 50234
rect 46440 50170 46492 50176
rect 47452 50228 47504 50234
rect 47452 50170 47504 50176
rect 45900 46686 46204 46714
rect 46176 46442 46204 46686
rect 45808 46414 46098 46442
rect 46176 46414 46834 46442
rect 47464 46428 47492 50170
rect 53352 47106 53380 66519
rect 59240 58433 59268 59892
rect 72580 58462 72608 59892
rect 79204 58530 79232 59892
rect 79192 58524 79244 58530
rect 79192 58466 79244 58472
rect 72568 58456 72620 58462
rect 59226 58424 59282 58433
rect 72568 58398 72620 58404
rect 59226 58359 59282 58368
rect 70544 57912 70596 57918
rect 70544 57854 70596 57860
rect 50396 47100 50448 47106
rect 50396 47042 50448 47048
rect 53340 47100 53392 47106
rect 53340 47042 53392 47048
rect 50408 46873 50436 47042
rect 50394 46864 50450 46873
rect 50394 46799 50450 46808
rect 50580 46488 50632 46494
rect 50580 46430 50632 46436
rect 61344 46488 61396 46494
rect 61344 46430 61396 46436
rect 13318 44144 13374 44153
rect 13318 44079 13374 44088
rect 50026 43736 50082 43745
rect 50026 43671 50082 43680
rect 50040 43570 50068 43671
rect 50028 43564 50080 43570
rect 50028 43506 50080 43512
rect 50210 42920 50266 42929
rect 50210 42855 50266 42864
rect 50224 42618 50252 42855
rect 50212 42612 50264 42618
rect 50212 42554 50264 42560
rect 18102 39384 18158 39393
rect 18102 39319 18158 39328
rect 18116 39218 18144 39319
rect 13320 39212 13372 39218
rect 13320 39154 13372 39160
rect 18104 39212 18156 39218
rect 18104 39154 18156 39160
rect 13332 20625 13360 39154
rect 50026 35712 50082 35721
rect 50026 35647 50082 35656
rect 50040 35274 50068 35647
rect 50028 35268 50080 35274
rect 50028 35210 50080 35216
rect 50210 34488 50266 34497
rect 50210 34423 50266 34432
rect 50224 33778 50252 34423
rect 50212 33772 50264 33778
rect 50212 33714 50264 33720
rect 50026 32720 50082 32729
rect 50026 32655 50082 32664
rect 50040 32350 50068 32655
rect 50028 32344 50080 32350
rect 50028 32286 50080 32292
rect 50486 26192 50542 26201
rect 50486 26127 50542 26136
rect 18102 25512 18158 25521
rect 50500 25482 50528 26127
rect 18102 25447 18158 25456
rect 50488 25476 50540 25482
rect 13318 20616 13374 20625
rect 13318 20551 13374 20560
rect 18116 18478 18144 25447
rect 50488 25418 50540 25424
rect 50210 23200 50266 23209
rect 50210 23135 50266 23144
rect 50224 22694 50252 23135
rect 50212 22688 50264 22694
rect 50212 22630 50264 22636
rect 50592 19265 50620 46430
rect 50764 46420 50816 46426
rect 50764 46362 50816 46368
rect 50672 46216 50724 46222
rect 50672 46158 50724 46164
rect 50684 21169 50712 46158
rect 50670 21160 50726 21169
rect 50670 21095 50726 21104
rect 50776 19809 50804 46362
rect 50856 46352 50908 46358
rect 50856 46294 50908 46300
rect 50868 20489 50896 46294
rect 51040 46284 51092 46290
rect 51040 46226 51092 46232
rect 50948 46148 51000 46154
rect 50948 46090 51000 46096
rect 50960 21849 50988 46090
rect 50946 21840 51002 21849
rect 50946 21775 51002 21784
rect 51052 21033 51080 46226
rect 51314 45232 51370 45241
rect 51314 45167 51370 45176
rect 51222 44824 51278 44833
rect 51222 44759 51224 44768
rect 51276 44759 51278 44768
rect 51224 44730 51276 44736
rect 51328 44658 51356 45167
rect 61356 44810 61384 46430
rect 62816 46420 62868 46426
rect 62816 46362 62868 46368
rect 62828 44810 62856 46362
rect 64288 46352 64340 46358
rect 64288 46294 64340 46300
rect 64300 44810 64328 46294
rect 65760 46284 65812 46290
rect 65760 46226 65812 46232
rect 65772 44810 65800 46226
rect 67324 46216 67376 46222
rect 67324 46158 67376 46164
rect 67336 44810 67364 46158
rect 68796 46148 68848 46154
rect 68796 46090 68848 46096
rect 68808 44810 68836 46090
rect 70556 44810 70584 57854
rect 72580 57850 72608 58398
rect 79204 58297 79232 58466
rect 79190 58288 79246 58297
rect 79190 58223 79246 58232
rect 92544 57918 92572 59892
rect 96132 58530 96160 151626
rect 98800 142986 98828 154375
rect 98880 151752 98932 151758
rect 98880 151694 98932 151700
rect 98788 142980 98840 142986
rect 98788 142922 98840 142928
rect 97408 137472 97460 137478
rect 97408 137414 97460 137420
rect 97420 137002 97448 137414
rect 98052 137268 98104 137274
rect 98052 137210 98104 137216
rect 97408 136996 97460 137002
rect 97408 136938 97460 136944
rect 97960 135908 98012 135914
rect 97960 135850 98012 135856
rect 97972 134282 98000 135850
rect 98064 135710 98092 137210
rect 98144 135840 98196 135846
rect 98144 135782 98196 135788
rect 98052 135704 98104 135710
rect 98052 135646 98104 135652
rect 98156 134350 98184 135782
rect 98144 134344 98196 134350
rect 98144 134286 98196 134292
rect 97960 134276 98012 134282
rect 97960 134218 98012 134224
rect 98052 126252 98104 126258
rect 98052 126194 98104 126200
rect 98064 124694 98092 126194
rect 98144 126184 98196 126190
rect 98144 126126 98196 126132
rect 98052 124688 98104 124694
rect 98052 124630 98104 124636
rect 98156 124626 98184 126126
rect 98144 124620 98196 124626
rect 98144 124562 98196 124568
rect 97500 120812 97552 120818
rect 97500 120754 97552 120760
rect 97512 119118 97540 120754
rect 97960 120744 98012 120750
rect 97960 120686 98012 120692
rect 97868 119384 97920 119390
rect 97868 119326 97920 119332
rect 97500 119112 97552 119118
rect 97500 119054 97552 119060
rect 97880 117758 97908 119326
rect 97972 119186 98000 120686
rect 98144 120676 98196 120682
rect 98144 120618 98196 120624
rect 98052 119316 98104 119322
rect 98052 119258 98104 119264
rect 97960 119180 98012 119186
rect 97960 119122 98012 119128
rect 97960 117956 98012 117962
rect 97960 117898 98012 117904
rect 97868 117752 97920 117758
rect 97868 117694 97920 117700
rect 97972 116330 98000 117898
rect 98064 117826 98092 119258
rect 98156 119254 98184 120618
rect 98144 119248 98196 119254
rect 98144 119190 98196 119196
rect 98144 117888 98196 117894
rect 98144 117830 98196 117836
rect 98052 117820 98104 117826
rect 98052 117762 98104 117768
rect 98156 116398 98184 117830
rect 98144 116392 98196 116398
rect 98144 116334 98196 116340
rect 97960 116324 98012 116330
rect 97960 116266 98012 116272
rect 98788 110272 98840 110278
rect 98788 110214 98840 110220
rect 98800 99777 98828 110214
rect 98786 99768 98842 99777
rect 98786 99703 98842 99712
rect 98788 97216 98840 97222
rect 98788 97158 98840 97164
rect 98696 93068 98748 93074
rect 98696 93010 98748 93016
rect 98708 87401 98736 93010
rect 98800 89985 98828 97158
rect 98786 89976 98842 89985
rect 98786 89911 98842 89920
rect 98694 87392 98750 87401
rect 98694 87327 98750 87336
rect 98234 75560 98290 75569
rect 98234 75495 98290 75504
rect 98248 75122 98276 75495
rect 98236 75116 98288 75122
rect 98236 75058 98288 75064
rect 96120 58524 96172 58530
rect 96120 58466 96172 58472
rect 98892 58462 98920 151694
rect 98984 143394 99012 162807
rect 99062 161648 99118 161657
rect 99062 161583 99118 161592
rect 99076 143462 99104 161583
rect 99154 160424 99210 160433
rect 99154 160359 99210 160368
rect 99168 143598 99196 160359
rect 99430 159200 99486 159209
rect 99430 159135 99486 159144
rect 99246 157976 99302 157985
rect 99246 157911 99302 157920
rect 99156 143592 99208 143598
rect 99156 143534 99208 143540
rect 99064 143456 99116 143462
rect 99064 143398 99116 143404
rect 98972 143388 99024 143394
rect 98972 143330 99024 143336
rect 99260 142918 99288 157911
rect 99338 156752 99394 156761
rect 99338 156687 99394 156696
rect 99248 142912 99300 142918
rect 99248 142854 99300 142860
rect 99352 142850 99380 156687
rect 99444 143530 99472 159135
rect 99522 155528 99578 155537
rect 99522 155463 99578 155472
rect 99432 143524 99484 143530
rect 99432 143466 99484 143472
rect 99340 142844 99392 142850
rect 99340 142786 99392 142792
rect 99536 142782 99564 155463
rect 104412 155090 104440 163390
rect 106896 161929 106924 167606
rect 183716 167602 183744 168791
rect 183794 167768 183850 167777
rect 183794 167703 183850 167712
rect 183704 167596 183756 167602
rect 183704 167538 183756 167544
rect 182874 166544 182930 166553
rect 182874 166479 182876 166488
rect 182928 166479 182930 166488
rect 182876 166450 182928 166456
rect 107252 166236 107304 166242
rect 107252 166178 107304 166184
rect 107160 164808 107212 164814
rect 107160 164750 107212 164756
rect 106882 161920 106938 161929
rect 106882 161855 106938 161864
rect 107172 157305 107200 164750
rect 107264 159617 107292 166178
rect 183702 165320 183758 165329
rect 183702 165255 183758 165264
rect 183716 165018 183744 165255
rect 183704 165012 183756 165018
rect 183704 164954 183756 164960
rect 183058 164096 183114 164105
rect 183058 164031 183114 164040
rect 128502 163824 128558 163833
rect 128502 163759 128558 163768
rect 128516 163454 128544 163759
rect 183072 163454 183100 164031
rect 128504 163448 128556 163454
rect 128504 163390 128556 163396
rect 137520 163448 137572 163454
rect 137520 163390 137572 163396
rect 183060 163448 183112 163454
rect 183060 163390 183112 163396
rect 137532 160569 137560 163390
rect 183808 163046 183836 167703
rect 191340 167596 191392 167602
rect 191340 167538 191392 167544
rect 187936 166508 187988 166514
rect 187936 166450 187988 166456
rect 183796 163040 183848 163046
rect 183796 162982 183848 162988
rect 183058 162872 183114 162881
rect 183058 162807 183114 162816
rect 137518 160560 137574 160569
rect 137518 160495 137574 160504
rect 107250 159608 107306 159617
rect 107250 159543 107306 159552
rect 107158 157296 107214 157305
rect 107158 157231 107214 157240
rect 137532 156761 137560 160495
rect 137518 156752 137574 156761
rect 137518 156687 137574 156696
rect 104400 155084 104452 155090
rect 104400 155026 104452 155032
rect 106516 155084 106568 155090
rect 106516 155026 106568 155032
rect 106528 154993 106556 155026
rect 106514 154984 106570 154993
rect 106514 154919 106570 154928
rect 110116 152098 110144 153868
rect 110208 153854 110498 153882
rect 110668 153854 110866 153882
rect 109184 152092 109236 152098
rect 109184 152034 109236 152040
rect 110104 152092 110156 152098
rect 110104 152034 110156 152040
rect 106700 143592 106752 143598
rect 106700 143534 106752 143540
rect 106608 143524 106660 143530
rect 106608 143466 106660 143472
rect 103940 142980 103992 142986
rect 103940 142922 103992 142928
rect 99524 142776 99576 142782
rect 99524 142718 99576 142724
rect 103952 140826 103980 142922
rect 105596 142912 105648 142918
rect 105596 142854 105648 142860
rect 105136 142844 105188 142850
rect 105136 142786 105188 142792
rect 104492 142776 104544 142782
rect 104492 142718 104544 142724
rect 104504 140826 104532 142718
rect 105148 140826 105176 142786
rect 105608 140826 105636 142854
rect 103952 140798 104242 140826
rect 104504 140798 104794 140826
rect 105148 140798 105346 140826
rect 105608 140798 105990 140826
rect 106620 140690 106648 143466
rect 106712 140826 106740 143534
rect 107436 143456 107488 143462
rect 107436 143398 107488 143404
rect 107448 140826 107476 143398
rect 107988 143388 108040 143394
rect 107988 143330 108040 143336
rect 108000 140826 108028 143330
rect 106712 140798 107094 140826
rect 107448 140798 107738 140826
rect 108000 140798 108290 140826
rect 109196 140690 109224 152034
rect 110208 151078 110236 153854
rect 110668 152250 110696 153854
rect 110932 152364 110984 152370
rect 110932 152306 110984 152312
rect 110484 152222 110696 152250
rect 109368 151072 109420 151078
rect 109368 151014 109420 151020
rect 110196 151072 110248 151078
rect 110196 151014 110248 151020
rect 109380 140826 109408 151014
rect 110484 143666 110512 152222
rect 110564 150936 110616 150942
rect 110944 150890 110972 152306
rect 111312 151010 111340 153868
rect 111680 152370 111708 153868
rect 111668 152364 111720 152370
rect 111668 152306 111720 152312
rect 111300 151004 111352 151010
rect 112048 150992 112076 153868
rect 112128 151888 112180 151894
rect 112128 151830 112180 151836
rect 111300 150946 111352 150952
rect 111956 150964 112076 150992
rect 110564 150878 110616 150884
rect 110196 143660 110248 143666
rect 110196 143602 110248 143608
rect 110472 143660 110524 143666
rect 110472 143602 110524 143608
rect 109380 140798 109486 140826
rect 110208 140690 110236 143602
rect 110576 140962 110604 150878
rect 110484 140934 110604 140962
rect 110668 150862 110972 150890
rect 110484 140826 110512 140934
rect 110484 140798 110590 140826
rect 106542 140662 106648 140690
rect 108842 140662 109224 140690
rect 110038 140662 110236 140690
rect 110668 140690 110696 150862
rect 111956 140690 111984 150964
rect 112140 143666 112168 151830
rect 112128 143660 112180 143666
rect 112128 143602 112180 143608
rect 112508 140690 112536 153868
rect 112876 151894 112904 153868
rect 112864 151888 112916 151894
rect 112864 151830 112916 151836
rect 112588 143660 112640 143666
rect 112588 143602 112640 143608
rect 112600 140826 112628 143602
rect 113244 142594 113272 153868
rect 113600 152364 113652 152370
rect 113600 152306 113652 152312
rect 113612 143530 113640 152306
rect 113600 143524 113652 143530
rect 113600 143466 113652 143472
rect 113244 142566 113456 142594
rect 113428 140826 113456 142566
rect 113704 140826 113732 153868
rect 114072 152370 114100 153868
rect 114060 152364 114112 152370
rect 114060 152306 114112 152312
rect 114440 143666 114468 153868
rect 114428 143660 114480 143666
rect 114428 143602 114480 143608
rect 114900 143598 114928 153868
rect 115268 151010 115296 153868
rect 115650 153854 115940 153882
rect 115256 151004 115308 151010
rect 115256 150946 115308 150952
rect 115808 151004 115860 151010
rect 115808 150946 115860 150952
rect 114980 143660 115032 143666
rect 114980 143602 115032 143608
rect 114888 143592 114940 143598
rect 114888 143534 114940 143540
rect 114428 143524 114480 143530
rect 114428 143466 114480 143472
rect 114440 140826 114468 143466
rect 114992 140826 115020 143602
rect 115532 143592 115584 143598
rect 115532 143534 115584 143540
rect 115544 140826 115572 143534
rect 115820 142866 115848 150946
rect 115912 143666 115940 153854
rect 115900 143660 115952 143666
rect 115900 143602 115952 143608
rect 116096 143598 116124 153868
rect 116464 151282 116492 153868
rect 116846 153854 117228 153882
rect 117306 153854 117504 153882
rect 117200 152386 117228 153854
rect 117200 152358 117412 152386
rect 116452 151276 116504 151282
rect 116452 151218 116504 151224
rect 117188 151276 117240 151282
rect 117188 151218 117240 151224
rect 116636 143660 116688 143666
rect 116636 143602 116688 143608
rect 116084 143592 116136 143598
rect 116084 143534 116136 143540
rect 115820 142838 116216 142866
rect 116188 140826 116216 142838
rect 116648 140826 116676 143602
rect 117200 142986 117228 151218
rect 117384 143122 117412 152358
rect 117476 143938 117504 153854
rect 117660 152370 117688 153868
rect 117648 152364 117700 152370
rect 117648 152306 117700 152312
rect 118120 151282 118148 153868
rect 118488 152302 118516 153868
rect 118764 153854 118870 153882
rect 118476 152296 118528 152302
rect 118476 152238 118528 152244
rect 118764 152234 118792 153854
rect 118844 152364 118896 152370
rect 118844 152306 118896 152312
rect 118752 152228 118804 152234
rect 118752 152170 118804 152176
rect 118108 151276 118160 151282
rect 118108 151218 118160 151224
rect 118856 144074 118884 152306
rect 119316 152098 119344 153868
rect 119684 152370 119712 153868
rect 119672 152364 119724 152370
rect 119672 152306 119724 152312
rect 120052 152166 120080 153868
rect 120040 152160 120092 152166
rect 120040 152102 120092 152108
rect 119304 152092 119356 152098
rect 119304 152034 119356 152040
rect 120512 151282 120540 153868
rect 120592 152296 120644 152302
rect 120592 152238 120644 152244
rect 120316 151276 120368 151282
rect 120316 151218 120368 151224
rect 120500 151276 120552 151282
rect 120500 151218 120552 151224
rect 118844 144068 118896 144074
rect 118844 144010 118896 144016
rect 119580 144068 119632 144074
rect 119580 144010 119632 144016
rect 117464 143932 117516 143938
rect 117464 143874 117516 143880
rect 119028 143932 119080 143938
rect 119028 143874 119080 143880
rect 117648 143592 117700 143598
rect 117648 143534 117700 143540
rect 117372 143116 117424 143122
rect 117372 143058 117424 143064
rect 117188 142980 117240 142986
rect 117188 142922 117240 142928
rect 112600 140798 112982 140826
rect 113428 140798 113534 140826
rect 113704 140798 114086 140826
rect 114440 140798 114730 140826
rect 114992 140798 115282 140826
rect 115544 140798 115834 140826
rect 116188 140798 116478 140826
rect 116648 140798 117030 140826
rect 117660 140690 117688 143534
rect 118476 143116 118528 143122
rect 118476 143058 118528 143064
rect 117924 142980 117976 142986
rect 117924 142922 117976 142928
rect 117936 140826 117964 142922
rect 118488 140826 118516 143058
rect 119040 140826 119068 143874
rect 119592 140826 119620 144010
rect 120328 140826 120356 151218
rect 120604 140826 120632 152238
rect 120880 151826 120908 153868
rect 120960 152228 121012 152234
rect 120960 152170 121012 152176
rect 120868 151820 120920 151826
rect 120868 151762 120920 151768
rect 120972 144074 121000 152170
rect 121248 151078 121276 153868
rect 121708 151418 121736 153868
rect 121972 152364 122024 152370
rect 121972 152306 122024 152312
rect 121788 152092 121840 152098
rect 121788 152034 121840 152040
rect 121696 151412 121748 151418
rect 121696 151354 121748 151360
rect 121236 151072 121288 151078
rect 121236 151014 121288 151020
rect 120960 144068 121012 144074
rect 120960 144010 121012 144016
rect 121696 144068 121748 144074
rect 121696 144010 121748 144016
rect 121708 140962 121736 144010
rect 121800 141098 121828 152034
rect 121984 149666 122012 152306
rect 122076 151010 122104 153868
rect 122444 151350 122472 153868
rect 122904 151962 122932 153868
rect 123168 152160 123220 152166
rect 123168 152102 123220 152108
rect 122892 151956 122944 151962
rect 122892 151898 122944 151904
rect 122432 151344 122484 151350
rect 122432 151286 122484 151292
rect 123076 151276 123128 151282
rect 123076 151218 123128 151224
rect 122064 151004 122116 151010
rect 122064 150946 122116 150952
rect 121984 149638 122472 149666
rect 121800 141070 122104 141098
rect 121708 140934 121828 140962
rect 117936 140798 118226 140826
rect 118488 140798 118778 140826
rect 119040 140798 119330 140826
rect 119592 140798 119974 140826
rect 120328 140798 120526 140826
rect 120604 140798 121078 140826
rect 121800 140690 121828 140934
rect 122076 140826 122104 141070
rect 122444 140826 122472 149638
rect 123088 146182 123116 151218
rect 123076 146176 123128 146182
rect 123076 146118 123128 146124
rect 123180 140826 123208 152102
rect 123272 151962 123300 153868
rect 123260 151956 123312 151962
rect 123260 151898 123312 151904
rect 123640 151622 123668 153868
rect 124100 152370 124128 153868
rect 124088 152364 124140 152370
rect 124088 152306 124140 152312
rect 124468 152098 124496 153868
rect 124836 152302 124864 153868
rect 124824 152296 124876 152302
rect 124824 152238 124876 152244
rect 124456 152092 124508 152098
rect 124456 152034 124508 152040
rect 123720 151820 123772 151826
rect 123720 151762 123772 151768
rect 123628 151616 123680 151622
rect 123628 151558 123680 151564
rect 123628 146176 123680 146182
rect 123628 146118 123680 146124
rect 123640 140826 123668 146118
rect 123732 144006 123760 151762
rect 124640 151412 124692 151418
rect 124640 151354 124692 151360
rect 123812 151072 123864 151078
rect 123812 151014 123864 151020
rect 123824 144074 123852 151014
rect 123812 144068 123864 144074
rect 123812 144010 123864 144016
rect 124548 144068 124600 144074
rect 124548 144010 124600 144016
rect 123720 144000 123772 144006
rect 123720 143942 123772 143948
rect 124456 144000 124508 144006
rect 124456 143942 124508 143948
rect 124468 140826 124496 143942
rect 124560 141098 124588 144010
rect 124652 143682 124680 151354
rect 125192 151344 125244 151350
rect 125192 151286 125244 151292
rect 125100 151004 125152 151010
rect 125100 150946 125152 150952
rect 125112 144074 125140 150946
rect 125100 144068 125152 144074
rect 125100 144010 125152 144016
rect 125204 144006 125232 151286
rect 125296 151078 125324 153868
rect 125664 151350 125692 153868
rect 127860 152364 127912 152370
rect 127860 152306 127912 152312
rect 127216 151956 127268 151962
rect 127216 151898 127268 151904
rect 125652 151344 125704 151350
rect 125652 151286 125704 151292
rect 125284 151072 125336 151078
rect 125284 151014 125336 151020
rect 127228 146182 127256 151898
rect 127308 151548 127360 151554
rect 127308 151490 127360 151496
rect 127216 146176 127268 146182
rect 127216 146118 127268 146124
rect 126020 144068 126072 144074
rect 126020 144010 126072 144016
rect 125192 144000 125244 144006
rect 125192 143942 125244 143948
rect 124652 143654 125416 143682
rect 124560 141070 124772 141098
rect 122076 140798 122274 140826
rect 122444 140798 122826 140826
rect 123180 140798 123470 140826
rect 123640 140798 124022 140826
rect 124468 140798 124574 140826
rect 110668 140662 111234 140690
rect 111786 140662 111984 140690
rect 112338 140662 112536 140690
rect 117582 140662 117688 140690
rect 121722 140662 121828 140690
rect 124744 140690 124772 141070
rect 125388 140826 125416 143654
rect 126032 140826 126060 144010
rect 126572 144000 126624 144006
rect 126572 143942 126624 143948
rect 126584 140826 126612 143942
rect 127320 140826 127348 151490
rect 127676 146176 127728 146182
rect 127676 146118 127728 146124
rect 127688 140826 127716 146118
rect 127872 144006 127900 152306
rect 129332 152296 129384 152302
rect 129332 152238 129384 152244
rect 128780 152092 128832 152098
rect 128780 152034 128832 152040
rect 127952 151616 128004 151622
rect 127952 151558 128004 151564
rect 127964 144074 127992 151558
rect 127952 144068 128004 144074
rect 127952 144010 128004 144016
rect 128596 144068 128648 144074
rect 128596 144010 128648 144016
rect 127860 144000 127912 144006
rect 127860 143942 127912 143948
rect 128608 140826 128636 144010
rect 128688 144000 128740 144006
rect 128688 143942 128740 143948
rect 128700 141098 128728 143942
rect 128792 143682 128820 152034
rect 129240 151072 129292 151078
rect 129240 151014 129292 151020
rect 129252 144006 129280 151014
rect 129344 144074 129372 152238
rect 131356 151344 131408 151350
rect 131356 151286 131408 151292
rect 129332 144068 129384 144074
rect 129332 144010 129384 144016
rect 130068 144068 130120 144074
rect 130068 144010 130120 144016
rect 129240 144000 129292 144006
rect 129240 143942 129292 143948
rect 128792 143654 129464 143682
rect 128700 141070 128820 141098
rect 125388 140798 125770 140826
rect 126032 140798 126322 140826
rect 126584 140798 126966 140826
rect 127320 140798 127518 140826
rect 127688 140798 128070 140826
rect 128608 140798 128714 140826
rect 128792 140690 128820 141070
rect 129436 140826 129464 143654
rect 130080 140826 130108 144010
rect 130620 144000 130672 144006
rect 130620 143942 130672 143948
rect 130632 140826 130660 143942
rect 131368 140826 131396 151286
rect 129436 140798 129818 140826
rect 130080 140798 130462 140826
rect 130632 140798 131014 140826
rect 131368 140798 131566 140826
rect 124744 140662 125218 140690
rect 128792 140662 129266 140690
rect 134850 140568 134906 140577
rect 134850 140503 134906 140512
rect 100810 140160 100866 140169
rect 100810 140095 100866 140104
rect 100824 138566 100852 140095
rect 134864 140062 134892 140503
rect 134852 140056 134904 140062
rect 100902 140024 100958 140033
rect 134852 139998 134904 140004
rect 135402 140024 135458 140033
rect 100902 139959 100958 139968
rect 135402 139959 135404 139968
rect 100812 138560 100864 138566
rect 100812 138502 100864 138508
rect 100916 138498 100944 139959
rect 135456 139959 135458 139968
rect 135404 139930 135456 139936
rect 134666 139480 134722 139489
rect 134666 139415 134722 139424
rect 101178 138936 101234 138945
rect 101178 138871 101234 138880
rect 101086 138800 101142 138809
rect 101086 138735 101142 138744
rect 100904 138492 100956 138498
rect 100904 138434 100956 138440
rect 101100 137070 101128 138735
rect 101192 137138 101220 138871
rect 134680 138634 134708 139415
rect 135402 138800 135458 138809
rect 135402 138735 135404 138744
rect 135456 138735 135458 138744
rect 135404 138706 135456 138712
rect 134668 138628 134720 138634
rect 134668 138570 134720 138576
rect 134666 138256 134722 138265
rect 134666 138191 134722 138200
rect 101822 137848 101878 137857
rect 101822 137783 101878 137792
rect 101270 137712 101326 137721
rect 101270 137647 101326 137656
rect 101284 137274 101312 137647
rect 101836 137478 101864 137783
rect 101824 137472 101876 137478
rect 101824 137414 101876 137420
rect 134680 137410 134708 138191
rect 135402 137712 135458 137721
rect 135402 137647 135458 137656
rect 134668 137404 134720 137410
rect 134668 137346 134720 137352
rect 101272 137268 101324 137274
rect 101272 137210 101324 137216
rect 135416 137206 135444 137647
rect 135404 137200 135456 137206
rect 135404 137142 135456 137148
rect 101180 137132 101232 137138
rect 101180 137074 101232 137080
rect 101088 137064 101140 137070
rect 101088 137006 101140 137012
rect 135034 137032 135090 137041
rect 135034 136967 135090 136976
rect 101178 136624 101234 136633
rect 101178 136559 101234 136568
rect 101192 135778 101220 136559
rect 101270 136080 101326 136089
rect 101270 136015 101326 136024
rect 101284 135914 101312 136015
rect 135048 135982 135076 136967
rect 135310 136488 135366 136497
rect 135310 136423 135366 136432
rect 135036 135976 135088 135982
rect 101730 135944 101786 135953
rect 101272 135908 101324 135914
rect 135036 135918 135088 135924
rect 135324 135914 135352 136423
rect 135402 135944 135458 135953
rect 101730 135879 101786 135888
rect 135312 135908 135364 135914
rect 101272 135850 101324 135856
rect 101744 135846 101772 135879
rect 135402 135879 135458 135888
rect 135312 135850 135364 135856
rect 135416 135846 135444 135879
rect 101732 135840 101784 135846
rect 101732 135782 101784 135788
rect 135404 135840 135456 135846
rect 135404 135782 135456 135788
rect 101180 135772 101232 135778
rect 101180 135714 101232 135720
rect 134850 135400 134906 135409
rect 134850 135335 134906 135344
rect 101822 134856 101878 134865
rect 101822 134791 101878 134800
rect 100902 134448 100958 134457
rect 101836 134418 101864 134791
rect 134482 134720 134538 134729
rect 134482 134655 134484 134664
rect 134536 134655 134538 134664
rect 134484 134626 134536 134632
rect 134864 134554 134892 135335
rect 136876 134684 136928 134690
rect 136876 134626 136928 134632
rect 134852 134548 134904 134554
rect 134852 134490 134904 134496
rect 100902 134383 100958 134392
rect 101824 134412 101876 134418
rect 100916 132922 100944 134383
rect 101824 134354 101876 134360
rect 135402 134176 135458 134185
rect 135402 134111 135458 134120
rect 101362 133768 101418 133777
rect 101362 133703 101418 133712
rect 101376 132990 101404 133703
rect 135034 133632 135090 133641
rect 135034 133567 135090 133576
rect 135048 133126 135076 133567
rect 135036 133120 135088 133126
rect 101730 133088 101786 133097
rect 135036 133062 135088 133068
rect 135416 133058 135444 134111
rect 101730 133023 101786 133032
rect 135404 133052 135456 133058
rect 101364 132984 101416 132990
rect 101364 132926 101416 132932
rect 100904 132916 100956 132922
rect 100904 132858 100956 132864
rect 101454 132000 101510 132009
rect 101454 131935 101510 131944
rect 101468 130202 101496 131935
rect 101638 131864 101694 131873
rect 101638 131799 101694 131808
rect 101652 130270 101680 131799
rect 101744 131562 101772 133023
rect 135404 132994 135456 133000
rect 135310 132952 135366 132961
rect 135310 132887 135366 132896
rect 101822 132544 101878 132553
rect 101822 132479 101878 132488
rect 101836 131630 101864 132479
rect 135034 131864 135090 131873
rect 135034 131799 135036 131808
rect 135088 131799 135090 131808
rect 135036 131770 135088 131776
rect 135324 131698 135352 132887
rect 136888 132854 136916 134626
rect 136876 132848 136928 132854
rect 136876 132790 136928 132796
rect 135402 132408 135458 132417
rect 135402 132343 135458 132352
rect 135416 132038 135444 132343
rect 135404 132032 135456 132038
rect 135404 131974 135456 131980
rect 137336 131828 137388 131834
rect 137336 131770 137388 131776
rect 135312 131692 135364 131698
rect 135312 131634 135364 131640
rect 101824 131624 101876 131630
rect 137348 131612 137376 131770
rect 101824 131566 101876 131572
rect 137256 131584 137376 131612
rect 101732 131556 101784 131562
rect 101732 131498 101784 131504
rect 135034 131320 135090 131329
rect 135034 131255 135090 131264
rect 101730 130776 101786 130785
rect 101730 130711 101786 130720
rect 101640 130264 101692 130270
rect 101640 130206 101692 130212
rect 101456 130196 101508 130202
rect 101456 130138 101508 130144
rect 101362 129688 101418 129697
rect 101362 129623 101418 129632
rect 101270 129008 101326 129017
rect 101270 128943 101326 128952
rect 100994 128464 101050 128473
rect 100994 128399 101050 128408
rect 101008 127482 101036 128399
rect 101178 127920 101234 127929
rect 101178 127855 101234 127864
rect 101086 127784 101142 127793
rect 101086 127719 101142 127728
rect 100996 127476 101048 127482
rect 100996 127418 101048 127424
rect 100994 126288 101050 126297
rect 100994 126223 101050 126232
rect 101008 126190 101036 126223
rect 100996 126184 101048 126190
rect 100996 126126 101048 126132
rect 101100 126054 101128 127719
rect 101192 126122 101220 127855
rect 101284 127414 101312 128943
rect 101376 128910 101404 129623
rect 101364 128904 101416 128910
rect 101364 128846 101416 128852
rect 101744 128774 101772 130711
rect 101822 130368 101878 130377
rect 135048 130338 135076 131255
rect 135402 130640 135458 130649
rect 135402 130575 135404 130584
rect 135456 130575 135458 130584
rect 135404 130546 135456 130552
rect 101822 130303 101878 130312
rect 135036 130332 135088 130338
rect 101836 128842 101864 130303
rect 135036 130274 135088 130280
rect 137256 130202 137284 131584
rect 137336 130332 137388 130338
rect 137336 130274 137388 130280
rect 137244 130196 137296 130202
rect 137244 130138 137296 130144
rect 135402 130096 135458 130105
rect 135402 130031 135458 130040
rect 135310 129552 135366 129561
rect 135310 129487 135366 129496
rect 135324 129386 135352 129487
rect 135312 129380 135364 129386
rect 135312 129322 135364 129328
rect 135416 128978 135444 130031
rect 135404 128972 135456 128978
rect 135404 128914 135456 128920
rect 135402 128872 135458 128881
rect 101824 128836 101876 128842
rect 137348 128842 137376 130274
rect 135402 128807 135458 128816
rect 137336 128836 137388 128842
rect 101824 128778 101876 128784
rect 101732 128768 101784 128774
rect 101732 128710 101784 128716
rect 134666 128328 134722 128337
rect 134666 128263 134722 128272
rect 134680 127618 134708 128263
rect 135310 127784 135366 127793
rect 135310 127719 135312 127728
rect 135364 127719 135366 127728
rect 135312 127690 135364 127696
rect 134668 127612 134720 127618
rect 134668 127554 134720 127560
rect 135416 127550 135444 128807
rect 137336 128778 137388 128784
rect 137428 127612 137480 127618
rect 137428 127554 137480 127560
rect 135404 127544 135456 127550
rect 135404 127486 135456 127492
rect 101272 127408 101324 127414
rect 101272 127350 101324 127356
rect 135402 127240 135458 127249
rect 135458 127198 135628 127226
rect 135402 127175 135458 127184
rect 101270 126696 101326 126705
rect 101270 126631 101326 126640
rect 101284 126258 101312 126631
rect 135402 126560 135458 126569
rect 135458 126518 135536 126546
rect 135402 126495 135458 126504
rect 101272 126252 101324 126258
rect 101272 126194 101324 126200
rect 101180 126116 101232 126122
rect 101180 126058 101232 126064
rect 101088 126048 101140 126054
rect 101088 125990 101140 125996
rect 135218 126016 135274 126025
rect 135218 125951 135274 125960
rect 100994 125608 101050 125617
rect 100994 125543 101050 125552
rect 101008 124762 101036 125543
rect 101270 125064 101326 125073
rect 101270 124999 101326 125008
rect 101086 124792 101142 124801
rect 100996 124756 101048 124762
rect 101086 124727 101142 124736
rect 100996 124698 101048 124704
rect 100994 123432 101050 123441
rect 100994 123367 101050 123376
rect 101008 121974 101036 123367
rect 101100 123334 101128 124727
rect 101178 123840 101234 123849
rect 101178 123775 101234 123784
rect 101088 123328 101140 123334
rect 101088 123270 101140 123276
rect 101086 122072 101142 122081
rect 101086 122007 101142 122016
rect 100996 121968 101048 121974
rect 100996 121910 101048 121916
rect 100994 121528 101050 121537
rect 100994 121463 101050 121472
rect 101008 120818 101036 121463
rect 100996 120812 101048 120818
rect 100996 120754 101048 120760
rect 100994 120712 101050 120721
rect 100994 120647 100996 120656
rect 101048 120647 101050 120656
rect 100996 120618 101048 120624
rect 101100 120614 101128 122007
rect 101192 121906 101220 123775
rect 101284 123266 101312 124999
rect 135232 124830 135260 125951
rect 135402 125472 135458 125481
rect 135402 125407 135404 125416
rect 135456 125407 135458 125416
rect 135404 125378 135456 125384
rect 135404 124892 135456 124898
rect 135404 124834 135456 124840
rect 135220 124824 135272 124830
rect 135416 124801 135444 124834
rect 135220 124766 135272 124772
rect 135402 124792 135458 124801
rect 135402 124727 135458 124736
rect 135508 124422 135536 126518
rect 135600 124762 135628 127198
rect 137440 126054 137468 127554
rect 137428 126048 137480 126054
rect 137428 125990 137480 125996
rect 136876 124892 136928 124898
rect 136876 124834 136928 124840
rect 135588 124756 135640 124762
rect 135588 124698 135640 124704
rect 135496 124416 135548 124422
rect 135496 124358 135548 124364
rect 134114 124248 134170 124257
rect 134114 124183 134170 124192
rect 134128 123402 134156 124183
rect 135034 123704 135090 123713
rect 135034 123639 135036 123648
rect 135088 123639 135090 123648
rect 135036 123610 135088 123616
rect 134116 123396 134168 123402
rect 134116 123338 134168 123344
rect 101272 123260 101324 123266
rect 101272 123202 101324 123208
rect 135218 123024 135274 123033
rect 135218 122959 135274 122968
rect 101270 122616 101326 122625
rect 135232 122586 135260 122959
rect 136888 122858 136916 124834
rect 137428 123668 137480 123674
rect 137428 123610 137480 123616
rect 136876 122852 136928 122858
rect 136876 122794 136928 122800
rect 101270 122551 101326 122560
rect 135220 122580 135272 122586
rect 101180 121900 101232 121906
rect 101180 121842 101232 121848
rect 101178 120848 101234 120857
rect 101178 120783 101234 120792
rect 101192 120750 101220 120783
rect 101180 120744 101232 120750
rect 101180 120686 101232 120692
rect 101088 120608 101140 120614
rect 101088 120550 101140 120556
rect 101284 120546 101312 122551
rect 135220 122522 135272 122528
rect 135218 122480 135274 122489
rect 135218 122415 135274 122424
rect 135232 122246 135260 122415
rect 135220 122240 135272 122246
rect 135220 122182 135272 122188
rect 137440 121974 137468 123610
rect 137428 121968 137480 121974
rect 134850 121936 134906 121945
rect 137428 121910 137480 121916
rect 134850 121871 134906 121880
rect 134666 121392 134722 121401
rect 134666 121327 134722 121336
rect 134680 120750 134708 121327
rect 134864 120818 134892 121871
rect 134852 120812 134904 120818
rect 134852 120754 134904 120760
rect 137336 120812 137388 120818
rect 137336 120754 137388 120760
rect 134668 120744 134720 120750
rect 134668 120686 134720 120692
rect 135402 120712 135458 120721
rect 135402 120647 135404 120656
rect 135456 120647 135458 120656
rect 136876 120676 136928 120682
rect 135404 120618 135456 120624
rect 136876 120618 136928 120624
rect 101272 120540 101324 120546
rect 101272 120482 101324 120488
rect 134298 120168 134354 120177
rect 134298 120103 134300 120112
rect 134352 120103 134354 120112
rect 134300 120074 134352 120080
rect 101086 119760 101142 119769
rect 101086 119695 101142 119704
rect 101100 119390 101128 119695
rect 135402 119624 135458 119633
rect 135402 119559 135404 119568
rect 135456 119559 135458 119568
rect 135404 119530 135456 119536
rect 101088 119384 101140 119390
rect 100994 119352 101050 119361
rect 101088 119326 101140 119332
rect 100994 119287 100996 119296
rect 101048 119287 101050 119296
rect 100996 119258 101048 119264
rect 136888 119118 136916 120618
rect 136968 120132 137020 120138
rect 136968 120074 137020 120080
rect 136876 119112 136928 119118
rect 136876 119054 136928 119060
rect 134850 118944 134906 118953
rect 134850 118879 134906 118888
rect 101086 118536 101142 118545
rect 101086 118471 101142 118480
rect 100994 117992 101050 118001
rect 101100 117962 101128 118471
rect 134482 118400 134538 118409
rect 134482 118335 134538 118344
rect 134496 118234 134524 118335
rect 134484 118228 134536 118234
rect 134484 118170 134536 118176
rect 134864 117962 134892 118879
rect 100994 117927 101050 117936
rect 101088 117956 101140 117962
rect 101008 117894 101036 117927
rect 101088 117898 101140 117904
rect 134852 117956 134904 117962
rect 134852 117898 134904 117904
rect 100996 117888 101048 117894
rect 100996 117830 101048 117836
rect 134850 117856 134906 117865
rect 136980 117826 137008 120074
rect 137348 119254 137376 120754
rect 137336 119248 137388 119254
rect 137336 119190 137388 119196
rect 137428 117956 137480 117962
rect 137428 117898 137480 117904
rect 134850 117791 134906 117800
rect 136968 117820 137020 117826
rect 101178 117448 101234 117457
rect 101178 117383 101234 117392
rect 101086 116768 101142 116777
rect 101086 116703 101142 116712
rect 100994 116632 101050 116641
rect 101100 116602 101128 116703
rect 100994 116567 101050 116576
rect 101088 116596 101140 116602
rect 101008 116534 101036 116567
rect 101088 116538 101140 116544
rect 100996 116528 101048 116534
rect 100996 116470 101048 116476
rect 101192 116466 101220 117383
rect 134758 116632 134814 116641
rect 134758 116567 134814 116576
rect 101180 116460 101232 116466
rect 101180 116402 101232 116408
rect 101086 115680 101142 115689
rect 101086 115615 101142 115624
rect 100994 115272 101050 115281
rect 101100 115242 101128 115615
rect 100994 115207 101050 115216
rect 101088 115236 101140 115242
rect 101008 115174 101036 115207
rect 101088 115178 101140 115184
rect 100996 115168 101048 115174
rect 100996 115110 101048 115116
rect 102006 114456 102062 114465
rect 102006 114391 102062 114400
rect 101638 113912 101694 113921
rect 101638 113847 101694 113856
rect 100994 112552 101050 112561
rect 100994 112487 101050 112496
rect 101008 112386 101036 112487
rect 100996 112380 101048 112386
rect 100996 112322 101048 112328
rect 99524 110476 99576 110482
rect 99524 110418 99576 110424
rect 99432 110340 99484 110346
rect 99432 110282 99484 110288
rect 99248 109864 99300 109870
rect 99248 109806 99300 109812
rect 99156 109796 99208 109802
rect 99156 109738 99208 109744
rect 99064 109728 99116 109734
rect 99064 109670 99116 109676
rect 98972 109660 99024 109666
rect 98972 109602 99024 109608
rect 98984 91209 99012 109602
rect 99076 92433 99104 109670
rect 99168 94337 99196 109738
rect 99260 95561 99288 109806
rect 99340 109592 99392 109598
rect 99340 109534 99392 109540
rect 99246 95552 99302 95561
rect 99246 95487 99302 95496
rect 99154 94328 99210 94337
rect 99154 94263 99210 94272
rect 99352 93657 99380 109534
rect 99444 97057 99472 110282
rect 99536 98553 99564 110418
rect 101652 102050 101680 113847
rect 101822 113776 101878 113785
rect 101822 113711 101878 113720
rect 101640 102044 101692 102050
rect 101640 101986 101692 101992
rect 101836 101982 101864 113711
rect 102020 102118 102048 114391
rect 104136 109666 104164 112932
rect 104596 109734 104624 112932
rect 104584 109728 104636 109734
rect 104584 109670 104636 109676
rect 104124 109660 104176 109666
rect 104124 109602 104176 109608
rect 105148 109598 105176 112932
rect 105700 109802 105728 112932
rect 106252 109870 106280 112932
rect 106804 110346 106832 112932
rect 107356 110482 107384 112932
rect 107344 110476 107396 110482
rect 107344 110418 107396 110424
rect 106792 110340 106844 110346
rect 106792 110282 106844 110288
rect 107908 110278 107936 112932
rect 108460 110958 108488 112932
rect 109012 110958 109040 112932
rect 108448 110952 108500 110958
rect 108448 110894 108500 110900
rect 109000 110952 109052 110958
rect 109000 110894 109052 110900
rect 108460 110278 108488 110894
rect 109564 110890 109592 112932
rect 109552 110884 109604 110890
rect 109552 110826 109604 110832
rect 107896 110272 107948 110278
rect 107896 110214 107948 110220
rect 108448 110272 108500 110278
rect 108448 110214 108500 110220
rect 106240 109864 106292 109870
rect 106240 109806 106292 109812
rect 105688 109796 105740 109802
rect 105688 109738 105740 109744
rect 105136 109592 105188 109598
rect 105136 109534 105188 109540
rect 102008 102112 102060 102118
rect 102008 102054 102060 102060
rect 101824 101976 101876 101982
rect 101824 101918 101876 101924
rect 110116 99740 110144 112932
rect 110668 110634 110696 112932
rect 110576 110606 110696 110634
rect 110576 99754 110604 110606
rect 111220 99754 111248 112932
rect 111772 102662 111800 112932
rect 111300 102656 111352 102662
rect 111300 102598 111352 102604
rect 111760 102656 111812 102662
rect 111760 102598 111812 102604
rect 110498 99726 110604 99754
rect 110866 99726 111248 99754
rect 111312 99740 111340 102598
rect 112324 102594 112352 112932
rect 112496 102656 112548 102662
rect 112496 102598 112548 102604
rect 111668 102588 111720 102594
rect 111668 102530 111720 102536
rect 112312 102588 112364 102594
rect 112312 102530 112364 102536
rect 111680 99740 111708 102530
rect 112036 101976 112088 101982
rect 112036 101918 112088 101924
rect 112048 99740 112076 101918
rect 112508 99740 112536 102598
rect 112876 101982 112904 112932
rect 113428 110634 113456 112932
rect 113336 110606 113456 110634
rect 113140 110544 113192 110550
rect 113140 110486 113192 110492
rect 113048 110204 113100 110210
rect 113048 110146 113100 110152
rect 112864 101976 112916 101982
rect 112864 101918 112916 101924
rect 113060 99754 113088 110146
rect 112890 99726 113088 99754
rect 113152 99754 113180 110486
rect 113336 102662 113364 110606
rect 113980 110210 114008 112932
rect 114532 110550 114560 112932
rect 115084 110634 115112 112932
rect 114716 110606 115112 110634
rect 114520 110544 114572 110550
rect 114520 110486 114572 110492
rect 114612 110544 114664 110550
rect 114612 110486 114664 110492
rect 113968 110204 114020 110210
rect 113968 110146 114020 110152
rect 113324 102656 113376 102662
rect 113324 102598 113376 102604
rect 113692 102656 113744 102662
rect 113692 102598 113744 102604
rect 113152 99726 113258 99754
rect 113704 99740 113732 102598
rect 114624 102594 114652 110486
rect 114716 102662 114744 110606
rect 115636 110550 115664 112932
rect 115624 110544 115676 110550
rect 115624 110486 115676 110492
rect 115992 110544 116044 110550
rect 115992 110486 116044 110492
rect 115716 110204 115768 110210
rect 115716 110146 115768 110152
rect 114704 102656 114756 102662
rect 114704 102598 114756 102604
rect 115624 102656 115676 102662
rect 115624 102598 115676 102604
rect 114060 102588 114112 102594
rect 114060 102530 114112 102536
rect 114612 102588 114664 102594
rect 114612 102530 114664 102536
rect 114888 102588 114940 102594
rect 114888 102530 114940 102536
rect 114072 99740 114100 102530
rect 114428 102248 114480 102254
rect 114428 102190 114480 102196
rect 114440 99740 114468 102190
rect 114900 99740 114928 102530
rect 115256 102520 115308 102526
rect 115256 102462 115308 102468
rect 115268 99740 115296 102462
rect 115636 99740 115664 102598
rect 115728 102594 115756 110146
rect 115808 110068 115860 110074
rect 115808 110010 115860 110016
rect 115716 102588 115768 102594
rect 115716 102530 115768 102536
rect 115820 99754 115848 110010
rect 115900 109728 115952 109734
rect 115900 109670 115952 109676
rect 115912 102662 115940 109670
rect 115900 102656 115952 102662
rect 115900 102598 115952 102604
rect 116004 102526 116032 110486
rect 115992 102520 116044 102526
rect 115992 102462 116044 102468
rect 116188 102254 116216 112932
rect 116740 110210 116768 112932
rect 117292 110550 117320 112932
rect 117280 110544 117332 110550
rect 117280 110486 117332 110492
rect 117464 110544 117516 110550
rect 117464 110486 117516 110492
rect 116728 110204 116780 110210
rect 116728 110146 116780 110152
rect 116176 102248 116228 102254
rect 116176 102190 116228 102196
rect 117476 101846 117504 110486
rect 117844 109734 117872 112932
rect 118304 110074 118332 112932
rect 118856 110550 118884 112932
rect 118844 110544 118896 110550
rect 118844 110486 118896 110492
rect 118292 110068 118344 110074
rect 118292 110010 118344 110016
rect 118936 109796 118988 109802
rect 118936 109738 118988 109744
rect 117832 109728 117884 109734
rect 117832 109670 117884 109676
rect 116452 101840 116504 101846
rect 116452 101782 116504 101788
rect 117464 101840 117516 101846
rect 117464 101782 117516 101788
rect 115820 99726 116110 99754
rect 116464 99740 116492 101782
rect 117648 101704 117700 101710
rect 117648 101646 117700 101652
rect 116820 101636 116872 101642
rect 116820 101578 116872 101584
rect 116832 99740 116860 101578
rect 117280 101432 117332 101438
rect 117280 101374 117332 101380
rect 117292 99740 117320 101374
rect 117660 99740 117688 101646
rect 118844 101568 118896 101574
rect 118844 101510 118896 101516
rect 118476 101500 118528 101506
rect 118476 101442 118528 101448
rect 118108 101364 118160 101370
rect 118108 101306 118160 101312
rect 118120 99740 118148 101306
rect 118488 99740 118516 101442
rect 118856 99740 118884 101510
rect 118948 101438 118976 109738
rect 119408 101642 119436 112932
rect 119764 109864 119816 109870
rect 119764 109806 119816 109812
rect 119580 109728 119632 109734
rect 119580 109670 119632 109676
rect 119396 101636 119448 101642
rect 119396 101578 119448 101584
rect 118936 101432 118988 101438
rect 118936 101374 118988 101380
rect 119304 101432 119356 101438
rect 119304 101374 119356 101380
rect 119316 99740 119344 101374
rect 119592 101370 119620 109670
rect 119672 102384 119724 102390
rect 119672 102326 119724 102332
rect 119580 101364 119632 101370
rect 119580 101306 119632 101312
rect 119684 99740 119712 102326
rect 119776 101506 119804 109806
rect 119960 109802 119988 112932
rect 119948 109796 120000 109802
rect 119948 109738 120000 109744
rect 119948 109660 120000 109666
rect 119948 109602 120000 109608
rect 119856 109592 119908 109598
rect 119856 109534 119908 109540
rect 119868 101710 119896 109534
rect 119856 101704 119908 101710
rect 119856 101646 119908 101652
rect 119960 101574 119988 109602
rect 120512 109598 120540 112932
rect 121064 109734 121092 112932
rect 121616 109870 121644 112932
rect 121604 109864 121656 109870
rect 121604 109806 121656 109812
rect 121052 109728 121104 109734
rect 121052 109670 121104 109676
rect 122168 109666 122196 112932
rect 122156 109660 122208 109666
rect 122156 109602 122208 109608
rect 122720 109598 122748 112932
rect 120500 109592 120552 109598
rect 120500 109534 120552 109540
rect 120960 109592 121012 109598
rect 120960 109534 121012 109540
rect 122708 109592 122760 109598
rect 122708 109534 122760 109540
rect 120500 102520 120552 102526
rect 120500 102462 120552 102468
rect 120040 102452 120092 102458
rect 120040 102394 120092 102400
rect 119948 101568 120000 101574
rect 119948 101510 120000 101516
rect 119764 101500 119816 101506
rect 119764 101442 119816 101448
rect 120052 99740 120080 102394
rect 120512 99740 120540 102462
rect 120868 101772 120920 101778
rect 120868 101714 120920 101720
rect 120880 99740 120908 101714
rect 120972 101438 121000 109534
rect 123272 102390 123300 112932
rect 123824 102458 123852 112932
rect 124376 102526 124404 112932
rect 124364 102520 124416 102526
rect 124364 102462 124416 102468
rect 123812 102452 123864 102458
rect 123812 102394 123864 102400
rect 123260 102384 123312 102390
rect 123260 102326 123312 102332
rect 122432 102248 122484 102254
rect 122432 102190 122484 102196
rect 121696 102180 121748 102186
rect 121696 102122 121748 102128
rect 121236 101976 121288 101982
rect 121236 101918 121288 101924
rect 120960 101432 121012 101438
rect 120960 101374 121012 101380
rect 121248 99740 121276 101918
rect 121708 99740 121736 102122
rect 122064 102044 122116 102050
rect 122064 101986 122116 101992
rect 122076 99740 122104 101986
rect 122444 99740 122472 102190
rect 122892 102112 122944 102118
rect 122892 102054 122944 102060
rect 122904 99740 122932 102054
rect 124456 101840 124508 101846
rect 124456 101782 124508 101788
rect 123260 101704 123312 101710
rect 123260 101646 123312 101652
rect 123272 99740 123300 101646
rect 123628 101636 123680 101642
rect 123628 101578 123680 101584
rect 123640 99740 123668 101578
rect 124088 101500 124140 101506
rect 124088 101442 124140 101448
rect 124100 99740 124128 101442
rect 124468 99740 124496 101782
rect 124928 101778 124956 112932
rect 125480 101982 125508 112932
rect 126032 102186 126060 112932
rect 126584 109954 126612 112932
rect 126124 109926 126612 109954
rect 126020 102180 126072 102186
rect 126020 102122 126072 102128
rect 126124 102050 126152 109926
rect 126664 109796 126716 109802
rect 126664 109738 126716 109744
rect 126572 109660 126624 109666
rect 126572 109602 126624 109608
rect 126480 109592 126532 109598
rect 126480 109534 126532 109540
rect 126112 102044 126164 102050
rect 126112 101986 126164 101992
rect 125468 101976 125520 101982
rect 125468 101918 125520 101924
rect 124916 101772 124968 101778
rect 124916 101714 124968 101720
rect 126492 101710 126520 109534
rect 126480 101704 126532 101710
rect 126480 101646 126532 101652
rect 126584 101642 126612 109602
rect 126572 101636 126624 101642
rect 126572 101578 126624 101584
rect 124824 101568 124876 101574
rect 124824 101510 124876 101516
rect 124836 99740 124864 101510
rect 126676 101506 126704 109738
rect 127136 102254 127164 112932
rect 127124 102248 127176 102254
rect 127124 102190 127176 102196
rect 127688 102118 127716 112932
rect 128240 109598 128268 112932
rect 128792 109666 128820 112932
rect 129344 109802 129372 112932
rect 129332 109796 129384 109802
rect 129332 109738 129384 109744
rect 128780 109660 128832 109666
rect 128780 109602 128832 109608
rect 129332 109660 129384 109666
rect 129332 109602 129384 109608
rect 128228 109592 128280 109598
rect 128228 109534 128280 109540
rect 129240 109592 129292 109598
rect 129240 109534 129292 109540
rect 127676 102112 127728 102118
rect 127676 102054 127728 102060
rect 129252 101574 129280 109534
rect 129240 101568 129292 101574
rect 129240 101510 129292 101516
rect 126664 101500 126716 101506
rect 126664 101442 126716 101448
rect 125652 101432 125704 101438
rect 125652 101374 125704 101380
rect 125284 101364 125336 101370
rect 125284 101306 125336 101312
rect 125296 99740 125324 101306
rect 125664 99740 125692 101374
rect 129344 101370 129372 109602
rect 129896 101846 129924 112932
rect 129976 111632 130028 111638
rect 129976 111574 130028 111580
rect 129988 110958 130016 111574
rect 129976 110952 130028 110958
rect 129976 110894 130028 110900
rect 130448 109598 130476 112932
rect 131000 109666 131028 112932
rect 130988 109660 131040 109666
rect 130988 109602 131040 109608
rect 130436 109592 130488 109598
rect 130436 109534 130488 109540
rect 129884 101840 129936 101846
rect 129884 101782 129936 101788
rect 131552 101438 131580 112932
rect 133380 110272 133432 110278
rect 133380 110214 133432 110220
rect 131540 101432 131592 101438
rect 131540 101374 131592 101380
rect 129332 101364 129384 101370
rect 129332 101306 129384 101312
rect 99522 98544 99578 98553
rect 99522 98479 99578 98488
rect 106790 98544 106846 98553
rect 106790 98479 106846 98488
rect 106804 97222 106832 98479
rect 106792 97216 106844 97222
rect 106792 97158 106844 97164
rect 99430 97048 99486 97057
rect 99430 96983 99486 96992
rect 106790 96232 106846 96241
rect 106790 96167 106846 96176
rect 106804 95862 106832 96167
rect 99524 95856 99576 95862
rect 99524 95798 99576 95804
rect 106792 95856 106844 95862
rect 106792 95798 106844 95804
rect 99338 93648 99394 93657
rect 99338 93583 99394 93592
rect 99062 92424 99118 92433
rect 99062 92359 99118 92368
rect 98970 91200 99026 91209
rect 98970 91135 99026 91144
rect 99536 88761 99564 95798
rect 106514 93920 106570 93929
rect 106514 93855 106570 93864
rect 106528 93074 106556 93855
rect 106516 93068 106568 93074
rect 106516 93010 106568 93016
rect 106790 91472 106846 91481
rect 106790 91407 106846 91416
rect 106804 90286 106832 91407
rect 105044 90280 105096 90286
rect 105044 90222 105096 90228
rect 106792 90280 106844 90286
rect 106792 90222 106844 90228
rect 104952 88920 105004 88926
rect 104952 88862 105004 88868
rect 99522 88752 99578 88761
rect 99522 88687 99578 88696
rect 99522 85352 99578 85361
rect 99522 85287 99578 85296
rect 99536 85254 99564 85287
rect 99524 85248 99576 85254
rect 99524 85190 99576 85196
rect 99432 84704 99484 84710
rect 99432 84646 99484 84652
rect 99522 84672 99578 84681
rect 99444 84001 99472 84646
rect 104964 84642 104992 88862
rect 105056 85254 105084 90222
rect 128502 89840 128558 89849
rect 128502 89775 128558 89784
rect 106790 89160 106846 89169
rect 106790 89095 106846 89104
rect 106804 88926 106832 89095
rect 128516 88926 128544 89775
rect 106792 88920 106844 88926
rect 106792 88862 106844 88868
rect 128504 88920 128556 88926
rect 128504 88862 128556 88868
rect 132000 88920 132052 88926
rect 132000 88862 132052 88868
rect 106790 86848 106846 86857
rect 106790 86783 106846 86792
rect 105044 85248 105096 85254
rect 105044 85190 105096 85196
rect 106804 84710 106832 86783
rect 106792 84704 106844 84710
rect 106792 84646 106844 84652
rect 99522 84607 99524 84616
rect 99576 84607 99578 84616
rect 104952 84636 105004 84642
rect 99524 84578 99576 84584
rect 104952 84578 105004 84584
rect 107802 84400 107858 84409
rect 107802 84335 107858 84344
rect 99430 83992 99486 84001
rect 99430 83927 99486 83936
rect 107816 83350 107844 84335
rect 99524 83344 99576 83350
rect 99524 83286 99576 83292
rect 107804 83344 107856 83350
rect 107804 83286 107856 83292
rect 99536 82777 99564 83286
rect 99522 82768 99578 82777
rect 99522 82703 99578 82712
rect 106792 82120 106844 82126
rect 106790 82088 106792 82097
rect 106844 82088 106846 82097
rect 106790 82023 106846 82032
rect 99524 81984 99576 81990
rect 99524 81926 99576 81932
rect 99536 81553 99564 81926
rect 99522 81544 99578 81553
rect 99522 81479 99578 81488
rect 132012 80562 132040 88862
rect 132000 80556 132052 80562
rect 132000 80498 132052 80504
rect 99524 79876 99576 79882
rect 99524 79818 99576 79824
rect 106792 79876 106844 79882
rect 106792 79818 106844 79824
rect 99536 79785 99564 79818
rect 106804 79785 106832 79818
rect 99522 79776 99578 79785
rect 99522 79711 99578 79720
rect 106790 79776 106846 79785
rect 106790 79711 106846 79720
rect 99522 78008 99578 78017
rect 99522 77943 99578 77952
rect 99536 77910 99564 77943
rect 99524 77904 99576 77910
rect 99524 77846 99576 77852
rect 106516 77904 106568 77910
rect 106516 77846 106568 77852
rect 106528 77473 106556 77846
rect 106514 77464 106570 77473
rect 106514 77399 106570 77408
rect 99522 76784 99578 76793
rect 99522 76719 99578 76728
rect 99536 76482 99564 76719
rect 99524 76476 99576 76482
rect 99524 76418 99576 76424
rect 100996 76476 101048 76482
rect 100996 76418 101048 76424
rect 101008 75054 101036 76418
rect 100996 75048 101048 75054
rect 106792 75048 106844 75054
rect 100996 74990 101048 74996
rect 106790 75016 106792 75025
rect 106844 75016 106846 75025
rect 106790 74951 106846 74960
rect 100996 74912 101048 74918
rect 100996 74854 101048 74860
rect 99430 74336 99486 74345
rect 99430 74271 99486 74280
rect 99444 73762 99472 74271
rect 99524 73892 99576 73898
rect 99524 73834 99576 73840
rect 99536 73801 99564 73834
rect 99522 73792 99578 73801
rect 99432 73756 99484 73762
rect 99522 73727 99578 73736
rect 99432 73698 99484 73704
rect 101008 73694 101036 74854
rect 105136 73892 105188 73898
rect 105136 73834 105188 73840
rect 100996 73688 101048 73694
rect 100996 73630 101048 73636
rect 99522 72568 99578 72577
rect 99522 72503 99578 72512
rect 99536 72402 99564 72503
rect 99524 72396 99576 72402
rect 99524 72338 99576 72344
rect 99522 71072 99578 71081
rect 99522 71007 99524 71016
rect 99576 71007 99578 71016
rect 104492 71036 104544 71042
rect 99524 70978 99576 70984
rect 104492 70978 104544 70984
rect 99522 69848 99578 69857
rect 99522 69783 99578 69792
rect 99536 69614 99564 69783
rect 99524 69608 99576 69614
rect 99524 69550 99576 69556
rect 104400 69608 104452 69614
rect 104400 69550 104452 69556
rect 98970 68352 99026 68361
rect 98970 68287 99026 68296
rect 98880 58456 98932 58462
rect 98880 58398 98932 58404
rect 92532 57912 92584 57918
rect 92532 57854 92584 57860
rect 72568 57844 72620 57850
rect 72568 57786 72620 57792
rect 98984 49554 99012 68287
rect 99062 67128 99118 67137
rect 99062 67063 99118 67072
rect 99076 49622 99104 67063
rect 99154 65904 99210 65913
rect 99154 65839 99210 65848
rect 99168 49690 99196 65839
rect 99246 64680 99302 64689
rect 99246 64615 99302 64624
rect 99260 49826 99288 64615
rect 99522 63456 99578 63465
rect 99522 63391 99578 63400
rect 99338 62776 99394 62785
rect 99338 62711 99394 62720
rect 99352 50166 99380 62711
rect 99536 61674 99564 63391
rect 99536 61646 99656 61674
rect 99522 61552 99578 61561
rect 99522 61487 99578 61496
rect 99536 61386 99564 61487
rect 99524 61380 99576 61386
rect 99524 61322 99576 61328
rect 99628 61266 99656 61646
rect 99536 61238 99656 61266
rect 104412 61250 104440 69550
rect 104504 63698 104532 70978
rect 105148 68186 105176 73834
rect 106700 73756 106752 73762
rect 106700 73698 106752 73704
rect 106516 72396 106568 72402
rect 106516 72338 106568 72344
rect 105136 68180 105188 68186
rect 105136 68122 105188 68128
rect 106528 65641 106556 72338
rect 106712 70401 106740 73698
rect 106792 73688 106844 73694
rect 106792 73630 106844 73636
rect 106804 72713 106832 73630
rect 106790 72704 106846 72713
rect 106790 72639 106846 72648
rect 106698 70392 106754 70401
rect 106698 70327 106754 70336
rect 133392 70226 133420 110214
rect 134772 102118 134800 116567
rect 134864 116534 134892 117791
rect 136968 117762 137020 117768
rect 134942 117312 134998 117321
rect 134942 117247 134998 117256
rect 134852 116528 134904 116534
rect 134852 116470 134904 116476
rect 134850 116088 134906 116097
rect 134850 116023 134906 116032
rect 134864 102186 134892 116023
rect 134852 102180 134904 102186
rect 134852 102122 134904 102128
rect 134760 102112 134812 102118
rect 134760 102054 134812 102060
rect 134956 102050 134984 117247
rect 137440 116398 137468 117898
rect 137428 116392 137480 116398
rect 137428 116334 137480 116340
rect 135034 115544 135090 115553
rect 135034 115479 135090 115488
rect 135048 102254 135076 115479
rect 135126 114864 135182 114873
rect 135126 114799 135182 114808
rect 135140 102390 135168 114799
rect 135310 114320 135366 114329
rect 135310 114255 135366 114264
rect 135218 113232 135274 113241
rect 135218 113167 135274 113176
rect 135128 102384 135180 102390
rect 135128 102326 135180 102332
rect 135036 102248 135088 102254
rect 135036 102190 135088 102196
rect 134944 102044 134996 102050
rect 134944 101986 134996 101992
rect 135232 101370 135260 113167
rect 135324 101982 135352 114255
rect 135402 113776 135458 113785
rect 135402 113711 135404 113720
rect 135456 113711 135458 113720
rect 135404 113682 135456 113688
rect 137532 110958 137560 156687
rect 182782 155528 182838 155537
rect 182782 155463 182784 155472
rect 182836 155463 182838 155472
rect 182784 155434 182836 155440
rect 143250 153854 143724 153882
rect 143592 140056 143644 140062
rect 143592 139998 143644 140004
rect 143316 139988 143368 139994
rect 143316 139930 143368 139936
rect 139820 138764 139872 138770
rect 139820 138706 139872 138712
rect 139636 138628 139688 138634
rect 139636 138570 139688 138576
rect 139648 137070 139676 138570
rect 139728 137404 139780 137410
rect 139728 137346 139780 137352
rect 139636 137064 139688 137070
rect 139636 137006 139688 137012
rect 139740 136662 139768 137346
rect 139832 137002 139860 138706
rect 143328 138265 143356 139930
rect 143604 138537 143632 139998
rect 143590 138528 143646 138537
rect 143590 138463 143646 138472
rect 143314 138256 143370 138265
rect 143314 138191 143370 138200
rect 143408 137200 143460 137206
rect 143408 137142 143460 137148
rect 143590 137168 143646 137177
rect 139820 136996 139872 137002
rect 139820 136938 139872 136944
rect 143132 136996 143184 137002
rect 143132 136938 143184 136944
rect 143144 136905 143172 136938
rect 143130 136896 143186 136905
rect 143130 136831 143186 136840
rect 139728 136656 139780 136662
rect 139728 136598 139780 136604
rect 143316 135976 143368 135982
rect 143316 135918 143368 135924
rect 143224 135840 143276 135846
rect 143224 135782 143276 135788
rect 139636 134548 139688 134554
rect 139636 134490 139688 134496
rect 139648 133806 139676 134490
rect 143236 134049 143264 135782
rect 143328 135273 143356 135918
rect 143420 135817 143448 137142
rect 143590 137103 143646 137112
rect 143604 137070 143632 137103
rect 143592 137064 143644 137070
rect 143592 137006 143644 137012
rect 143500 136656 143552 136662
rect 143500 136598 143552 136604
rect 143512 136361 143540 136598
rect 143498 136352 143554 136361
rect 143498 136287 143554 136296
rect 143592 135908 143644 135914
rect 143592 135850 143644 135856
rect 143406 135808 143462 135817
rect 143406 135743 143462 135752
rect 143314 135264 143370 135273
rect 143314 135199 143370 135208
rect 143604 134321 143632 135850
rect 143590 134312 143646 134321
rect 143590 134247 143646 134256
rect 143222 134040 143278 134049
rect 143222 133975 143278 133984
rect 139636 133800 139688 133806
rect 139636 133742 139688 133748
rect 142948 133800 143000 133806
rect 142948 133742 143000 133748
rect 142960 133369 142988 133742
rect 142946 133360 143002 133369
rect 142946 133295 143002 133304
rect 138164 133120 138216 133126
rect 138164 133062 138216 133068
rect 138072 132032 138124 132038
rect 138072 131974 138124 131980
rect 137612 130604 137664 130610
rect 137612 130546 137664 130552
rect 137624 128774 137652 130546
rect 138084 130270 138112 131974
rect 138176 131562 138204 133062
rect 143224 132984 143276 132990
rect 143224 132926 143276 132932
rect 143236 132281 143264 132926
rect 143592 132848 143644 132854
rect 143590 132816 143592 132825
rect 143644 132816 143646 132825
rect 143590 132751 143646 132760
rect 143222 132272 143278 132281
rect 143222 132207 143278 132216
rect 142488 131624 142540 131630
rect 142488 131566 142540 131572
rect 138164 131556 138216 131562
rect 138164 131498 138216 131504
rect 142500 131057 142528 131566
rect 143592 131556 143644 131562
rect 143592 131498 143644 131504
rect 143604 131465 143632 131498
rect 143590 131456 143646 131465
rect 143590 131391 143646 131400
rect 142486 131048 142542 131057
rect 142486 130983 142542 130992
rect 138072 130264 138124 130270
rect 143592 130264 143644 130270
rect 138072 130206 138124 130212
rect 143590 130232 143592 130241
rect 143644 130232 143646 130241
rect 143040 130196 143092 130202
rect 143590 130167 143646 130176
rect 143040 130138 143092 130144
rect 143052 129969 143080 130138
rect 143038 129960 143094 129969
rect 143038 129895 143094 129904
rect 137704 129380 137756 129386
rect 137704 129322 137756 129328
rect 137612 128768 137664 128774
rect 137612 128710 137664 128716
rect 137612 127748 137664 127754
rect 137612 127690 137664 127696
rect 137624 126122 137652 127690
rect 137716 127414 137744 129322
rect 143132 128904 143184 128910
rect 142762 128872 142818 128881
rect 143132 128846 143184 128852
rect 142762 128807 142764 128816
rect 142816 128807 142818 128816
rect 142764 128778 142816 128784
rect 143144 128065 143172 128846
rect 143592 128768 143644 128774
rect 143590 128736 143592 128745
rect 143644 128736 143646 128745
rect 143590 128671 143646 128680
rect 143130 128056 143186 128065
rect 143130 127991 143186 128000
rect 143316 127476 143368 127482
rect 143316 127418 143368 127424
rect 137704 127408 137756 127414
rect 142488 127408 142540 127414
rect 137704 127350 137756 127356
rect 142486 127376 142488 127385
rect 142540 127376 142542 127385
rect 142486 127311 142542 127320
rect 143328 126977 143356 127418
rect 143314 126968 143370 126977
rect 143314 126903 143370 126912
rect 137612 126116 137664 126122
rect 137612 126058 137664 126064
rect 143500 126116 143552 126122
rect 143500 126058 143552 126064
rect 143512 125617 143540 126058
rect 143592 126048 143644 126054
rect 143590 126016 143592 126025
rect 143644 126016 143646 126025
rect 143590 125951 143646 125960
rect 143498 125608 143554 125617
rect 143498 125543 143554 125552
rect 137612 125436 137664 125442
rect 137612 125378 137664 125384
rect 137624 123334 137652 125378
rect 142764 124824 142816 124830
rect 142764 124766 142816 124772
rect 142488 124416 142540 124422
rect 142486 124384 142488 124393
rect 142540 124384 142542 124393
rect 142486 124319 142542 124328
rect 142776 123985 142804 124766
rect 143592 124756 143644 124762
rect 143592 124698 143644 124704
rect 143604 124665 143632 124698
rect 143590 124656 143646 124665
rect 143590 124591 143646 124600
rect 142762 123976 142818 123985
rect 142762 123911 142818 123920
rect 138164 123396 138216 123402
rect 138164 123338 138216 123344
rect 137612 123328 137664 123334
rect 137612 123270 137664 123276
rect 137888 122580 137940 122586
rect 137888 122522 137940 122528
rect 137796 122240 137848 122246
rect 137796 122182 137848 122188
rect 137612 120744 137664 120750
rect 137612 120686 137664 120692
rect 137624 119186 137652 120686
rect 137808 120546 137836 122182
rect 137900 120614 137928 122522
rect 138176 121906 138204 123338
rect 143592 123328 143644 123334
rect 143590 123296 143592 123305
rect 143644 123296 143646 123305
rect 143590 123231 143646 123240
rect 143592 122852 143644 122858
rect 143592 122794 143644 122800
rect 143604 122489 143632 122794
rect 143590 122480 143646 122489
rect 143590 122415 143646 122424
rect 142764 121968 142816 121974
rect 142764 121910 142816 121916
rect 138164 121900 138216 121906
rect 138164 121842 138216 121848
rect 142776 121537 142804 121910
rect 143040 121900 143092 121906
rect 143040 121842 143092 121848
rect 143052 121809 143080 121842
rect 143038 121800 143094 121809
rect 143038 121735 143094 121744
rect 142762 121528 142818 121537
rect 142762 121463 142818 121472
rect 137888 120608 137940 120614
rect 142948 120608 143000 120614
rect 137888 120550 137940 120556
rect 142946 120576 142948 120585
rect 143000 120576 143002 120585
rect 137796 120540 137848 120546
rect 142946 120511 143002 120520
rect 143592 120540 143644 120546
rect 137796 120482 137848 120488
rect 143592 120482 143644 120488
rect 143604 120313 143632 120482
rect 143590 120304 143646 120313
rect 143590 120239 143646 120248
rect 137704 119588 137756 119594
rect 137704 119530 137756 119536
rect 137612 119180 137664 119186
rect 137612 119122 137664 119128
rect 137612 118228 137664 118234
rect 137612 118170 137664 118176
rect 137624 116330 137652 118170
rect 137716 117758 137744 119530
rect 143592 119248 143644 119254
rect 143590 119216 143592 119225
rect 143644 119216 143646 119225
rect 143040 119180 143092 119186
rect 143590 119151 143646 119160
rect 143040 119122 143092 119128
rect 143052 118953 143080 119122
rect 143316 119112 143368 119118
rect 143316 119054 143368 119060
rect 143038 118944 143094 118953
rect 143038 118879 143094 118888
rect 143328 118545 143356 119054
rect 143314 118536 143370 118545
rect 143314 118471 143370 118480
rect 142580 117820 142632 117826
rect 142580 117762 142632 117768
rect 137704 117752 137756 117758
rect 142592 117729 142620 117762
rect 143224 117752 143276 117758
rect 137704 117694 137756 117700
rect 142578 117720 142634 117729
rect 143224 117694 143276 117700
rect 142578 117655 142634 117664
rect 143236 117321 143264 117694
rect 143222 117312 143278 117321
rect 143222 117247 143278 117256
rect 142764 116460 142816 116466
rect 142764 116402 142816 116408
rect 137612 116324 137664 116330
rect 137612 116266 137664 116272
rect 142776 115553 142804 116402
rect 142948 116392 143000 116398
rect 142946 116360 142948 116369
rect 143000 116360 143002 116369
rect 142946 116295 143002 116304
rect 143592 116324 143644 116330
rect 143592 116266 143644 116272
rect 143604 116097 143632 116266
rect 143590 116088 143646 116097
rect 143590 116023 143646 116032
rect 142762 115544 142818 115553
rect 142762 115479 142818 115488
rect 141568 113740 141620 113746
rect 141568 113682 141620 113688
rect 137520 110952 137572 110958
rect 137520 110894 137572 110900
rect 137532 110278 137560 110894
rect 137520 110272 137572 110278
rect 137520 110214 137572 110220
rect 135312 101976 135364 101982
rect 135312 101918 135364 101924
rect 135220 101364 135272 101370
rect 135220 101306 135272 101312
rect 140464 101364 140516 101370
rect 140464 101306 140516 101312
rect 140476 99740 140504 101306
rect 141580 99740 141608 113682
rect 143696 102322 143724 153854
rect 156576 151758 156604 153868
rect 156564 151752 156616 151758
rect 156564 151694 156616 151700
rect 163200 151690 163228 153868
rect 163188 151684 163240 151690
rect 163188 151626 163240 151632
rect 169916 142510 169944 153868
rect 183072 143462 183100 162807
rect 187948 162026 187976 166450
rect 190052 165012 190104 165018
rect 190052 164954 190104 164960
rect 189960 163448 190012 163454
rect 189960 163390 190012 163396
rect 187936 162020 187988 162026
rect 187936 161962 187988 161968
rect 183150 161648 183206 161657
rect 183150 161583 183206 161592
rect 183060 143456 183112 143462
rect 183060 143398 183112 143404
rect 183164 143394 183192 161583
rect 183242 160424 183298 160433
rect 183242 160359 183298 160368
rect 183256 143530 183284 160359
rect 183518 159200 183574 159209
rect 183518 159135 183574 159144
rect 183334 157976 183390 157985
rect 183334 157911 183390 157920
rect 183348 143870 183376 157911
rect 183426 156752 183482 156761
rect 183426 156687 183482 156696
rect 183440 144006 183468 156687
rect 183428 144000 183480 144006
rect 183428 143942 183480 143948
rect 183532 143938 183560 159135
rect 189972 156761 190000 163390
rect 190064 158801 190092 164954
rect 191352 164785 191380 167538
rect 191904 166825 191932 168898
rect 191984 168888 192036 168894
rect 191984 168830 192036 168836
rect 191996 168729 192024 168830
rect 191982 168720 192038 168729
rect 191982 168655 192038 168664
rect 191890 166816 191946 166825
rect 191890 166751 191946 166760
rect 191338 164776 191394 164785
rect 191338 164711 191394 164720
rect 211762 163824 211818 163833
rect 211762 163759 211818 163768
rect 211776 163658 211804 163759
rect 211764 163652 211816 163658
rect 211764 163594 211816 163600
rect 191524 163040 191576 163046
rect 191524 162982 191576 162988
rect 191536 162745 191564 162982
rect 191522 162736 191578 162745
rect 191522 162671 191578 162680
rect 191984 162020 192036 162026
rect 191984 161962 192036 161968
rect 191996 160841 192024 161962
rect 191982 160832 192038 160841
rect 191982 160767 192038 160776
rect 190050 158792 190106 158801
rect 190050 158727 190106 158736
rect 189958 156752 190014 156761
rect 189958 156687 190014 156696
rect 188028 155492 188080 155498
rect 188028 155434 188080 155440
rect 183610 154440 183666 154449
rect 183610 154375 183666 154384
rect 183624 144074 183652 154375
rect 183612 144068 183664 144074
rect 183612 144010 183664 144016
rect 187936 144068 187988 144074
rect 187936 144010 187988 144016
rect 183520 143932 183572 143938
rect 183520 143874 183572 143880
rect 183336 143864 183388 143870
rect 183336 143806 183388 143812
rect 183244 143524 183296 143530
rect 183244 143466 183296 143472
rect 183152 143388 183204 143394
rect 183152 143330 183204 143336
rect 167696 142504 167748 142510
rect 167696 142446 167748 142452
rect 169904 142504 169956 142510
rect 169904 142446 169956 142452
rect 167708 138786 167736 142446
rect 187948 140826 187976 144010
rect 188040 140962 188068 155434
rect 191982 154848 192038 154857
rect 191982 154783 192038 154792
rect 189408 144000 189460 144006
rect 189408 143942 189460 143948
rect 188040 140934 188528 140962
rect 188500 140826 188528 140934
rect 187948 140798 188238 140826
rect 188500 140798 188790 140826
rect 189420 140690 189448 143942
rect 190052 143932 190104 143938
rect 190052 143874 190104 143880
rect 189500 143864 189552 143870
rect 189500 143806 189552 143812
rect 189512 140826 189540 143806
rect 190064 140826 190092 143874
rect 190788 143524 190840 143530
rect 190788 143466 190840 143472
rect 190800 140826 190828 143466
rect 191996 143394 192024 154783
rect 199646 153990 200028 154018
rect 193364 151072 193416 151078
rect 193364 151014 193416 151020
rect 193272 151004 193324 151010
rect 193272 150946 193324 150952
rect 193284 143666 193312 150946
rect 192996 143660 193048 143666
rect 192996 143602 193048 143608
rect 193272 143660 193324 143666
rect 193272 143602 193324 143608
rect 192076 143456 192128 143462
rect 192076 143398 192128 143404
rect 191340 143388 191392 143394
rect 191340 143330 191392 143336
rect 191984 143388 192036 143394
rect 191984 143330 192036 143336
rect 191352 140826 191380 143330
rect 192088 140826 192116 143398
rect 189512 140798 189894 140826
rect 190064 140798 190446 140826
rect 190800 140798 191090 140826
rect 191352 140798 191642 140826
rect 192088 140798 192194 140826
rect 193008 140690 193036 143602
rect 193376 140690 193404 151014
rect 194112 151010 194140 153868
rect 194480 151078 194508 153868
rect 194468 151072 194520 151078
rect 194468 151014 194520 151020
rect 194100 151004 194152 151010
rect 194848 150992 194876 153868
rect 194100 150946 194152 150952
rect 194664 150964 194876 150992
rect 194940 153854 195322 153882
rect 195400 153854 195690 153882
rect 194664 143666 194692 150964
rect 194940 150890 194968 153854
rect 194756 150862 194968 150890
rect 194192 143660 194244 143666
rect 194192 143602 194244 143608
rect 194652 143660 194704 143666
rect 194652 143602 194704 143608
rect 194204 140690 194232 143602
rect 194756 140690 194784 150862
rect 195400 150346 195428 153854
rect 196044 151010 196072 153868
rect 196228 153854 196518 153882
rect 196228 152352 196256 153854
rect 196136 152324 196256 152352
rect 195480 151004 195532 151010
rect 195480 150946 195532 150952
rect 196032 151004 196084 151010
rect 196032 150946 196084 150952
rect 195124 150318 195428 150346
rect 195124 140690 195152 150318
rect 195492 150210 195520 150946
rect 195216 150182 195520 150210
rect 195216 140826 195244 150182
rect 196136 140962 196164 152324
rect 196216 152228 196268 152234
rect 196216 152170 196268 152176
rect 196228 148358 196256 152170
rect 196872 151010 196900 153868
rect 197240 152234 197268 153868
rect 197596 152364 197648 152370
rect 197596 152306 197648 152312
rect 197228 152228 197280 152234
rect 197228 152170 197280 152176
rect 196308 151004 196360 151010
rect 196308 150946 196360 150952
rect 196860 151004 196912 151010
rect 196860 150946 196912 150952
rect 196216 148352 196268 148358
rect 196216 148294 196268 148300
rect 196320 140962 196348 150946
rect 197044 148352 197096 148358
rect 197044 148294 197096 148300
rect 196136 140934 196256 140962
rect 196320 140934 196532 140962
rect 195216 140798 195598 140826
rect 196228 140690 196256 140934
rect 196504 140826 196532 140934
rect 197056 140826 197084 148294
rect 197608 146182 197636 152306
rect 197596 146176 197648 146182
rect 197596 146118 197648 146124
rect 197700 140826 197728 153868
rect 198068 152370 198096 153868
rect 198056 152364 198108 152370
rect 198056 152306 198108 152312
rect 198148 146176 198200 146182
rect 198148 146118 198200 146124
rect 198160 140826 198188 146118
rect 198436 144074 198464 153868
rect 198424 144068 198476 144074
rect 198424 144010 198476 144016
rect 198896 144006 198924 153868
rect 199264 146130 199292 153868
rect 200000 152386 200028 153990
rect 200106 153854 200304 153882
rect 200000 152358 200212 152386
rect 199264 146102 199752 146130
rect 199068 144068 199120 144074
rect 199068 144010 199120 144016
rect 198884 144000 198936 144006
rect 198884 143942 198936 143948
rect 196504 140798 196794 140826
rect 197056 140798 197346 140826
rect 197700 140798 197898 140826
rect 198160 140798 198450 140826
rect 199080 140690 199108 144010
rect 199252 144000 199304 144006
rect 199252 143942 199304 143948
rect 199264 140826 199292 143942
rect 199724 140826 199752 146102
rect 200184 142730 200212 152358
rect 200276 142850 200304 153854
rect 200460 152370 200488 153868
rect 200448 152364 200500 152370
rect 200448 152306 200500 152312
rect 200828 151282 200856 153868
rect 201302 153854 201500 153882
rect 201184 152364 201236 152370
rect 201184 152306 201236 152312
rect 201368 152364 201420 152370
rect 201368 152306 201420 152312
rect 200816 151276 200868 151282
rect 200816 151218 200868 151224
rect 201196 144006 201224 152306
rect 201184 144000 201236 144006
rect 201184 143942 201236 143948
rect 201380 143802 201408 152306
rect 201472 143870 201500 153854
rect 201656 152370 201684 153868
rect 201644 152364 201696 152370
rect 201644 152306 201696 152312
rect 201552 151276 201604 151282
rect 201552 151218 201604 151224
rect 201564 144074 201592 151218
rect 202116 151010 202144 153868
rect 202484 151418 202512 153868
rect 202472 151412 202524 151418
rect 202472 151354 202524 151360
rect 202104 151004 202156 151010
rect 202104 150946 202156 150952
rect 202748 151004 202800 151010
rect 202748 150946 202800 150952
rect 201552 144068 201604 144074
rect 201552 144010 201604 144016
rect 202196 144068 202248 144074
rect 202196 144010 202248 144016
rect 201736 144000 201788 144006
rect 201736 143942 201788 143948
rect 201460 143864 201512 143870
rect 201460 143806 201512 143812
rect 201368 143796 201420 143802
rect 201368 143738 201420 143744
rect 200264 142844 200316 142850
rect 200264 142786 200316 142792
rect 200908 142844 200960 142850
rect 200908 142786 200960 142792
rect 200184 142702 200396 142730
rect 200368 140826 200396 142702
rect 200920 140826 200948 142786
rect 201748 140826 201776 143942
rect 202208 140826 202236 144010
rect 202760 144006 202788 150946
rect 202748 144000 202800 144006
rect 202748 143942 202800 143948
rect 202852 143938 202880 153868
rect 203312 152302 203340 153868
rect 203680 152370 203708 153868
rect 203668 152364 203720 152370
rect 203668 152306 203720 152312
rect 203300 152296 203352 152302
rect 203300 152238 203352 152244
rect 204048 151486 204076 153868
rect 204508 152166 204536 153868
rect 204876 152234 204904 153868
rect 204864 152228 204916 152234
rect 204864 152170 204916 152176
rect 204496 152160 204548 152166
rect 204496 152102 204548 152108
rect 205244 151962 205272 153868
rect 205704 152098 205732 153868
rect 206086 153854 206376 153882
rect 205968 152364 206020 152370
rect 205968 152306 206020 152312
rect 205876 152296 205928 152302
rect 205876 152238 205928 152244
rect 205692 152092 205744 152098
rect 205692 152034 205744 152040
rect 205232 151956 205284 151962
rect 205232 151898 205284 151904
rect 204036 151480 204088 151486
rect 204036 151422 204088 151428
rect 203024 151412 203076 151418
rect 203024 151354 203076 151360
rect 203036 144074 203064 151354
rect 203024 144068 203076 144074
rect 203024 144010 203076 144016
rect 204496 144068 204548 144074
rect 204496 144010 204548 144016
rect 203852 144000 203904 144006
rect 203852 143942 203904 143948
rect 202840 143932 202892 143938
rect 202840 143874 202892 143880
rect 202748 143864 202800 143870
rect 202748 143806 202800 143812
rect 202760 140826 202788 143806
rect 203300 143796 203352 143802
rect 203300 143738 203352 143744
rect 203312 140826 203340 143738
rect 203864 140826 203892 143942
rect 204508 140826 204536 144010
rect 204956 143932 205008 143938
rect 204956 143874 205008 143880
rect 204968 140826 204996 143874
rect 205888 140962 205916 152238
rect 205980 141098 206008 152306
rect 206060 151480 206112 151486
rect 206060 151422 206112 151428
rect 206072 141234 206100 151422
rect 206348 151010 206376 153854
rect 206440 151486 206468 153868
rect 206428 151480 206480 151486
rect 206428 151422 206480 151428
rect 206900 151418 206928 153868
rect 207268 152302 207296 153868
rect 207256 152296 207308 152302
rect 207256 152238 207308 152244
rect 207348 152228 207400 152234
rect 207348 152170 207400 152176
rect 207256 152160 207308 152166
rect 207256 152102 207308 152108
rect 206888 151412 206940 151418
rect 206888 151354 206940 151360
rect 206336 151004 206388 151010
rect 206336 150946 206388 150952
rect 206072 141206 206744 141234
rect 205980 141070 206100 141098
rect 205888 140934 206008 140962
rect 199264 140798 199646 140826
rect 199724 140798 200198 140826
rect 200368 140798 200750 140826
rect 200920 140798 201302 140826
rect 201748 140798 201854 140826
rect 202208 140798 202498 140826
rect 202760 140798 203050 140826
rect 203312 140798 203602 140826
rect 203864 140798 204154 140826
rect 204508 140798 204706 140826
rect 204968 140798 205350 140826
rect 205980 140690 206008 140934
rect 206072 140826 206100 141070
rect 206716 140826 206744 141206
rect 207268 140826 207296 152102
rect 207360 140962 207388 152170
rect 207636 151350 207664 153868
rect 207992 152092 208044 152098
rect 207992 152034 208044 152040
rect 207900 151956 207952 151962
rect 207900 151898 207952 151904
rect 207624 151344 207676 151350
rect 207624 151286 207676 151292
rect 207912 144006 207940 151898
rect 208004 144074 208032 152034
rect 208096 151214 208124 153868
rect 208084 151208 208136 151214
rect 208084 151150 208136 151156
rect 208464 151146 208492 153868
rect 208832 151282 208860 153868
rect 208820 151276 208872 151282
rect 208820 151218 208872 151224
rect 208452 151140 208504 151146
rect 208452 151082 208504 151088
rect 209292 151078 209320 153868
rect 209280 151072 209332 151078
rect 209280 151014 209332 151020
rect 209660 151010 209688 153868
rect 212052 153730 212080 183751
rect 212144 179910 212172 190415
rect 212132 179904 212184 179910
rect 212132 179846 212184 179852
rect 216180 175892 216232 175898
rect 216180 175834 216232 175840
rect 212682 157160 212738 157169
rect 212682 157095 212684 157104
rect 212736 157095 212738 157104
rect 212684 157066 212736 157072
rect 212040 153724 212092 153730
rect 212040 153666 212092 153672
rect 210752 152296 210804 152302
rect 210752 152238 210804 152244
rect 210016 151480 210068 151486
rect 210016 151422 210068 151428
rect 208820 151004 208872 151010
rect 208820 150946 208872 150952
rect 209648 151004 209700 151010
rect 209648 150946 209700 150952
rect 207992 144068 208044 144074
rect 207992 144010 208044 144016
rect 208728 144068 208780 144074
rect 208728 144010 208780 144016
rect 207900 144000 207952 144006
rect 207900 143942 207952 143948
rect 208636 144000 208688 144006
rect 208636 143942 208688 143948
rect 207360 140934 207756 140962
rect 206072 140798 206454 140826
rect 206716 140798 207006 140826
rect 207268 140798 207558 140826
rect 189342 140662 189448 140690
rect 192746 140662 193036 140690
rect 193298 140662 193404 140690
rect 193942 140662 194232 140690
rect 194494 140662 194784 140690
rect 195046 140662 195152 140690
rect 196150 140662 196256 140690
rect 199002 140662 199108 140690
rect 205902 140662 206008 140690
rect 207728 140690 207756 140934
rect 208648 140826 208676 143942
rect 208740 141098 208768 144010
rect 208832 141234 208860 150946
rect 208832 141206 209412 141234
rect 208740 141070 208952 141098
rect 208924 140826 208952 141070
rect 208648 140798 208754 140826
rect 208924 140798 209306 140826
rect 209384 140690 209412 141206
rect 210028 140826 210056 151422
rect 210108 151412 210160 151418
rect 210108 151354 210160 151360
rect 210120 140962 210148 151354
rect 210660 151344 210712 151350
rect 210660 151286 210712 151292
rect 210672 143938 210700 151286
rect 210764 144074 210792 152238
rect 212868 151276 212920 151282
rect 212868 151218 212920 151224
rect 210844 151208 210896 151214
rect 210844 151150 210896 151156
rect 210752 144068 210804 144074
rect 210752 144010 210804 144016
rect 210856 144006 210884 151150
rect 210936 151140 210988 151146
rect 210936 151082 210988 151088
rect 210844 144000 210896 144006
rect 210844 143942 210896 143948
rect 210660 143932 210712 143938
rect 210660 143874 210712 143880
rect 210948 143870 210976 151082
rect 212880 146266 212908 151218
rect 214156 151072 214208 151078
rect 214156 151014 214208 151020
rect 212880 146238 213184 146266
rect 211396 144068 211448 144074
rect 211396 144010 211448 144016
rect 210936 143864 210988 143870
rect 210936 143806 210988 143812
rect 210120 140934 210516 140962
rect 210028 140798 210410 140826
rect 210488 140690 210516 140934
rect 211408 140826 211436 144010
rect 212316 144000 212368 144006
rect 212316 143942 212368 143948
rect 211764 143932 211816 143938
rect 211764 143874 211816 143880
rect 211776 140826 211804 143874
rect 212328 140826 212356 143942
rect 212960 143864 213012 143870
rect 212960 143806 213012 143812
rect 212972 140826 213000 143806
rect 213156 141370 213184 146238
rect 213156 141342 213552 141370
rect 213524 140826 213552 141342
rect 214168 140826 214196 151014
rect 214248 151004 214300 151010
rect 214248 150946 214300 150952
rect 214260 140962 214288 150946
rect 215628 143388 215680 143394
rect 215628 143330 215680 143336
rect 214260 140934 214564 140962
rect 211408 140798 211606 140826
rect 211776 140798 212158 140826
rect 212328 140798 212710 140826
rect 212972 140798 213262 140826
rect 213524 140798 213906 140826
rect 214168 140798 214458 140826
rect 214536 140690 214564 140934
rect 215640 140690 215668 143330
rect 207728 140662 208202 140690
rect 209384 140662 209858 140690
rect 210488 140662 211054 140690
rect 214536 140662 215010 140690
rect 215562 140662 215668 140690
rect 184990 140160 185046 140169
rect 184990 140095 185046 140104
rect 167400 138758 167736 138786
rect 177632 138560 177684 138566
rect 177632 138502 177684 138508
rect 177722 138528 177778 138537
rect 177644 138265 177672 138502
rect 185004 138498 185032 140095
rect 185082 140024 185138 140033
rect 185082 139959 185138 139968
rect 185096 138566 185124 139959
rect 185358 138936 185414 138945
rect 185358 138871 185414 138880
rect 185266 138664 185322 138673
rect 185266 138599 185322 138608
rect 185084 138560 185136 138566
rect 185084 138502 185136 138508
rect 177722 138463 177724 138472
rect 177776 138463 177778 138472
rect 184992 138492 185044 138498
rect 177724 138434 177776 138440
rect 184992 138434 185044 138440
rect 177630 138256 177686 138265
rect 177630 138191 177686 138200
rect 185174 137848 185230 137857
rect 185174 137783 185230 137792
rect 185188 137274 185216 137783
rect 181588 137268 181640 137274
rect 181588 137210 181640 137216
rect 185176 137268 185228 137274
rect 185176 137210 185228 137216
rect 177724 137132 177776 137138
rect 177724 137074 177776 137080
rect 177632 137064 177684 137070
rect 177736 137041 177764 137074
rect 177632 137006 177684 137012
rect 177722 137032 177778 137041
rect 177644 136905 177672 137006
rect 177722 136967 177778 136976
rect 177630 136896 177686 136905
rect 177630 136831 177686 136840
rect 181600 136662 181628 137210
rect 182232 137200 182284 137206
rect 182232 137142 182284 137148
rect 177724 136656 177776 136662
rect 177724 136598 177776 136604
rect 181588 136656 181640 136662
rect 181588 136598 181640 136604
rect 177736 136361 177764 136598
rect 177722 136352 177778 136361
rect 177722 136287 177778 136296
rect 181956 135840 182008 135846
rect 181956 135782 182008 135788
rect 177632 135772 177684 135778
rect 177632 135714 177684 135720
rect 177644 135273 177672 135714
rect 177724 135704 177776 135710
rect 177724 135646 177776 135652
rect 177736 135545 177764 135646
rect 177722 135536 177778 135545
rect 177722 135471 177778 135480
rect 177630 135264 177686 135273
rect 177630 135199 177686 135208
rect 177632 134412 177684 134418
rect 177632 134354 177684 134360
rect 177644 133505 177672 134354
rect 181968 134350 181996 135782
rect 182244 135710 182272 137142
rect 185280 137070 185308 138599
rect 185372 137138 185400 138871
rect 185450 137304 185506 137313
rect 185450 137239 185506 137248
rect 185464 137206 185492 137239
rect 185452 137200 185504 137206
rect 185452 137142 185504 137148
rect 185360 137132 185412 137138
rect 185360 137074 185412 137080
rect 185268 137064 185320 137070
rect 185268 137006 185320 137012
rect 185174 136624 185230 136633
rect 185174 136559 185230 136568
rect 182324 135908 182376 135914
rect 182324 135850 182376 135856
rect 182232 135704 182284 135710
rect 182232 135646 182284 135652
rect 177724 134344 177776 134350
rect 177722 134312 177724 134321
rect 181956 134344 182008 134350
rect 177776 134312 177778 134321
rect 181956 134286 182008 134292
rect 177722 134247 177778 134256
rect 182336 134078 182364 135850
rect 185188 135778 185216 136559
rect 185266 136080 185322 136089
rect 185266 136015 185322 136024
rect 185280 135846 185308 136015
rect 185358 135944 185414 135953
rect 185358 135879 185360 135888
rect 185412 135879 185414 135888
rect 185360 135850 185412 135856
rect 185268 135840 185320 135846
rect 185268 135782 185320 135788
rect 185176 135772 185228 135778
rect 185176 135714 185228 135720
rect 185174 134856 185230 134865
rect 185174 134791 185230 134800
rect 185082 134448 185138 134457
rect 185188 134418 185216 134791
rect 185082 134383 185138 134392
rect 185176 134412 185228 134418
rect 177724 134072 177776 134078
rect 177724 134014 177776 134020
rect 182324 134072 182376 134078
rect 182324 134014 182376 134020
rect 177736 133913 177764 134014
rect 177722 133904 177778 133913
rect 177722 133839 177778 133848
rect 177630 133496 177686 133505
rect 177630 133431 177686 133440
rect 177632 132984 177684 132990
rect 177632 132926 177684 132932
rect 177644 132281 177672 132926
rect 185096 132922 185124 134383
rect 185176 134354 185228 134360
rect 185174 133768 185230 133777
rect 185174 133703 185230 133712
rect 185188 132990 185216 133703
rect 185818 133088 185874 133097
rect 185818 133023 185874 133032
rect 185176 132984 185228 132990
rect 185176 132926 185228 132932
rect 177724 132916 177776 132922
rect 177724 132858 177776 132864
rect 185084 132916 185136 132922
rect 185084 132858 185136 132864
rect 177736 132689 177764 132858
rect 177722 132680 177778 132689
rect 177722 132615 177778 132624
rect 185450 132544 185506 132553
rect 185450 132479 185506 132488
rect 177630 132272 177686 132281
rect 177630 132207 177686 132216
rect 185464 131630 185492 132479
rect 185726 132000 185782 132009
rect 185726 131935 185782 131944
rect 185542 131728 185598 131737
rect 185542 131663 185598 131672
rect 177632 131624 177684 131630
rect 177632 131566 177684 131572
rect 185452 131624 185504 131630
rect 185452 131566 185504 131572
rect 177644 131057 177672 131566
rect 177724 131556 177776 131562
rect 177724 131498 177776 131504
rect 177736 131329 177764 131498
rect 177722 131320 177778 131329
rect 177722 131255 177778 131264
rect 177630 131048 177686 131057
rect 177630 130983 177686 130992
rect 185266 130776 185322 130785
rect 185266 130711 185322 130720
rect 177632 130264 177684 130270
rect 177632 130206 177684 130212
rect 177722 130232 177778 130241
rect 177644 129833 177672 130206
rect 177722 130167 177724 130176
rect 177776 130167 177778 130176
rect 177724 130138 177776 130144
rect 177630 129824 177686 129833
rect 177630 129759 177686 129768
rect 185174 129688 185230 129697
rect 185174 129623 185230 129632
rect 177724 128904 177776 128910
rect 177724 128846 177776 128852
rect 177632 128768 177684 128774
rect 177736 128745 177764 128846
rect 185188 128842 185216 129623
rect 185280 128910 185308 130711
rect 185358 130368 185414 130377
rect 185358 130303 185414 130312
rect 185268 128904 185320 128910
rect 185268 128846 185320 128852
rect 177816 128836 177868 128842
rect 177816 128778 177868 128784
rect 185176 128836 185228 128842
rect 185176 128778 185228 128784
rect 177632 128710 177684 128716
rect 177722 128736 177778 128745
rect 177644 128473 177672 128710
rect 177722 128671 177778 128680
rect 177630 128464 177686 128473
rect 177630 128399 177686 128408
rect 177828 128065 177856 128778
rect 185372 128774 185400 130303
rect 185556 130270 185584 131663
rect 185544 130264 185596 130270
rect 185544 130206 185596 130212
rect 185740 130202 185768 131935
rect 185832 131562 185860 133023
rect 185820 131556 185872 131562
rect 185820 131498 185872 131504
rect 185728 130196 185780 130202
rect 185728 130138 185780 130144
rect 185450 129008 185506 129017
rect 185450 128943 185506 128952
rect 185360 128768 185412 128774
rect 185360 128710 185412 128716
rect 185174 128464 185230 128473
rect 185174 128399 185230 128408
rect 177814 128056 177870 128065
rect 177814 127991 177870 128000
rect 185188 127482 185216 128399
rect 185358 127920 185414 127929
rect 185358 127855 185414 127864
rect 185266 127648 185322 127657
rect 185266 127583 185322 127592
rect 177724 127476 177776 127482
rect 177724 127418 177776 127424
rect 185176 127476 185228 127482
rect 185176 127418 185228 127424
rect 177172 127408 177224 127414
rect 177172 127350 177224 127356
rect 177184 127249 177212 127350
rect 177170 127240 177226 127249
rect 177170 127175 177226 127184
rect 177736 126977 177764 127418
rect 177722 126968 177778 126977
rect 177722 126903 177778 126912
rect 185174 126288 185230 126297
rect 182232 126252 182284 126258
rect 185174 126223 185230 126232
rect 182232 126194 182284 126200
rect 177724 126116 177776 126122
rect 177724 126058 177776 126064
rect 177632 126048 177684 126054
rect 177736 126025 177764 126058
rect 177632 125990 177684 125996
rect 177722 126016 177778 126025
rect 177644 125617 177672 125990
rect 177722 125951 177778 125960
rect 177630 125608 177686 125617
rect 177630 125543 177686 125552
rect 177632 124756 177684 124762
rect 177632 124698 177684 124704
rect 177172 124416 177224 124422
rect 177172 124358 177224 124364
rect 177184 124257 177212 124358
rect 177170 124248 177226 124257
rect 177170 124183 177226 124192
rect 177644 123985 177672 124698
rect 182244 124694 182272 126194
rect 185188 126190 185216 126223
rect 182324 126184 182376 126190
rect 182324 126126 182376 126132
rect 185176 126184 185228 126190
rect 185176 126126 185228 126132
rect 177724 124688 177776 124694
rect 177724 124630 177776 124636
rect 182232 124688 182284 124694
rect 182232 124630 182284 124636
rect 177736 124529 177764 124630
rect 177722 124520 177778 124529
rect 177722 124455 177778 124464
rect 182336 124422 182364 126126
rect 185280 126054 185308 127583
rect 185372 126122 185400 127855
rect 185464 127414 185492 128943
rect 216192 127482 216220 175834
rect 216928 157130 216956 211495
rect 220332 205449 220360 220743
rect 220318 205440 220374 205449
rect 220318 205375 220374 205384
rect 222344 179904 222396 179910
rect 222344 179846 222396 179852
rect 222356 179201 222384 179846
rect 222342 179192 222398 179201
rect 222342 179127 222398 179136
rect 217008 163652 217060 163658
rect 217008 163594 217060 163600
rect 216916 157124 216968 157130
rect 216916 157066 216968 157072
rect 216928 156518 216956 157066
rect 216916 156512 216968 156518
rect 216916 156454 216968 156460
rect 216180 127476 216232 127482
rect 216180 127418 216232 127424
rect 185452 127408 185504 127414
rect 217020 127385 217048 163594
rect 218296 156512 218348 156518
rect 218296 156454 218348 156460
rect 185452 127350 185504 127356
rect 217006 127376 217062 127385
rect 217006 127311 217062 127320
rect 185450 126696 185506 126705
rect 185450 126631 185506 126640
rect 185464 126258 185492 126631
rect 185452 126252 185504 126258
rect 185452 126194 185504 126200
rect 185360 126116 185412 126122
rect 185360 126058 185412 126064
rect 185268 126048 185320 126054
rect 185268 125990 185320 125996
rect 185174 125608 185230 125617
rect 185174 125543 185230 125552
rect 185188 124762 185216 125543
rect 185450 124928 185506 124937
rect 185450 124863 185506 124872
rect 185358 124792 185414 124801
rect 185176 124756 185228 124762
rect 185358 124727 185414 124736
rect 185176 124698 185228 124704
rect 182324 124416 182376 124422
rect 182324 124358 182376 124364
rect 177630 123976 177686 123985
rect 177630 123911 177686 123920
rect 185266 123432 185322 123441
rect 185266 123367 185322 123376
rect 177632 123328 177684 123334
rect 177632 123270 177684 123276
rect 177644 122761 177672 123270
rect 177724 123260 177776 123266
rect 177724 123202 177776 123208
rect 177736 123033 177764 123202
rect 177722 123024 177778 123033
rect 177722 122959 177778 122968
rect 177630 122752 177686 122761
rect 177630 122687 177686 122696
rect 177724 121968 177776 121974
rect 177724 121910 177776 121916
rect 177356 121900 177408 121906
rect 177356 121842 177408 121848
rect 177368 121537 177396 121842
rect 177736 121809 177764 121910
rect 185280 121906 185308 123367
rect 185372 123334 185400 124727
rect 185360 123328 185412 123334
rect 185360 123270 185412 123276
rect 185464 123266 185492 124863
rect 185818 123840 185874 123849
rect 185818 123775 185874 123784
rect 185452 123260 185504 123266
rect 185452 123202 185504 123208
rect 185634 122616 185690 122625
rect 185634 122551 185690 122560
rect 185268 121900 185320 121906
rect 185268 121842 185320 121848
rect 177722 121800 177778 121809
rect 177722 121735 177778 121744
rect 177354 121528 177410 121537
rect 177354 121463 177410 121472
rect 185358 121528 185414 121537
rect 185358 121463 185414 121472
rect 185174 120848 185230 120857
rect 182048 120812 182100 120818
rect 185372 120818 185400 121463
rect 185174 120783 185230 120792
rect 185360 120812 185412 120818
rect 182048 120754 182100 120760
rect 181588 120676 181640 120682
rect 181588 120618 181640 120624
rect 177632 120608 177684 120614
rect 177632 120550 177684 120556
rect 177722 120576 177778 120585
rect 177644 120313 177672 120550
rect 177722 120511 177724 120520
rect 177776 120511 177778 120520
rect 177724 120482 177776 120488
rect 177630 120304 177686 120313
rect 177630 120239 177686 120248
rect 177724 119112 177776 119118
rect 177722 119080 177724 119089
rect 177776 119080 177778 119089
rect 177722 119015 177778 119024
rect 181600 118982 181628 120618
rect 182060 119118 182088 120754
rect 182324 120744 182376 120750
rect 182324 120686 182376 120692
rect 182140 119384 182192 119390
rect 182140 119326 182192 119332
rect 182048 119112 182100 119118
rect 182048 119054 182100 119060
rect 177724 118976 177776 118982
rect 177724 118918 177776 118924
rect 181588 118976 181640 118982
rect 181588 118918 181640 118924
rect 177632 118840 177684 118846
rect 177736 118817 177764 118918
rect 177632 118782 177684 118788
rect 177722 118808 177778 118817
rect 177644 118545 177672 118782
rect 177722 118743 177778 118752
rect 177630 118536 177686 118545
rect 177630 118471 177686 118480
rect 182048 117956 182100 117962
rect 182048 117898 182100 117904
rect 177724 117752 177776 117758
rect 177724 117694 177776 117700
rect 177736 117593 177764 117694
rect 177722 117584 177778 117593
rect 177722 117519 177778 117528
rect 177172 117480 177224 117486
rect 177172 117422 177224 117428
rect 177184 117185 177212 117422
rect 177170 117176 177226 117185
rect 177170 117111 177226 117120
rect 178184 116596 178236 116602
rect 178184 116538 178236 116544
rect 176804 116528 176856 116534
rect 176804 116470 176856 116476
rect 175424 115236 175476 115242
rect 175424 115178 175476 115184
rect 174780 115168 174832 115174
rect 174780 115110 174832 115116
rect 145352 114822 145596 114850
rect 146976 114822 147312 114850
rect 145352 110958 145380 114822
rect 147284 113338 147312 114822
rect 148112 114822 148448 114850
rect 149308 114822 149828 114850
rect 150688 114822 151300 114850
rect 152068 114822 152680 114850
rect 153448 114822 154152 114850
rect 154828 114822 155532 114850
rect 156208 114822 157004 114850
rect 158048 114822 158384 114850
rect 159520 114822 159856 114850
rect 160900 114822 161236 114850
rect 161728 114822 162708 114850
rect 163752 114822 164088 114850
rect 164488 114822 165560 114850
rect 166604 114822 166940 114850
rect 168076 114822 168412 114850
rect 169456 114822 169792 114850
rect 170928 114822 171264 114850
rect 172644 114822 172704 114850
rect 147272 113332 147324 113338
rect 147272 113274 147324 113280
rect 148112 111638 148140 114822
rect 148100 111632 148152 111638
rect 148100 111574 148152 111580
rect 145340 110952 145392 110958
rect 145340 110894 145392 110900
rect 143776 102384 143828 102390
rect 143776 102326 143828 102332
rect 143684 102316 143736 102322
rect 143684 102258 143736 102264
rect 142672 101976 142724 101982
rect 142672 101918 142724 101924
rect 142684 99740 142712 101918
rect 143788 99740 143816 102326
rect 144880 102248 144932 102254
rect 144880 102190 144932 102196
rect 144892 99740 144920 102190
rect 145984 102180 146036 102186
rect 145984 102122 146036 102128
rect 145996 99740 146024 102122
rect 147088 102112 147140 102118
rect 147088 102054 147140 102060
rect 147100 99740 147128 102054
rect 148192 102044 148244 102050
rect 148192 101986 148244 101992
rect 148204 99740 148232 101986
rect 149308 99740 149336 114822
rect 150688 101386 150716 114822
rect 152068 101386 152096 114822
rect 150504 101358 150716 101386
rect 151976 101358 152096 101386
rect 153448 101370 153476 114822
rect 154828 101370 154856 114822
rect 156208 101438 156236 114822
rect 158048 111026 158076 114822
rect 158864 111088 158916 111094
rect 158864 111030 158916 111036
rect 156840 111020 156892 111026
rect 156840 110962 156892 110968
rect 158036 111020 158088 111026
rect 158036 110962 158088 110968
rect 158312 111020 158364 111026
rect 158312 110962 158364 110968
rect 154908 101432 154960 101438
rect 154908 101374 154960 101380
rect 156196 101432 156248 101438
rect 156196 101374 156248 101380
rect 152608 101364 152660 101370
rect 150504 99754 150532 101358
rect 151976 99754 152004 101358
rect 152608 101306 152660 101312
rect 153436 101364 153488 101370
rect 153436 101306 153488 101312
rect 153804 101364 153856 101370
rect 153804 101306 153856 101312
rect 154816 101364 154868 101370
rect 154816 101306 154868 101312
rect 150426 99726 150532 99754
rect 151530 99726 152004 99754
rect 152620 99740 152648 101306
rect 153816 99740 153844 101306
rect 154920 99740 154948 101374
rect 156852 101370 156880 110962
rect 158220 101432 158272 101438
rect 158220 101374 158272 101380
rect 156012 101364 156064 101370
rect 156012 101306 156064 101312
rect 156840 101364 156892 101370
rect 156840 101306 156892 101312
rect 157116 101364 157168 101370
rect 157116 101306 157168 101312
rect 156024 99740 156052 101306
rect 157128 99740 157156 101306
rect 158232 99740 158260 101374
rect 158324 101370 158352 110962
rect 158876 101438 158904 111030
rect 159520 111026 159548 114822
rect 160900 111094 160928 114822
rect 160888 111088 160940 111094
rect 160888 111030 160940 111036
rect 159508 111020 159560 111026
rect 159508 110962 159560 110968
rect 161624 111020 161676 111026
rect 161624 110962 161676 110968
rect 161532 102044 161584 102050
rect 161532 101986 161584 101992
rect 159324 101636 159376 101642
rect 159324 101578 159376 101584
rect 158864 101432 158916 101438
rect 158864 101374 158916 101380
rect 158312 101364 158364 101370
rect 158312 101306 158364 101312
rect 159336 99740 159364 101578
rect 160428 101364 160480 101370
rect 160428 101306 160480 101312
rect 160440 99740 160468 101306
rect 161544 99740 161572 101986
rect 161636 101370 161664 110962
rect 161728 101642 161756 114822
rect 163752 111026 163780 114822
rect 163832 111156 163884 111162
rect 163832 111098 163884 111104
rect 163740 111020 163792 111026
rect 163740 110962 163792 110968
rect 161716 101636 161768 101642
rect 161716 101578 161768 101584
rect 163740 101432 163792 101438
rect 163740 101374 163792 101380
rect 161624 101364 161676 101370
rect 161624 101306 161676 101312
rect 162636 101364 162688 101370
rect 162636 101306 162688 101312
rect 162648 99740 162676 101306
rect 163752 99740 163780 101374
rect 163844 101370 163872 111098
rect 164488 102050 164516 114822
rect 166604 111162 166632 114822
rect 166592 111156 166644 111162
rect 166592 111098 166644 111104
rect 167880 111156 167932 111162
rect 167880 111098 167932 111104
rect 166500 111088 166552 111094
rect 166500 111030 166552 111036
rect 165120 111020 165172 111026
rect 165120 110962 165172 110968
rect 164476 102044 164528 102050
rect 164476 101986 164528 101992
rect 165132 101438 165160 110962
rect 165120 101432 165172 101438
rect 165120 101374 165172 101380
rect 165948 101432 166000 101438
rect 165948 101374 166000 101380
rect 163832 101364 163884 101370
rect 163832 101306 163884 101312
rect 164844 101364 164896 101370
rect 164844 101306 164896 101312
rect 164856 99740 164884 101306
rect 165960 99740 165988 101374
rect 166512 101370 166540 111030
rect 167144 102316 167196 102322
rect 167144 102258 167196 102264
rect 166500 101364 166552 101370
rect 166500 101306 166552 101312
rect 167156 99740 167184 102258
rect 167892 101438 167920 111098
rect 168076 111026 168104 114822
rect 169456 111094 169484 114822
rect 169904 112380 169956 112386
rect 169904 112322 169956 112328
rect 169444 111088 169496 111094
rect 169444 111030 169496 111036
rect 168064 111020 168116 111026
rect 168064 110962 168116 110968
rect 167880 101432 167932 101438
rect 167880 101374 167932 101380
rect 169916 99890 169944 112322
rect 170928 111162 170956 114822
rect 170916 111156 170968 111162
rect 170916 111098 170968 111104
rect 172676 111026 172704 114822
rect 172664 111020 172716 111026
rect 172664 110962 172716 110968
rect 172664 102112 172716 102118
rect 172664 102054 172716 102060
rect 171560 102044 171612 102050
rect 171560 101986 171612 101992
rect 170456 101976 170508 101982
rect 170456 101918 170508 101924
rect 169824 99862 169944 99890
rect 169824 99754 169852 99862
rect 169378 99726 169852 99754
rect 170468 99740 170496 101918
rect 171572 99740 171600 101986
rect 172676 99740 172704 102054
rect 174792 101370 174820 115110
rect 173768 101364 173820 101370
rect 173768 101306 173820 101312
rect 174780 101364 174832 101370
rect 174780 101306 174832 101312
rect 173780 99740 173808 101306
rect 175436 99618 175464 115178
rect 176160 111020 176212 111026
rect 176160 110962 176212 110968
rect 176172 101438 176200 110962
rect 176160 101432 176212 101438
rect 176160 101374 176212 101380
rect 176816 101370 176844 116470
rect 177080 116460 177132 116466
rect 177080 116402 177132 116408
rect 177092 115553 177120 116402
rect 177724 116392 177776 116398
rect 177722 116360 177724 116369
rect 177776 116360 177778 116369
rect 177722 116295 177778 116304
rect 177724 116120 177776 116126
rect 177724 116062 177776 116068
rect 177736 115961 177764 116062
rect 177722 115952 177778 115961
rect 177722 115887 177778 115896
rect 177078 115544 177134 115553
rect 177078 115479 177134 115488
rect 178196 101370 178224 116538
rect 182060 116398 182088 117898
rect 182152 117758 182180 119326
rect 182232 119316 182284 119322
rect 182232 119258 182284 119264
rect 182140 117752 182192 117758
rect 182140 117694 182192 117700
rect 182244 117486 182272 119258
rect 182336 118846 182364 120686
rect 185188 120682 185216 120783
rect 185360 120754 185412 120760
rect 185268 120744 185320 120750
rect 185266 120712 185268 120721
rect 185320 120712 185322 120721
rect 185176 120676 185228 120682
rect 185266 120647 185322 120656
rect 185176 120618 185228 120624
rect 185648 120546 185676 122551
rect 185832 121974 185860 123775
rect 185910 122208 185966 122217
rect 185910 122143 185966 122152
rect 185820 121968 185872 121974
rect 185820 121910 185872 121916
rect 185924 120614 185952 122143
rect 185912 120608 185964 120614
rect 185912 120550 185964 120556
rect 185636 120540 185688 120546
rect 185636 120482 185688 120488
rect 185266 119760 185322 119769
rect 185266 119695 185322 119704
rect 185280 119390 185308 119695
rect 185268 119384 185320 119390
rect 185174 119352 185230 119361
rect 185268 119326 185320 119332
rect 185174 119287 185176 119296
rect 185228 119287 185230 119296
rect 185176 119258 185228 119264
rect 182324 118840 182376 118846
rect 182324 118782 182376 118788
rect 185266 118536 185322 118545
rect 185266 118471 185322 118480
rect 185174 117992 185230 118001
rect 185280 117962 185308 118471
rect 185174 117927 185230 117936
rect 185268 117956 185320 117962
rect 185188 117894 185216 117927
rect 185268 117898 185320 117904
rect 182324 117888 182376 117894
rect 182324 117830 182376 117836
rect 185176 117888 185228 117894
rect 218308 117865 218336 156454
rect 222252 153724 222304 153730
rect 222252 153666 222304 153672
rect 222264 152953 222292 153666
rect 222250 152944 222306 152953
rect 222250 152879 222306 152888
rect 218386 135944 218442 135953
rect 218386 135879 218442 135888
rect 185176 117830 185228 117836
rect 218294 117856 218350 117865
rect 182232 117480 182284 117486
rect 182232 117422 182284 117428
rect 182048 116392 182100 116398
rect 182048 116334 182100 116340
rect 182336 116126 182364 117830
rect 218294 117791 218350 117800
rect 185358 117448 185414 117457
rect 185358 117383 185414 117392
rect 185266 116768 185322 116777
rect 185266 116703 185322 116712
rect 185280 116602 185308 116703
rect 185268 116596 185320 116602
rect 185268 116538 185320 116544
rect 185176 116528 185228 116534
rect 185174 116496 185176 116505
rect 185228 116496 185230 116505
rect 185372 116466 185400 117383
rect 185174 116431 185230 116440
rect 185360 116460 185412 116466
rect 185360 116402 185412 116408
rect 182324 116120 182376 116126
rect 182324 116062 182376 116068
rect 185266 115680 185322 115689
rect 185266 115615 185322 115624
rect 185174 115272 185230 115281
rect 185280 115242 185308 115615
rect 185174 115207 185230 115216
rect 185268 115236 185320 115242
rect 185188 115174 185216 115207
rect 185268 115178 185320 115184
rect 185176 115168 185228 115174
rect 185176 115110 185228 115116
rect 186002 114456 186058 114465
rect 186002 114391 186058 114400
rect 185818 113912 185874 113921
rect 185818 113847 185874 113856
rect 185174 112688 185230 112697
rect 185174 112623 185230 112632
rect 185188 112386 185216 112623
rect 185176 112380 185228 112386
rect 185176 112322 185228 112328
rect 183612 110408 183664 110414
rect 183612 110350 183664 110356
rect 183520 110272 183572 110278
rect 183520 110214 183572 110220
rect 183336 109864 183388 109870
rect 183336 109806 183388 109812
rect 183244 109796 183296 109802
rect 183244 109738 183296 109744
rect 183152 109728 183204 109734
rect 183152 109670 183204 109676
rect 183060 109660 183112 109666
rect 183060 109602 183112 109608
rect 179288 101432 179340 101438
rect 179288 101374 179340 101380
rect 175976 101364 176028 101370
rect 175976 101306 176028 101312
rect 176804 101364 176856 101370
rect 176804 101306 176856 101312
rect 177080 101364 177132 101370
rect 177080 101306 177132 101312
rect 178184 101364 178236 101370
rect 178184 101306 178236 101312
rect 175988 99740 176016 101306
rect 177092 99740 177120 101306
rect 179300 99740 179328 101374
rect 174898 99590 175464 99618
rect 183072 90665 183100 109602
rect 183164 91889 183192 109670
rect 183256 94337 183284 109738
rect 183348 95561 183376 109806
rect 183428 109592 183480 109598
rect 183428 109534 183480 109540
rect 183334 95552 183390 95561
rect 183334 95487 183390 95496
rect 183242 94328 183298 94337
rect 183242 94263 183298 94272
rect 183440 93113 183468 109534
rect 183532 96785 183560 110214
rect 183624 98009 183652 110350
rect 183704 110340 183756 110346
rect 183704 110282 183756 110288
rect 183716 99233 183744 110282
rect 185832 102050 185860 113847
rect 186016 102118 186044 114391
rect 186186 113776 186242 113785
rect 186186 113711 186242 113720
rect 186004 102112 186056 102118
rect 186004 102054 186056 102060
rect 185820 102044 185872 102050
rect 185820 101986 185872 101992
rect 186200 101982 186228 113711
rect 218400 113338 218428 135879
rect 222344 127476 222396 127482
rect 222344 127418 222396 127424
rect 222356 126841 222384 127418
rect 222342 126832 222398 126841
rect 222342 126767 222398 126776
rect 218388 113332 218440 113338
rect 218388 113274 218440 113280
rect 199816 113054 200198 113082
rect 207636 113054 208202 113082
rect 188224 109666 188252 112932
rect 188776 109734 188804 112932
rect 188764 109728 188816 109734
rect 188764 109670 188816 109676
rect 188212 109660 188264 109666
rect 188212 109602 188264 109608
rect 189328 109598 189356 112932
rect 189880 109802 189908 112932
rect 190432 109870 190460 112932
rect 191076 110278 191104 112932
rect 191628 110414 191656 112932
rect 191616 110408 191668 110414
rect 191616 110350 191668 110356
rect 192180 110346 192208 112932
rect 192746 112918 193036 112946
rect 193298 112918 193404 112946
rect 193008 112538 193036 112918
rect 193008 112510 193312 112538
rect 192168 110340 192220 110346
rect 192168 110282 192220 110288
rect 191064 110272 191116 110278
rect 191064 110214 191116 110220
rect 191984 110272 192036 110278
rect 191984 110214 192036 110220
rect 190420 109864 190472 109870
rect 190420 109806 190472 109812
rect 189868 109796 189920 109802
rect 189868 109738 189920 109744
rect 189316 109592 189368 109598
rect 189316 109534 189368 109540
rect 186188 101976 186240 101982
rect 186188 101918 186240 101924
rect 183702 99224 183758 99233
rect 183702 99159 183758 99168
rect 191996 98825 192024 110214
rect 193284 102662 193312 112510
rect 193272 102656 193324 102662
rect 193272 102598 193324 102604
rect 193376 101438 193404 112918
rect 193928 109598 193956 112932
rect 194494 112918 194692 112946
rect 193916 109592 193968 109598
rect 193916 109534 193968 109540
rect 194100 102656 194152 102662
rect 194100 102598 194152 102604
rect 193364 101432 193416 101438
rect 193364 101374 193416 101380
rect 194112 99740 194140 102598
rect 194468 101432 194520 101438
rect 194468 101374 194520 101380
rect 194480 99740 194508 101374
rect 194664 101370 194692 112918
rect 194744 109592 194796 109598
rect 194744 109534 194796 109540
rect 194652 101364 194704 101370
rect 194652 101306 194704 101312
rect 194756 99618 194784 109534
rect 194928 102724 194980 102730
rect 194928 102666 194980 102672
rect 194940 101370 194968 102666
rect 194928 101364 194980 101370
rect 194928 101306 194980 101312
rect 194928 101228 194980 101234
rect 194928 101170 194980 101176
rect 194940 99754 194968 101170
rect 195032 100842 195060 112932
rect 195124 112918 195598 112946
rect 195124 102730 195152 112918
rect 195112 102724 195164 102730
rect 195112 102666 195164 102672
rect 196136 101386 196164 112932
rect 196320 112918 196794 112946
rect 197056 112918 197346 112946
rect 197700 112918 197898 112946
rect 198160 112918 198450 112946
rect 199002 112918 199108 112946
rect 196320 102662 196348 112918
rect 196308 102656 196360 102662
rect 196308 102598 196360 102604
rect 196860 102656 196912 102662
rect 196860 102598 196912 102604
rect 196032 101364 196084 101370
rect 196136 101358 196256 101386
rect 196032 101306 196084 101312
rect 195032 100814 195428 100842
rect 195400 99754 195428 100814
rect 194940 99726 195322 99754
rect 195400 99726 195690 99754
rect 196044 99740 196072 101306
rect 196228 99754 196256 101358
rect 196228 99726 196518 99754
rect 196872 99740 196900 102598
rect 197056 99754 197084 112918
rect 197056 99726 197254 99754
rect 197700 99740 197728 112918
rect 198160 99754 198188 112918
rect 199080 102730 199108 112918
rect 199172 112918 199646 112946
rect 199068 102724 199120 102730
rect 199068 102666 199120 102672
rect 198424 102656 198476 102662
rect 199172 102610 199200 112918
rect 199816 112674 199844 113054
rect 199724 112646 199844 112674
rect 200368 112918 200750 112946
rect 201012 112918 201302 112946
rect 201748 112918 201854 112946
rect 198424 102598 198476 102604
rect 198082 99726 198188 99754
rect 198436 99740 198464 102598
rect 198896 102582 199200 102610
rect 199620 102656 199672 102662
rect 199620 102598 199672 102604
rect 199252 102588 199304 102594
rect 198896 99740 198924 102582
rect 199252 102530 199304 102536
rect 199264 99740 199292 102530
rect 199632 99740 199660 102598
rect 199724 102594 199752 112646
rect 200368 102662 200396 112918
rect 201012 112674 201040 112918
rect 200644 112646 201040 112674
rect 200356 102656 200408 102662
rect 200356 102598 200408 102604
rect 199712 102588 199764 102594
rect 199712 102530 199764 102536
rect 200644 102066 200672 112646
rect 201748 109682 201776 112918
rect 201460 109660 201512 109666
rect 201460 109602 201512 109608
rect 201564 109654 201776 109682
rect 200816 102656 200868 102662
rect 200816 102598 200868 102604
rect 200276 102038 200672 102066
rect 200276 99754 200304 102038
rect 200448 101908 200500 101914
rect 200448 101850 200500 101856
rect 200106 99726 200304 99754
rect 200460 99740 200488 101850
rect 200828 99740 200856 102598
rect 201472 99754 201500 109602
rect 201564 101914 201592 109654
rect 202484 109598 202512 112932
rect 203036 109666 203064 112932
rect 203128 112918 203602 112946
rect 203772 112918 204154 112946
rect 203024 109660 203076 109666
rect 203024 109602 203076 109608
rect 201644 109592 201696 109598
rect 201644 109534 201696 109540
rect 202472 109592 202524 109598
rect 202472 109534 202524 109540
rect 201656 102662 201684 109534
rect 201644 102656 201696 102662
rect 201644 102598 201696 102604
rect 202840 102656 202892 102662
rect 202840 102598 202892 102604
rect 202472 102588 202524 102594
rect 202472 102530 202524 102536
rect 201644 102520 201696 102526
rect 201644 102462 201696 102468
rect 201552 101908 201604 101914
rect 201552 101850 201604 101856
rect 201302 99726 201500 99754
rect 201656 99740 201684 102462
rect 202104 102044 202156 102050
rect 202104 101986 202156 101992
rect 202116 99740 202144 101986
rect 202484 99740 202512 102530
rect 202852 99740 202880 102598
rect 203128 102526 203156 112918
rect 203772 112674 203800 112918
rect 203220 112646 203800 112674
rect 203116 102520 203168 102526
rect 203116 102462 203168 102468
rect 203220 102050 203248 112646
rect 203760 109864 203812 109870
rect 203760 109806 203812 109812
rect 203772 102662 203800 109806
rect 204692 109598 204720 112932
rect 205336 109870 205364 112932
rect 205324 109864 205376 109870
rect 205324 109806 205376 109812
rect 205324 109728 205376 109734
rect 205324 109670 205376 109676
rect 205140 109660 205192 109666
rect 205140 109602 205192 109608
rect 203852 109592 203904 109598
rect 203852 109534 203904 109540
rect 204680 109592 204732 109598
rect 204680 109534 204732 109540
rect 203760 102656 203812 102662
rect 203760 102598 203812 102604
rect 203864 102594 203892 109534
rect 204864 102656 204916 102662
rect 204864 102598 204916 102604
rect 203852 102588 203904 102594
rect 203852 102530 203904 102536
rect 204036 102588 204088 102594
rect 204036 102530 204088 102536
rect 203300 102520 203352 102526
rect 203300 102462 203352 102468
rect 203208 102044 203260 102050
rect 203208 101986 203260 101992
rect 203312 99740 203340 102462
rect 203668 102180 203720 102186
rect 203668 102122 203720 102128
rect 203680 99740 203708 102122
rect 204048 99740 204076 102530
rect 204496 101704 204548 101710
rect 204496 101646 204548 101652
rect 204508 99740 204536 101646
rect 204876 99740 204904 102598
rect 205152 102526 205180 109602
rect 205140 102520 205192 102526
rect 205140 102462 205192 102468
rect 205232 102452 205284 102458
rect 205232 102394 205284 102400
rect 205244 99740 205272 102394
rect 205336 102186 205364 109670
rect 205888 109666 205916 112932
rect 206440 109734 206468 112932
rect 206428 109728 206480 109734
rect 206428 109670 206480 109676
rect 205876 109660 205928 109666
rect 205876 109602 205928 109608
rect 206992 109598 207020 112932
rect 207268 112918 207558 112946
rect 205416 109592 205468 109598
rect 205416 109534 205468 109540
rect 206980 109592 207032 109598
rect 206980 109534 207032 109540
rect 205428 102594 205456 109534
rect 205416 102588 205468 102594
rect 205416 102530 205468 102536
rect 206428 102384 206480 102390
rect 206428 102326 206480 102332
rect 205324 102180 205376 102186
rect 205324 102122 205376 102128
rect 205692 101636 205744 101642
rect 205692 101578 205744 101584
rect 205704 99740 205732 101578
rect 206060 101500 206112 101506
rect 206060 101442 206112 101448
rect 206072 99740 206100 101442
rect 206440 99740 206468 102326
rect 206888 101840 206940 101846
rect 206888 101782 206940 101788
rect 206900 99740 206928 101782
rect 207268 101710 207296 112918
rect 207636 112674 207664 113054
rect 208754 112918 208860 112946
rect 207360 112646 207664 112674
rect 207360 102662 207388 112646
rect 208268 110340 208320 110346
rect 208268 110282 208320 110288
rect 208176 109728 208228 109734
rect 208176 109670 208228 109676
rect 207348 102656 207400 102662
rect 207348 102598 207400 102604
rect 207256 101704 207308 101710
rect 207256 101646 207308 101652
rect 208188 101574 208216 109670
rect 207624 101568 207676 101574
rect 207624 101510 207676 101516
rect 208176 101568 208228 101574
rect 208176 101510 208228 101516
rect 207256 101432 207308 101438
rect 207256 101374 207308 101380
rect 207268 99740 207296 101374
rect 207636 99740 207664 101510
rect 208084 101364 208136 101370
rect 208084 101306 208136 101312
rect 208096 99740 208124 101306
rect 208280 99754 208308 110282
rect 208544 109660 208596 109666
rect 208544 109602 208596 109608
rect 208360 109592 208412 109598
rect 208360 109534 208412 109540
rect 208372 101438 208400 109534
rect 208360 101432 208412 101438
rect 208360 101374 208412 101380
rect 208556 101370 208584 109602
rect 208636 107552 208688 107558
rect 208636 107494 208688 107500
rect 208648 101506 208676 107494
rect 208832 102458 208860 112918
rect 208924 112918 209306 112946
rect 209568 112918 209858 112946
rect 210120 112918 210410 112946
rect 210672 112918 211054 112946
rect 208820 102452 208872 102458
rect 208820 102394 208872 102400
rect 208820 102248 208872 102254
rect 208820 102190 208872 102196
rect 208636 101500 208688 101506
rect 208636 101442 208688 101448
rect 208544 101364 208596 101370
rect 208544 101306 208596 101312
rect 208280 99726 208478 99754
rect 208832 99740 208860 102190
rect 208924 101642 208952 112918
rect 209568 107558 209596 112918
rect 209556 107552 209608 107558
rect 209556 107494 209608 107500
rect 210016 107552 210068 107558
rect 210016 107494 210068 107500
rect 209280 102112 209332 102118
rect 209280 102054 209332 102060
rect 208912 101636 208964 101642
rect 208912 101578 208964 101584
rect 209292 99740 209320 102054
rect 209648 101976 209700 101982
rect 209648 101918 209700 101924
rect 209660 99740 209688 101918
rect 210028 101846 210056 107494
rect 210120 102390 210148 112918
rect 210672 107558 210700 112918
rect 211592 109598 211620 112932
rect 212144 109734 212172 112932
rect 212132 109728 212184 109734
rect 212132 109670 212184 109676
rect 212696 109666 212724 112932
rect 213248 110346 213276 112932
rect 213340 112918 213906 112946
rect 213236 110340 213288 110346
rect 213236 110282 213288 110288
rect 212684 109660 212736 109666
rect 212684 109602 212736 109608
rect 211580 109592 211632 109598
rect 211580 109534 211632 109540
rect 210660 107552 210712 107558
rect 213340 107506 213368 112918
rect 213512 109660 213564 109666
rect 213512 109602 213564 109608
rect 213420 109592 213472 109598
rect 213420 109534 213472 109540
rect 210660 107494 210712 107500
rect 212880 107478 213368 107506
rect 210108 102384 210160 102390
rect 210108 102326 210160 102332
rect 212880 102254 212908 107478
rect 212868 102248 212920 102254
rect 212868 102190 212920 102196
rect 213432 102118 213460 109534
rect 213420 102112 213472 102118
rect 213420 102054 213472 102060
rect 213524 101982 213552 109602
rect 214444 109598 214472 112932
rect 214996 109666 215024 112932
rect 215548 110278 215576 112932
rect 215536 110272 215588 110278
rect 215536 110214 215588 110220
rect 214984 109660 215036 109666
rect 214984 109602 215036 109608
rect 214432 109592 214484 109598
rect 214432 109534 214484 109540
rect 213512 101976 213564 101982
rect 213512 101918 213564 101924
rect 210016 101840 210068 101846
rect 210016 101782 210068 101788
rect 220962 100584 221018 100593
rect 220962 100519 221018 100528
rect 194756 99590 194862 99618
rect 191982 98816 192038 98825
rect 191982 98751 192038 98760
rect 183610 98000 183666 98009
rect 183610 97935 183666 97944
rect 220976 97154 221004 100519
rect 212316 97148 212368 97154
rect 212316 97090 212368 97096
rect 220964 97148 221016 97154
rect 220964 97090 221016 97096
rect 209830 96912 209886 96921
rect 209752 96870 209830 96898
rect 183518 96776 183574 96785
rect 183518 96711 183574 96720
rect 191982 94736 192038 94745
rect 191982 94671 192038 94680
rect 191996 94434 192024 94671
rect 188580 94428 188632 94434
rect 188580 94370 188632 94376
rect 191984 94428 192036 94434
rect 191984 94370 192036 94376
rect 183426 93104 183482 93113
rect 183426 93039 183482 93048
rect 183150 91880 183206 91889
rect 183150 91815 183206 91824
rect 183058 90656 183114 90665
rect 183058 90591 183114 90600
rect 188592 90218 188620 94370
rect 191154 92832 191210 92841
rect 191154 92767 191210 92776
rect 190786 90792 190842 90801
rect 190786 90727 190842 90736
rect 182876 90212 182928 90218
rect 182876 90154 182928 90160
rect 188580 90212 188632 90218
rect 188580 90154 188632 90160
rect 182888 89441 182916 90154
rect 182874 89432 182930 89441
rect 182874 89367 182930 89376
rect 183520 88852 183572 88858
rect 183520 88794 183572 88800
rect 183532 88217 183560 88794
rect 183518 88208 183574 88217
rect 183518 88143 183574 88152
rect 190800 87498 190828 90727
rect 191168 88858 191196 92767
rect 191156 88852 191208 88858
rect 191156 88794 191208 88800
rect 191706 88752 191762 88761
rect 191706 88687 191762 88696
rect 183704 87492 183756 87498
rect 183704 87434 183756 87440
rect 190788 87492 190840 87498
rect 190788 87434 190840 87440
rect 183716 87129 183744 87434
rect 183702 87120 183758 87129
rect 183702 87055 183758 87064
rect 191614 86848 191670 86857
rect 191614 86783 191670 86792
rect 183704 86064 183756 86070
rect 183704 86006 183756 86012
rect 183716 85905 183744 86006
rect 183702 85896 183758 85905
rect 183702 85831 183758 85840
rect 182508 84704 182560 84710
rect 182508 84646 182560 84652
rect 183702 84672 183758 84681
rect 182520 83457 182548 84646
rect 191628 84642 191656 86783
rect 191720 86070 191748 88687
rect 191708 86064 191760 86070
rect 191708 86006 191760 86012
rect 191982 84808 192038 84817
rect 191982 84743 192038 84752
rect 191996 84710 192024 84743
rect 191984 84704 192036 84710
rect 191984 84646 192036 84652
rect 183702 84607 183704 84616
rect 183756 84607 183758 84616
rect 191616 84636 191668 84642
rect 183704 84578 183756 84584
rect 191616 84578 191668 84584
rect 182506 83448 182562 83457
rect 182506 83383 182562 83392
rect 191982 82768 192038 82777
rect 191982 82703 192038 82712
rect 191996 82670 192024 82703
rect 183704 82664 183756 82670
rect 183704 82606 183756 82612
rect 191984 82664 192036 82670
rect 191984 82606 192036 82612
rect 183716 82233 183744 82606
rect 183702 82224 183758 82233
rect 183702 82159 183758 82168
rect 183244 81304 183296 81310
rect 183244 81246 183296 81252
rect 191892 81304 191944 81310
rect 191892 81246 191944 81252
rect 183256 81009 183284 81246
rect 183242 81000 183298 81009
rect 183242 80935 183298 80944
rect 191904 80873 191932 81246
rect 191890 80864 191946 80873
rect 191890 80799 191946 80808
rect 136876 80556 136928 80562
rect 136876 80498 136928 80504
rect 136888 80465 136916 80498
rect 136874 80456 136930 80465
rect 136874 80391 136930 80400
rect 183702 79776 183758 79785
rect 183702 79711 183758 79720
rect 183716 79270 183744 79711
rect 183704 79264 183756 79270
rect 183704 79206 183756 79212
rect 191984 79196 192036 79202
rect 191984 79138 192036 79144
rect 191996 78833 192024 79138
rect 191982 78824 192038 78833
rect 191982 78759 192038 78768
rect 183518 78552 183574 78561
rect 183518 78487 183574 78496
rect 183532 77910 183560 78487
rect 183520 77904 183572 77910
rect 183520 77846 183572 77852
rect 191984 77904 192036 77910
rect 191984 77846 192036 77852
rect 183058 77328 183114 77337
rect 183058 77263 183114 77272
rect 183072 76482 183100 77263
rect 191996 76793 192024 77846
rect 209752 76906 209780 96870
rect 209830 96847 209886 96856
rect 212328 96513 212356 97090
rect 212314 96504 212370 96513
rect 212314 96439 212370 96448
rect 212130 89840 212186 89849
rect 212130 89775 212186 89784
rect 212038 83176 212094 83185
rect 212038 83111 212094 83120
rect 209830 76920 209886 76929
rect 209752 76878 209830 76906
rect 209830 76855 209886 76864
rect 191982 76784 192038 76793
rect 191982 76719 192038 76728
rect 183060 76476 183112 76482
rect 183060 76418 183112 76424
rect 185176 76476 185228 76482
rect 185176 76418 185228 76424
rect 183242 76104 183298 76113
rect 183242 76039 183298 76048
rect 183256 75122 183284 76039
rect 183244 75116 183296 75122
rect 183244 75058 183296 75064
rect 185188 75054 185216 76418
rect 186188 75116 186240 75122
rect 186188 75058 186240 75064
rect 185176 75048 185228 75054
rect 185176 74990 185228 74996
rect 183702 74880 183758 74889
rect 183702 74815 183758 74824
rect 183716 73898 183744 74815
rect 183704 73892 183756 73898
rect 183704 73834 183756 73840
rect 183702 73792 183758 73801
rect 183702 73727 183704 73736
rect 183756 73727 183758 73736
rect 183704 73698 183756 73704
rect 186200 73694 186228 75058
rect 191524 75048 191576 75054
rect 191524 74990 191576 74996
rect 191536 74753 191564 74990
rect 191522 74744 191578 74753
rect 191522 74679 191578 74688
rect 188488 73756 188540 73762
rect 188488 73698 188540 73704
rect 190788 73756 190840 73762
rect 190788 73698 190840 73704
rect 186188 73688 186240 73694
rect 186188 73630 186240 73636
rect 183702 72568 183758 72577
rect 183758 72526 183836 72554
rect 183702 72503 183758 72512
rect 183702 71344 183758 71353
rect 183702 71279 183758 71288
rect 183716 70974 183744 71279
rect 183704 70968 183756 70974
rect 183704 70910 183756 70916
rect 128504 70220 128556 70226
rect 128504 70162 128556 70168
rect 133380 70220 133432 70226
rect 133380 70162 133432 70168
rect 136876 70220 136928 70226
rect 136876 70162 136928 70168
rect 128516 69857 128544 70162
rect 128502 69848 128558 69857
rect 128502 69783 128558 69792
rect 106608 68180 106660 68186
rect 106608 68122 106660 68128
rect 106620 67953 106648 68122
rect 106606 67944 106662 67953
rect 106606 67879 106662 67888
rect 136888 66593 136916 70162
rect 182874 70120 182930 70129
rect 182874 70055 182930 70064
rect 182888 69954 182916 70055
rect 182876 69948 182928 69954
rect 182876 69890 182928 69896
rect 183058 68896 183114 68905
rect 183058 68831 183114 68840
rect 136874 66584 136930 66593
rect 136874 66519 136930 66528
rect 137978 66584 138034 66593
rect 137978 66519 138034 66528
rect 106514 65632 106570 65641
rect 106514 65567 106570 65576
rect 104492 63692 104544 63698
rect 104492 63634 104544 63640
rect 106608 63692 106660 63698
rect 106608 63634 106660 63640
rect 106620 63329 106648 63634
rect 106606 63320 106662 63329
rect 106606 63255 106662 63264
rect 105320 61380 105372 61386
rect 105320 61322 105372 61328
rect 104400 61244 104452 61250
rect 99340 50160 99392 50166
rect 99340 50102 99392 50108
rect 99536 50098 99564 61238
rect 104400 61186 104452 61192
rect 100258 59920 100314 59929
rect 100258 59855 100314 59864
rect 100272 50234 100300 59855
rect 100260 50228 100312 50234
rect 100260 50170 100312 50176
rect 104768 50228 104820 50234
rect 104768 50170 104820 50176
rect 99524 50092 99576 50098
rect 99524 50034 99576 50040
rect 99248 49820 99300 49826
rect 99248 49762 99300 49768
rect 99156 49684 99208 49690
rect 99156 49626 99208 49632
rect 99064 49616 99116 49622
rect 99064 49558 99116 49564
rect 98972 49548 99024 49554
rect 98972 49490 99024 49496
rect 90692 48936 90744 48942
rect 90692 48878 90744 48884
rect 104216 48936 104268 48942
rect 104216 48878 104268 48884
rect 79282 46864 79338 46873
rect 79282 46799 79338 46808
rect 73394 46592 73450 46601
rect 73394 46527 73450 46536
rect 73408 44810 73436 46527
rect 76338 46456 76394 46465
rect 76338 46391 76394 46400
rect 74866 46320 74922 46329
rect 74866 46255 74922 46264
rect 74880 44810 74908 46255
rect 76352 44810 76380 46391
rect 77810 46184 77866 46193
rect 77810 46119 77866 46128
rect 77824 44810 77852 46119
rect 79296 44810 79324 46799
rect 80754 46728 80810 46737
rect 80754 46663 80810 46672
rect 80768 44810 80796 46663
rect 85722 46320 85778 46329
rect 82964 46284 83016 46290
rect 85722 46255 85778 46264
rect 82964 46226 83016 46232
rect 82976 44810 83004 46226
rect 84068 46216 84120 46222
rect 84068 46158 84120 46164
rect 61356 44782 61692 44810
rect 62828 44782 63164 44810
rect 64300 44782 64636 44810
rect 65772 44782 66108 44810
rect 67336 44782 67672 44810
rect 68808 44782 69144 44810
rect 70556 44782 70616 44810
rect 73408 44782 73652 44810
rect 74880 44782 75124 44810
rect 76352 44782 76688 44810
rect 77824 44782 78160 44810
rect 79296 44782 79632 44810
rect 80768 44782 81104 44810
rect 82668 44782 83004 44810
rect 84080 44810 84108 46158
rect 85736 44810 85764 46255
rect 87102 46184 87158 46193
rect 87102 46119 87158 46128
rect 88944 46148 88996 46154
rect 84080 44782 84140 44810
rect 85612 44782 85764 44810
rect 58308 44720 58360 44726
rect 58308 44662 58360 44668
rect 87116 44674 87144 46119
rect 88944 46090 88996 46096
rect 88956 44810 88984 46090
rect 88648 44782 88984 44810
rect 51316 44652 51368 44658
rect 51316 44594 51368 44600
rect 58216 44652 58268 44658
rect 58216 44594 58268 44600
rect 58228 44425 58256 44594
rect 58214 44416 58270 44425
rect 58214 44351 58270 44360
rect 51222 44144 51278 44153
rect 51222 44079 51278 44088
rect 51236 43366 51264 44079
rect 58320 43881 58348 44662
rect 87116 44646 87176 44674
rect 90324 44584 90376 44590
rect 90120 44532 90324 44538
rect 90120 44526 90376 44532
rect 90120 44510 90364 44526
rect 90704 44522 90732 48878
rect 104228 46700 104256 48878
rect 104780 46700 104808 50170
rect 105332 46700 105360 61322
rect 107160 61244 107212 61250
rect 107160 61186 107212 61192
rect 107172 61017 107200 61186
rect 107158 61008 107214 61017
rect 107158 60943 107214 60952
rect 109276 57232 109328 57238
rect 109276 57174 109328 57180
rect 109184 57164 109236 57170
rect 109184 57106 109236 57112
rect 105872 50160 105924 50166
rect 105872 50102 105924 50108
rect 105884 46700 105912 50102
rect 106424 50092 106476 50098
rect 106424 50034 106476 50040
rect 106436 46700 106464 50034
rect 106976 49820 107028 49826
rect 106976 49762 107028 49768
rect 106988 46700 107016 49762
rect 107528 49684 107580 49690
rect 107528 49626 107580 49632
rect 107540 46700 107568 49626
rect 108080 49616 108132 49622
rect 108080 49558 108132 49564
rect 108092 46700 108120 49558
rect 108632 49548 108684 49554
rect 108632 49490 108684 49496
rect 108644 46700 108672 49490
rect 109196 46700 109224 57106
rect 109288 46850 109316 57174
rect 110116 57170 110144 59892
rect 110484 57238 110512 59892
rect 110760 59878 110866 59906
rect 111128 59878 111326 59906
rect 110472 57232 110524 57238
rect 110472 57174 110524 57180
rect 110104 57164 110156 57170
rect 110104 57106 110156 57112
rect 110760 57050 110788 59878
rect 111128 58546 111156 59878
rect 110576 57022 110788 57050
rect 110944 58518 111156 58546
rect 109288 46822 109500 46850
rect 109472 46714 109500 46822
rect 110576 46714 110604 57022
rect 110944 54874 110972 58518
rect 111680 57170 111708 59892
rect 112062 59878 112260 59906
rect 111116 57164 111168 57170
rect 111116 57106 111168 57112
rect 111668 57164 111720 57170
rect 111668 57106 111720 57112
rect 110760 54846 110972 54874
rect 110760 46970 110788 54846
rect 110748 46964 110800 46970
rect 110748 46906 110800 46912
rect 110932 46964 110984 46970
rect 110932 46906 110984 46912
rect 110944 46714 110972 46906
rect 109472 46686 109762 46714
rect 110314 46686 110604 46714
rect 110866 46686 110972 46714
rect 111128 46714 111156 57106
rect 112232 46714 112260 59878
rect 112404 58592 112456 58598
rect 112404 58534 112456 58540
rect 112312 50296 112364 50302
rect 112312 50238 112364 50244
rect 111128 46686 111510 46714
rect 112062 46686 112260 46714
rect 112324 46714 112352 50238
rect 112416 46986 112444 58534
rect 112508 50302 112536 59892
rect 112876 58598 112904 59892
rect 112864 58592 112916 58598
rect 112864 58534 112916 58540
rect 113244 57186 113272 59892
rect 113718 59878 113824 59906
rect 113244 57158 113548 57186
rect 112496 50296 112548 50302
rect 112496 50238 112548 50244
rect 112416 46958 112904 46986
rect 112876 46714 112904 46958
rect 113520 46714 113548 57158
rect 113796 46714 113824 59878
rect 114072 57782 114100 59892
rect 114060 57776 114112 57782
rect 114060 57718 114112 57724
rect 114440 57238 114468 59892
rect 114428 57232 114480 57238
rect 114428 57174 114480 57180
rect 114900 57170 114928 59892
rect 114980 57776 115032 57782
rect 114980 57718 115032 57724
rect 114888 57164 114940 57170
rect 114888 57106 114940 57112
rect 114992 46714 115020 57718
rect 115268 57306 115296 59892
rect 115650 59878 116032 59906
rect 115256 57300 115308 57306
rect 115256 57242 115308 57248
rect 115348 57232 115400 57238
rect 115348 57174 115400 57180
rect 112324 46686 112614 46714
rect 112876 46686 113166 46714
rect 113520 46686 113718 46714
rect 113796 46686 114270 46714
rect 114822 46686 115020 46714
rect 115360 46700 115388 57174
rect 116004 57170 116032 59878
rect 116096 57646 116124 59892
rect 116084 57640 116136 57646
rect 116084 57582 116136 57588
rect 116268 57300 116320 57306
rect 116268 57242 116320 57248
rect 115532 57164 115584 57170
rect 115532 57106 115584 57112
rect 115992 57164 116044 57170
rect 115992 57106 116044 57112
rect 115544 46714 115572 57106
rect 116280 46714 116308 57242
rect 116464 57238 116492 59892
rect 116832 57714 116860 59892
rect 116820 57708 116872 57714
rect 116820 57650 116872 57656
rect 116452 57232 116504 57238
rect 116452 57174 116504 57180
rect 117292 57170 117320 59892
rect 117660 57306 117688 59892
rect 117740 57640 117792 57646
rect 117740 57582 117792 57588
rect 117648 57300 117700 57306
rect 117648 57242 117700 57248
rect 116636 57164 116688 57170
rect 116636 57106 116688 57112
rect 117280 57164 117332 57170
rect 117280 57106 117332 57112
rect 116648 46714 116676 57106
rect 117752 46714 117780 57582
rect 118120 57510 118148 59892
rect 118384 57708 118436 57714
rect 118384 57650 118436 57656
rect 118108 57504 118160 57510
rect 118108 57446 118160 57452
rect 118396 57322 118424 57650
rect 118488 57442 118516 59892
rect 118856 57578 118884 59892
rect 118844 57572 118896 57578
rect 118844 57514 118896 57520
rect 118476 57436 118528 57442
rect 118476 57378 118528 57384
rect 118396 57294 118516 57322
rect 119316 57306 119344 59892
rect 118108 57232 118160 57238
rect 118108 57174 118160 57180
rect 118120 48346 118148 57174
rect 118200 57164 118252 57170
rect 118200 57106 118252 57112
rect 118212 50234 118240 57106
rect 118200 50228 118252 50234
rect 118200 50170 118252 50176
rect 118120 48318 118240 48346
rect 115544 46686 115926 46714
rect 116280 46686 116478 46714
rect 116648 46686 117030 46714
rect 117582 46686 117780 46714
rect 118212 46700 118240 48318
rect 118488 46714 118516 57294
rect 118844 57300 118896 57306
rect 118844 57242 118896 57248
rect 119304 57300 119356 57306
rect 119304 57242 119356 57248
rect 118856 49146 118884 57242
rect 119684 57170 119712 59892
rect 120052 57238 120080 59892
rect 120512 58122 120540 59892
rect 120500 58116 120552 58122
rect 120500 58058 120552 58064
rect 120880 57986 120908 59892
rect 121248 58394 121276 59892
rect 121236 58388 121288 58394
rect 121236 58330 121288 58336
rect 120868 57980 120920 57986
rect 120868 57922 120920 57928
rect 121236 57572 121288 57578
rect 121236 57514 121288 57520
rect 120500 57504 120552 57510
rect 120500 57446 120552 57452
rect 120040 57232 120092 57238
rect 120040 57174 120092 57180
rect 119672 57164 119724 57170
rect 119672 57106 119724 57112
rect 119304 50228 119356 50234
rect 119304 50170 119356 50176
rect 118844 49140 118896 49146
rect 118844 49082 118896 49088
rect 118488 46686 118778 46714
rect 119316 46700 119344 50170
rect 119856 49140 119908 49146
rect 119856 49082 119908 49088
rect 119868 46700 119896 49082
rect 120512 46714 120540 57446
rect 120776 57436 120828 57442
rect 120776 57378 120828 57384
rect 120434 46686 120540 46714
rect 120788 46714 120816 57378
rect 121052 57300 121104 57306
rect 121052 57242 121104 57248
rect 120960 57164 121012 57170
rect 120960 57106 121012 57112
rect 120972 50234 121000 57106
rect 120960 50228 121012 50234
rect 120960 50170 121012 50176
rect 121064 49758 121092 57242
rect 121144 57232 121196 57238
rect 121144 57174 121196 57180
rect 121156 50098 121184 57174
rect 121144 50092 121196 50098
rect 121144 50034 121196 50040
rect 121052 49752 121104 49758
rect 121052 49694 121104 49700
rect 121248 46714 121276 57514
rect 121708 57442 121736 59892
rect 122076 57850 122104 59892
rect 122444 58326 122472 59892
rect 122432 58320 122484 58326
rect 122432 58262 122484 58268
rect 122064 57844 122116 57850
rect 122064 57786 122116 57792
rect 122904 57578 122932 59892
rect 123272 58258 123300 59892
rect 123260 58252 123312 58258
rect 123260 58194 123312 58200
rect 123260 58116 123312 58122
rect 123260 58058 123312 58064
rect 122892 57572 122944 57578
rect 122892 57514 122944 57520
rect 121696 57436 121748 57442
rect 121696 57378 121748 57384
rect 122616 50228 122668 50234
rect 122616 50170 122668 50176
rect 122064 49752 122116 49758
rect 122064 49694 122116 49700
rect 120788 46686 120986 46714
rect 121248 46686 121538 46714
rect 122076 46700 122104 49694
rect 122628 46700 122656 50170
rect 123168 50092 123220 50098
rect 123168 50034 123220 50040
rect 123180 46700 123208 50034
rect 123272 46714 123300 58058
rect 123444 57980 123496 57986
rect 123444 57922 123496 57928
rect 123456 47802 123484 57922
rect 123640 57306 123668 59892
rect 123720 58388 123772 58394
rect 123720 58330 123772 58336
rect 123628 57300 123680 57306
rect 123628 57242 123680 57248
rect 123732 50234 123760 58330
rect 124100 57510 124128 59892
rect 124088 57504 124140 57510
rect 124088 57446 124140 57452
rect 124468 57374 124496 59892
rect 124456 57368 124508 57374
rect 124456 57310 124508 57316
rect 124836 57238 124864 59892
rect 125100 58320 125152 58326
rect 125100 58262 125152 58268
rect 124916 57436 124968 57442
rect 124916 57378 124968 57384
rect 124824 57232 124876 57238
rect 124824 57174 124876 57180
rect 123720 50228 123772 50234
rect 123720 50170 123772 50176
rect 124824 50228 124876 50234
rect 124824 50170 124876 50176
rect 123456 47774 123944 47802
rect 123916 46714 123944 47774
rect 123272 46686 123746 46714
rect 123916 46686 124298 46714
rect 124836 46700 124864 50170
rect 124928 46850 124956 57378
rect 125112 49554 125140 58262
rect 125192 57844 125244 57850
rect 125192 57786 125244 57792
rect 125204 49962 125232 57786
rect 125296 57714 125324 59892
rect 125284 57708 125336 57714
rect 125284 57650 125336 57656
rect 125284 57572 125336 57578
rect 125284 57514 125336 57520
rect 125192 49956 125244 49962
rect 125192 49898 125244 49904
rect 125100 49548 125152 49554
rect 125100 49490 125152 49496
rect 125296 49214 125324 57514
rect 125664 57170 125692 59892
rect 137992 59890 138020 66519
rect 182690 60464 182746 60473
rect 182690 60399 182692 60408
rect 182744 60399 182746 60408
rect 182692 60370 182744 60376
rect 137980 59884 138032 59890
rect 137980 59826 138032 59832
rect 138164 59884 138216 59890
rect 138164 59826 138216 59832
rect 127308 58252 127360 58258
rect 127308 58194 127360 58200
rect 127216 57300 127268 57306
rect 127216 57242 127268 57248
rect 125652 57164 125704 57170
rect 125652 57106 125704 57112
rect 127228 50438 127256 57242
rect 127216 50432 127268 50438
rect 127216 50374 127268 50380
rect 126020 49956 126072 49962
rect 126020 49898 126072 49904
rect 125284 49208 125336 49214
rect 125284 49150 125336 49156
rect 124928 46822 125140 46850
rect 125112 46714 125140 46822
rect 125112 46686 125494 46714
rect 126032 46700 126060 49898
rect 126572 49548 126624 49554
rect 126572 49490 126624 49496
rect 126584 46700 126612 49490
rect 127124 49208 127176 49214
rect 127124 49150 127176 49156
rect 127136 46700 127164 49150
rect 127320 46714 127348 58194
rect 129976 57708 130028 57714
rect 129976 57650 130028 57656
rect 128780 57504 128832 57510
rect 128780 57446 128832 57452
rect 127860 50432 127912 50438
rect 127860 50374 127912 50380
rect 127872 46714 127900 50374
rect 127320 46686 127702 46714
rect 127872 46686 128254 46714
rect 128792 46700 128820 57446
rect 128872 57368 128924 57374
rect 128872 57310 128924 57316
rect 128884 46714 128912 57310
rect 129516 57232 129568 57238
rect 129516 57174 129568 57180
rect 129528 46714 129556 57174
rect 129988 46714 130016 57650
rect 130068 57164 130120 57170
rect 130068 57106 130120 57112
rect 130080 47122 130108 57106
rect 138176 55742 138204 59826
rect 156576 58462 156604 59892
rect 163200 58530 163228 59892
rect 163188 58524 163240 58530
rect 163188 58466 163240 58472
rect 156564 58456 156616 58462
rect 156564 58398 156616 58404
rect 169916 57850 169944 59892
rect 156104 57844 156156 57850
rect 156104 57786 156156 57792
rect 169904 57844 169956 57850
rect 169904 57786 169956 57792
rect 138164 55736 138216 55742
rect 138164 55678 138216 55684
rect 138348 55736 138400 55742
rect 138348 55678 138400 55684
rect 130080 47094 130568 47122
rect 130540 46714 130568 47094
rect 128884 46686 129358 46714
rect 129528 46686 129910 46714
rect 129988 46686 130462 46714
rect 130540 46686 131014 46714
rect 134576 46556 134628 46562
rect 134576 46498 134628 46504
rect 93360 46284 93412 46290
rect 93360 46226 93412 46232
rect 90416 44516 90468 44522
rect 90416 44458 90468 44464
rect 90692 44516 90744 44522
rect 90692 44458 90744 44464
rect 58306 43872 58362 43881
rect 58306 43807 58362 43816
rect 56744 43564 56796 43570
rect 56744 43506 56796 43512
rect 51224 43360 51276 43366
rect 51224 43302 51276 43308
rect 56652 43360 56704 43366
rect 56652 43302 56704 43308
rect 56664 43230 56692 43302
rect 56652 43224 56704 43230
rect 56652 43166 56704 43172
rect 56756 43162 56784 43506
rect 58216 43224 58268 43230
rect 58214 43192 58216 43201
rect 58268 43192 58270 43201
rect 56744 43156 56796 43162
rect 58214 43127 58270 43136
rect 58308 43156 58360 43162
rect 56744 43098 56796 43104
rect 58308 43098 58360 43104
rect 58320 42657 58348 43098
rect 58306 42648 58362 42657
rect 58216 42612 58268 42618
rect 58306 42583 58362 42592
rect 58216 42554 58268 42560
rect 51130 42376 51186 42385
rect 51130 42311 51186 42320
rect 51144 42074 51172 42311
rect 58228 42113 58256 42554
rect 51222 42104 51278 42113
rect 51132 42068 51184 42074
rect 51222 42039 51278 42048
rect 58214 42104 58270 42113
rect 58214 42039 58270 42048
rect 51132 42010 51184 42016
rect 51236 42006 51264 42039
rect 51224 42000 51276 42006
rect 51224 41942 51276 41948
rect 58216 41932 58268 41938
rect 58216 41874 58268 41880
rect 58228 41433 58256 41874
rect 58308 41796 58360 41802
rect 58308 41738 58360 41744
rect 58214 41424 58270 41433
rect 58214 41359 58270 41368
rect 51130 41152 51186 41161
rect 51130 41087 51186 41096
rect 51144 40646 51172 41087
rect 58320 40889 58348 41738
rect 51222 40880 51278 40889
rect 51222 40815 51278 40824
rect 58306 40880 58362 40889
rect 58306 40815 58362 40824
rect 51236 40714 51264 40815
rect 51224 40708 51276 40714
rect 51224 40650 51276 40656
rect 55732 40708 55784 40714
rect 55732 40650 55784 40656
rect 51132 40640 51184 40646
rect 51132 40582 51184 40588
rect 55744 40170 55772 40650
rect 56560 40640 56612 40646
rect 56560 40582 56612 40588
rect 56572 40442 56600 40582
rect 56560 40436 56612 40442
rect 56560 40378 56612 40384
rect 58216 40436 58268 40442
rect 58216 40378 58268 40384
rect 58228 40209 58256 40378
rect 58214 40200 58270 40209
rect 55732 40164 55784 40170
rect 58214 40135 58270 40144
rect 58308 40164 58360 40170
rect 55732 40106 55784 40112
rect 58308 40106 58360 40112
rect 51130 39928 51186 39937
rect 51130 39863 51186 39872
rect 51144 39286 51172 39863
rect 58320 39665 58348 40106
rect 58306 39656 58362 39665
rect 58306 39591 58362 39600
rect 51222 39520 51278 39529
rect 51222 39455 51278 39464
rect 51132 39280 51184 39286
rect 51132 39222 51184 39228
rect 51236 39218 51264 39455
rect 51224 39212 51276 39218
rect 51224 39154 51276 39160
rect 58216 39144 58268 39150
rect 58214 39112 58216 39121
rect 58268 39112 58270 39121
rect 58214 39047 58270 39056
rect 58400 39076 58452 39082
rect 58400 39018 58452 39024
rect 51222 38840 51278 38849
rect 51222 38775 51278 38784
rect 51236 38470 51264 38775
rect 51224 38464 51276 38470
rect 51224 38406 51276 38412
rect 58308 38464 58360 38470
rect 58412 38441 58440 39018
rect 58308 38406 58360 38412
rect 58398 38432 58454 38441
rect 51130 38160 51186 38169
rect 51130 38095 51186 38104
rect 51144 37926 51172 38095
rect 51132 37920 51184 37926
rect 58320 37897 58348 38406
rect 58398 38367 58454 38376
rect 58400 37920 58452 37926
rect 51132 37862 51184 37868
rect 51222 37888 51278 37897
rect 58306 37888 58362 37897
rect 51222 37823 51224 37832
rect 51276 37823 51278 37832
rect 58216 37852 58268 37858
rect 51224 37794 51276 37800
rect 58400 37862 58452 37868
rect 58306 37823 58362 37832
rect 58216 37794 58268 37800
rect 51130 36936 51186 36945
rect 51130 36871 51186 36880
rect 51144 36498 51172 36871
rect 58228 36673 58256 37794
rect 58412 37217 58440 37862
rect 58398 37208 58454 37217
rect 58398 37143 58454 37152
rect 51222 36664 51278 36673
rect 51222 36599 51278 36608
rect 58214 36664 58270 36673
rect 58214 36599 58270 36608
rect 51236 36566 51264 36599
rect 51224 36560 51276 36566
rect 51224 36502 51276 36508
rect 58308 36560 58360 36566
rect 58308 36502 58360 36508
rect 51132 36492 51184 36498
rect 51132 36434 51184 36440
rect 58216 36492 58268 36498
rect 58216 36434 58268 36440
rect 58228 36129 58256 36434
rect 58214 36120 58270 36129
rect 58214 36055 58270 36064
rect 58320 35449 58348 36502
rect 58306 35440 58362 35449
rect 58306 35375 58362 35384
rect 51222 35304 51278 35313
rect 51222 35239 51278 35248
rect 55456 35268 55508 35274
rect 51236 35138 51264 35239
rect 55456 35210 55508 35216
rect 51224 35132 51276 35138
rect 51224 35074 51276 35080
rect 55468 35002 55496 35210
rect 58308 35064 58360 35070
rect 58308 35006 58360 35012
rect 55456 34996 55508 35002
rect 55456 34938 55508 34944
rect 58216 34996 58268 35002
rect 58216 34938 58268 34944
rect 58228 34905 58256 34938
rect 58214 34896 58270 34905
rect 58214 34831 58270 34840
rect 58320 34225 58348 35006
rect 51222 34216 51278 34225
rect 51222 34151 51278 34160
rect 58306 34216 58362 34225
rect 58306 34151 58362 34160
rect 51236 34050 51264 34151
rect 51224 34044 51276 34050
rect 51224 33986 51276 33992
rect 56744 34044 56796 34050
rect 56744 33986 56796 33992
rect 51222 33808 51278 33817
rect 51222 33743 51278 33752
rect 51236 33710 51264 33743
rect 51224 33704 51276 33710
rect 51224 33646 51276 33652
rect 56008 33704 56060 33710
rect 56008 33646 56060 33652
rect 56020 33030 56048 33646
rect 56756 33506 56784 33986
rect 58214 33672 58270 33681
rect 58214 33607 58216 33616
rect 58268 33607 58270 33616
rect 58216 33578 58268 33584
rect 56744 33500 56796 33506
rect 56744 33442 56796 33448
rect 58216 33500 58268 33506
rect 58216 33442 58268 33448
rect 58228 33137 58256 33442
rect 58214 33128 58270 33137
rect 58214 33063 58270 33072
rect 56008 33024 56060 33030
rect 56008 32966 56060 32972
rect 58216 33024 58268 33030
rect 58216 32966 58268 32972
rect 58228 32457 58256 32966
rect 51222 32448 51278 32457
rect 58214 32448 58270 32457
rect 51222 32383 51224 32392
rect 51276 32383 51278 32392
rect 56744 32412 56796 32418
rect 51224 32354 51276 32360
rect 58214 32383 58270 32392
rect 56744 32354 56796 32360
rect 56652 32344 56704 32350
rect 56652 32286 56704 32292
rect 56664 32214 56692 32286
rect 56652 32208 56704 32214
rect 56652 32150 56704 32156
rect 56756 31874 56784 32354
rect 58216 32208 58268 32214
rect 58216 32150 58268 32156
rect 58228 31913 58256 32150
rect 58214 31904 58270 31913
rect 56744 31868 56796 31874
rect 58214 31839 58270 31848
rect 58308 31868 58360 31874
rect 56744 31810 56796 31816
rect 58308 31810 58360 31816
rect 51130 31632 51186 31641
rect 51130 31567 51186 31576
rect 51144 31058 51172 31567
rect 58320 31233 58348 31810
rect 51222 31224 51278 31233
rect 51222 31159 51278 31168
rect 58306 31224 58362 31233
rect 58306 31159 58362 31168
rect 51132 31052 51184 31058
rect 51132 30994 51184 31000
rect 51236 30990 51264 31159
rect 51224 30984 51276 30990
rect 51224 30926 51276 30932
rect 58216 30916 58268 30922
rect 58216 30858 58268 30864
rect 58228 30689 58256 30858
rect 58308 30780 58360 30786
rect 58308 30722 58360 30728
rect 58214 30680 58270 30689
rect 58214 30615 58270 30624
rect 51130 30408 51186 30417
rect 51130 30343 51186 30352
rect 51144 29630 51172 30343
rect 58320 30145 58348 30722
rect 58306 30136 58362 30145
rect 58306 30071 58362 30080
rect 51222 29864 51278 29873
rect 51222 29799 51278 29808
rect 51132 29624 51184 29630
rect 51132 29566 51184 29572
rect 51236 29562 51264 29799
rect 51224 29556 51276 29562
rect 51224 29498 51276 29504
rect 56652 29556 56704 29562
rect 56652 29498 56704 29504
rect 56664 29290 56692 29498
rect 58216 29488 58268 29494
rect 58214 29456 58216 29465
rect 58268 29456 58270 29465
rect 58214 29391 58270 29400
rect 56652 29284 56704 29290
rect 56652 29226 56704 29232
rect 58216 29284 58268 29290
rect 58216 29226 58268 29232
rect 51130 29184 51186 29193
rect 51130 29119 51186 29128
rect 51144 28814 51172 29119
rect 58228 28921 58256 29226
rect 58214 28912 58270 28921
rect 58214 28847 58270 28856
rect 51132 28808 51184 28814
rect 58216 28808 58268 28814
rect 51132 28750 51184 28756
rect 51222 28776 51278 28785
rect 58216 28750 58268 28756
rect 51222 28711 51278 28720
rect 51236 28610 51264 28711
rect 51224 28604 51276 28610
rect 51224 28546 51276 28552
rect 56744 28604 56796 28610
rect 56744 28546 56796 28552
rect 51222 28368 51278 28377
rect 51222 28303 51224 28312
rect 51276 28303 51278 28312
rect 56008 28332 56060 28338
rect 51224 28274 51276 28280
rect 56008 28274 56060 28280
rect 56020 27726 56048 28274
rect 56756 28134 56784 28546
rect 58228 28241 58256 28750
rect 58214 28232 58270 28241
rect 58214 28167 58270 28176
rect 56744 28128 56796 28134
rect 56744 28070 56796 28076
rect 58216 28128 58268 28134
rect 58216 28070 58268 28076
rect 56008 27720 56060 27726
rect 58228 27697 58256 28070
rect 58308 27720 58360 27726
rect 56008 27662 56060 27668
rect 58214 27688 58270 27697
rect 58308 27662 58360 27668
rect 58214 27623 58270 27632
rect 51130 27416 51186 27425
rect 51130 27351 51186 27360
rect 51144 26842 51172 27351
rect 58320 27153 58348 27662
rect 58306 27144 58362 27153
rect 58306 27079 58362 27088
rect 51222 27008 51278 27017
rect 51222 26943 51278 26952
rect 51236 26910 51264 26943
rect 51224 26904 51276 26910
rect 51224 26846 51276 26852
rect 58308 26904 58360 26910
rect 58308 26846 58360 26852
rect 51132 26836 51184 26842
rect 51132 26778 51184 26784
rect 58216 26836 58268 26842
rect 58216 26778 58268 26784
rect 58228 26473 58256 26778
rect 58214 26464 58270 26473
rect 58214 26399 58270 26408
rect 58320 25929 58348 26846
rect 58306 25920 58362 25929
rect 58306 25855 58362 25864
rect 51222 25784 51278 25793
rect 51222 25719 51278 25728
rect 51132 25612 51184 25618
rect 51132 25554 51184 25560
rect 51144 25521 51172 25554
rect 51236 25550 51264 25719
rect 59320 25612 59372 25618
rect 59320 25554 59372 25560
rect 51224 25544 51276 25550
rect 51130 25512 51186 25521
rect 51224 25486 51276 25492
rect 51130 25447 51186 25456
rect 51130 24424 51186 24433
rect 51130 24359 51186 24368
rect 51144 24122 51172 24359
rect 59332 24161 59360 25554
rect 59412 25544 59464 25550
rect 59412 25486 59464 25492
rect 59424 24705 59452 25486
rect 59504 25476 59556 25482
rect 59504 25418 59556 25424
rect 59516 25249 59544 25418
rect 59502 25240 59558 25249
rect 59502 25175 59558 25184
rect 59410 24696 59466 24705
rect 59410 24631 59466 24640
rect 51222 24152 51278 24161
rect 51132 24116 51184 24122
rect 51222 24087 51278 24096
rect 59318 24152 59374 24161
rect 59318 24087 59374 24096
rect 51132 24058 51184 24064
rect 51236 24054 51264 24087
rect 51224 24048 51276 24054
rect 51224 23990 51276 23996
rect 58216 23980 58268 23986
rect 58216 23922 58268 23928
rect 58228 23481 58256 23922
rect 58308 23912 58360 23918
rect 58308 23854 58360 23860
rect 58214 23472 58270 23481
rect 58214 23407 58270 23416
rect 58320 22937 58348 23854
rect 51222 22928 51278 22937
rect 51222 22863 51278 22872
rect 58306 22928 58362 22937
rect 58306 22863 58362 22872
rect 51236 22762 51264 22863
rect 51224 22756 51276 22762
rect 51224 22698 51276 22704
rect 55916 22756 55968 22762
rect 55916 22698 55968 22704
rect 55928 22218 55956 22698
rect 58216 22620 58268 22626
rect 58216 22562 58268 22568
rect 58228 22257 58256 22562
rect 58214 22248 58270 22257
rect 55916 22212 55968 22218
rect 58214 22183 58270 22192
rect 58308 22212 58360 22218
rect 55916 22154 55968 22160
rect 58308 22154 58360 22160
rect 51222 21976 51278 21985
rect 51222 21911 51278 21920
rect 51236 21334 51264 21911
rect 58320 21713 58348 22154
rect 58306 21704 58362 21713
rect 58306 21639 58362 21648
rect 51224 21328 51276 21334
rect 90428 21282 90456 44458
rect 92716 41932 92768 41938
rect 92716 41874 92768 41880
rect 92728 41297 92756 41874
rect 92714 41288 92770 41297
rect 92714 41223 92770 41232
rect 92716 40572 92768 40578
rect 92716 40514 92768 40520
rect 92728 40073 92756 40514
rect 92714 40064 92770 40073
rect 92714 39999 92770 40008
rect 92900 39144 92952 39150
rect 92900 39086 92952 39092
rect 92912 38305 92940 39086
rect 92898 38296 92954 38305
rect 92898 38231 92954 38240
rect 90600 37852 90652 37858
rect 90600 37794 90652 37800
rect 90612 28116 90640 37794
rect 92900 36424 92952 36430
rect 92900 36366 92952 36372
rect 92912 35993 92940 36366
rect 92898 35984 92954 35993
rect 92898 35919 92954 35928
rect 92716 30916 92768 30922
rect 92716 30858 92768 30864
rect 92728 30553 92756 30858
rect 92714 30544 92770 30553
rect 92714 30479 92770 30488
rect 92716 29420 92768 29426
rect 92716 29362 92768 29368
rect 92728 28785 92756 29362
rect 92714 28776 92770 28785
rect 92714 28711 92770 28720
rect 90692 28128 90744 28134
rect 90612 28088 90692 28116
rect 90692 28070 90744 28076
rect 92716 28060 92768 28066
rect 92716 28002 92768 28008
rect 92728 27561 92756 28002
rect 92714 27552 92770 27561
rect 92714 27487 92770 27496
rect 92900 23980 92952 23986
rect 92900 23922 92952 23928
rect 92912 23345 92940 23922
rect 92898 23336 92954 23345
rect 92898 23271 92954 23280
rect 51224 21270 51276 21276
rect 58216 21260 58268 21266
rect 90304 21254 90456 21282
rect 58216 21202 58268 21208
rect 58228 21169 58256 21202
rect 58214 21160 58270 21169
rect 58214 21095 58270 21104
rect 51038 21024 51094 21033
rect 61710 21024 61766 21033
rect 61416 20982 61710 21010
rect 51038 20959 51094 20968
rect 61710 20959 61766 20968
rect 63182 21024 63238 21033
rect 64746 21024 64802 21033
rect 63238 20982 63440 21010
rect 64452 20982 64746 21010
rect 63182 20959 63238 20968
rect 64746 20959 64802 20968
rect 65114 21024 65170 21033
rect 65170 20982 65464 21010
rect 65114 20959 65170 20968
rect 62722 20888 62778 20897
rect 62428 20846 62722 20874
rect 62722 20823 62778 20832
rect 66508 20846 66568 20874
rect 67580 20846 67824 20874
rect 50854 20480 50910 20489
rect 50854 20415 50910 20424
rect 50762 19800 50818 19809
rect 50762 19735 50818 19744
rect 50578 19256 50634 19265
rect 50578 19191 50634 19200
rect 18104 18472 18156 18478
rect 18104 18414 18156 18420
rect 60792 18336 60844 18342
rect 66508 18313 66536 20846
rect 60792 18278 60844 18284
rect 66494 18304 66550 18313
rect 54812 18268 54864 18274
rect 54812 18210 54864 18216
rect 42852 18200 42904 18206
rect 42852 18142 42904 18148
rect 36780 18064 36832 18070
rect 36780 18006 36832 18012
rect 30800 17996 30852 18002
rect 30800 17938 30852 17944
rect 18840 17928 18892 17934
rect 18840 17870 18892 17876
rect 12860 17792 12912 17798
rect 12860 17734 12912 17740
rect 12872 9304 12900 17734
rect 18852 9304 18880 17870
rect 24820 17860 24872 17866
rect 24820 17802 24872 17808
rect 24832 9304 24860 17802
rect 30812 9304 30840 17938
rect 36792 9304 36820 18006
rect 42864 9304 42892 18142
rect 48832 18132 48884 18138
rect 48832 18074 48884 18080
rect 48844 9304 48872 18074
rect 54824 9304 54852 18210
rect 60804 9304 60832 18278
rect 66494 18239 66550 18248
rect 67796 17118 67824 20846
rect 68256 20846 68592 20874
rect 69604 20846 69940 20874
rect 68256 18478 68284 20846
rect 68244 18472 68296 18478
rect 68244 18414 68296 18420
rect 69912 18410 69940 20846
rect 70648 20846 70708 20874
rect 71384 20846 71720 20874
rect 72396 20846 72732 20874
rect 73408 20846 73744 20874
rect 74788 20846 74848 20874
rect 75524 20846 75860 20874
rect 76872 20846 77208 20874
rect 69900 18404 69952 18410
rect 69900 18346 69952 18352
rect 70648 18206 70676 20846
rect 70636 18200 70688 18206
rect 70636 18142 70688 18148
rect 71384 18070 71412 20846
rect 71372 18064 71424 18070
rect 71372 18006 71424 18012
rect 72396 18002 72424 20846
rect 72384 17996 72436 18002
rect 72384 17938 72436 17944
rect 73408 17866 73436 20846
rect 74788 17934 74816 20846
rect 74776 17928 74828 17934
rect 74776 17870 74828 17876
rect 73396 17860 73448 17866
rect 73396 17802 73448 17808
rect 75524 17798 75552 20846
rect 76248 18336 76300 18342
rect 76248 18278 76300 18284
rect 75512 17792 75564 17798
rect 75512 17734 75564 17740
rect 76156 17520 76208 17526
rect 76156 17462 76208 17468
rect 67784 17112 67836 17118
rect 67784 17054 67836 17060
rect 66864 12284 66916 12290
rect 66864 12226 66916 12232
rect 66876 9304 66904 12226
rect 76168 12154 76196 17462
rect 76260 12290 76288 18278
rect 77180 17594 77208 20846
rect 77548 20846 77884 20874
rect 78928 20846 78988 20874
rect 79664 20846 80000 20874
rect 80676 20846 81012 20874
rect 81688 20846 82024 20874
rect 83128 20846 83464 20874
rect 84140 20846 84384 20874
rect 85152 20846 85488 20874
rect 86164 20846 86500 20874
rect 87268 20846 87604 20874
rect 77168 17588 77220 17594
rect 77168 17530 77220 17536
rect 77548 17526 77576 20846
rect 78928 18342 78956 20846
rect 78916 18336 78968 18342
rect 78916 18278 78968 18284
rect 79664 18274 79692 20846
rect 80676 18478 80704 20846
rect 80664 18472 80716 18478
rect 80664 18414 80716 18420
rect 79652 18268 79704 18274
rect 79652 18210 79704 18216
rect 81688 18138 81716 20846
rect 81676 18132 81728 18138
rect 81676 18074 81728 18080
rect 78824 17588 78876 17594
rect 78824 17530 78876 17536
rect 77536 17520 77588 17526
rect 77536 17462 77588 17468
rect 76248 12284 76300 12290
rect 76248 12226 76300 12232
rect 72844 12148 72896 12154
rect 72844 12090 72896 12096
rect 76156 12148 76208 12154
rect 76156 12090 76208 12096
rect 72856 9304 72884 12090
rect 78836 9304 78864 17530
rect 83436 12290 83464 20846
rect 84356 12358 84384 20846
rect 84804 17180 84856 17186
rect 84804 17122 84856 17128
rect 84344 12352 84396 12358
rect 84344 12294 84396 12300
rect 83424 12284 83476 12290
rect 83424 12226 83476 12232
rect 84816 9304 84844 17122
rect 85460 12562 85488 20846
rect 86472 17798 86500 20846
rect 86460 17792 86512 17798
rect 86460 17734 86512 17740
rect 87576 17254 87604 20846
rect 87944 20846 88280 20874
rect 87564 17248 87616 17254
rect 87564 17190 87616 17196
rect 87944 17186 87972 20846
rect 93372 19838 93400 46226
rect 94740 46216 94792 46222
rect 94740 46158 94792 46164
rect 101178 46184 101234 46193
rect 93912 44720 93964 44726
rect 93912 44662 93964 44668
rect 93924 44289 93952 44662
rect 94004 44652 94056 44658
rect 94004 44594 94056 44600
rect 94016 44425 94044 44594
rect 94002 44416 94058 44425
rect 94002 44351 94058 44360
rect 93910 44280 93966 44289
rect 93910 44215 93966 44224
rect 93912 43292 93964 43298
rect 93912 43234 93964 43240
rect 93924 42929 93952 43234
rect 94004 43224 94056 43230
rect 94002 43192 94004 43201
rect 94056 43192 94058 43201
rect 94002 43127 94058 43136
rect 93910 42920 93966 42929
rect 93910 42855 93966 42864
rect 94004 42612 94056 42618
rect 94004 42554 94056 42560
rect 94016 42521 94044 42554
rect 94002 42512 94058 42521
rect 94002 42447 94058 42456
rect 94004 41864 94056 41870
rect 94004 41806 94056 41812
rect 94016 41705 94044 41806
rect 94002 41696 94058 41705
rect 94002 41631 94058 41640
rect 94004 40504 94056 40510
rect 94004 40446 94056 40452
rect 94016 40209 94044 40446
rect 94002 40200 94058 40209
rect 94002 40135 94058 40144
rect 94002 39112 94058 39121
rect 93912 39076 93964 39082
rect 94002 39047 94058 39056
rect 93912 39018 93964 39024
rect 93924 38713 93952 39018
rect 94016 39014 94044 39047
rect 94004 39008 94056 39014
rect 94004 38950 94056 38956
rect 93910 38704 93966 38713
rect 93910 38639 93966 38648
rect 94004 37648 94056 37654
rect 94002 37616 94004 37625
rect 94056 37616 94058 37625
rect 94002 37551 94058 37560
rect 94004 37104 94056 37110
rect 94002 37072 94004 37081
rect 94056 37072 94058 37081
rect 94002 37007 94058 37016
rect 94004 36356 94056 36362
rect 94004 36298 94056 36304
rect 94016 36129 94044 36298
rect 94002 36120 94058 36129
rect 94002 36055 94058 36064
rect 93452 35064 93504 35070
rect 93452 35006 93504 35012
rect 93464 34633 93492 35006
rect 94004 34996 94056 35002
rect 94004 34938 94056 34944
rect 94016 34905 94044 34938
rect 94002 34896 94058 34905
rect 94002 34831 94058 34840
rect 93450 34624 93506 34633
rect 93450 34559 93506 34568
rect 93910 33672 93966 33681
rect 93820 33636 93872 33642
rect 93910 33607 93966 33616
rect 93820 33578 93872 33584
rect 93832 33001 93860 33578
rect 93924 33506 93952 33607
rect 94004 33568 94056 33574
rect 94004 33510 94056 33516
rect 93912 33500 93964 33506
rect 93912 33442 93964 33448
rect 94016 33409 94044 33510
rect 94002 33400 94058 33409
rect 94002 33335 94058 33344
rect 93818 32992 93874 33001
rect 93818 32927 93874 32936
rect 93912 32276 93964 32282
rect 93912 32218 93964 32224
rect 93924 31777 93952 32218
rect 94004 32208 94056 32214
rect 94004 32150 94056 32156
rect 94016 31913 94044 32150
rect 94002 31904 94058 31913
rect 94002 31839 94058 31848
rect 93910 31768 93966 31777
rect 93910 31703 93966 31712
rect 94004 30848 94056 30854
rect 94004 30790 94056 30796
rect 94016 30689 94044 30790
rect 94002 30680 94058 30689
rect 94002 30615 94058 30624
rect 93912 29488 93964 29494
rect 93912 29430 93964 29436
rect 94002 29456 94058 29465
rect 93924 29193 93952 29430
rect 94002 29391 94058 29400
rect 94016 29358 94044 29391
rect 94004 29352 94056 29358
rect 94004 29294 94056 29300
rect 93910 29184 93966 29193
rect 93910 29119 93966 29128
rect 93912 28196 93964 28202
rect 93912 28138 93964 28144
rect 93924 26745 93952 28138
rect 94004 28128 94056 28134
rect 94004 28070 94056 28076
rect 94016 27969 94044 28070
rect 94002 27960 94058 27969
rect 94002 27895 94058 27904
rect 93910 26736 93966 26745
rect 93910 26671 93966 26680
rect 94004 26360 94056 26366
rect 94002 26328 94004 26337
rect 94056 26328 94058 26337
rect 94002 26263 94058 26272
rect 93820 25408 93872 25414
rect 93820 25350 93872 25356
rect 93832 24569 93860 25350
rect 93912 25340 93964 25346
rect 93912 25282 93964 25288
rect 93924 24977 93952 25282
rect 94004 25272 94056 25278
rect 94002 25240 94004 25249
rect 94056 25240 94058 25249
rect 94002 25175 94058 25184
rect 93910 24968 93966 24977
rect 93910 24903 93966 24912
rect 93818 24560 93874 24569
rect 93818 24495 93874 24504
rect 94004 23912 94056 23918
rect 94004 23854 94056 23860
rect 94016 23753 94044 23854
rect 94002 23744 94058 23753
rect 94002 23679 94058 23688
rect 94004 22620 94056 22626
rect 94004 22562 94056 22568
rect 93912 22552 93964 22558
rect 94016 22529 94044 22562
rect 93912 22494 93964 22500
rect 94002 22520 94058 22529
rect 93924 22121 93952 22494
rect 94002 22455 94058 22464
rect 93910 22112 93966 22121
rect 93910 22047 93966 22056
rect 94004 21260 94056 21266
rect 94004 21202 94056 21208
rect 94016 21169 94044 21202
rect 94002 21160 94058 21169
rect 94002 21095 94058 21104
rect 93360 19832 93412 19838
rect 93360 19774 93412 19780
rect 94752 19770 94780 46158
rect 96120 46148 96172 46154
rect 101178 46119 101234 46128
rect 96120 46090 96172 46096
rect 96132 22354 96160 46090
rect 100994 45504 101050 45513
rect 100994 45439 101050 45448
rect 101008 44726 101036 45439
rect 101086 44824 101142 44833
rect 101086 44759 101142 44768
rect 100996 44720 101048 44726
rect 100996 44662 101048 44668
rect 100994 43736 101050 43745
rect 100994 43671 101050 43680
rect 100810 43464 100866 43473
rect 100810 43399 100866 43408
rect 96856 43360 96908 43366
rect 96856 43302 96908 43308
rect 96868 42618 96896 43302
rect 96856 42612 96908 42618
rect 96856 42554 96908 42560
rect 100824 41870 100852 43399
rect 101008 43366 101036 43671
rect 100996 43360 101048 43366
rect 100996 43302 101048 43308
rect 101100 43298 101128 44759
rect 101192 44658 101220 46119
rect 134298 45096 134354 45105
rect 134298 45031 134354 45040
rect 101270 44960 101326 44969
rect 101270 44895 101326 44904
rect 101180 44652 101232 44658
rect 101180 44594 101232 44600
rect 101088 43292 101140 43298
rect 101088 43234 101140 43240
rect 101284 43230 101312 44895
rect 134312 44862 134340 45031
rect 134300 44856 134352 44862
rect 134300 44798 134352 44804
rect 101272 43224 101324 43230
rect 101272 43166 101324 43172
rect 100994 42512 101050 42521
rect 100994 42447 101050 42456
rect 100902 42104 100958 42113
rect 100902 42039 100958 42048
rect 100812 41864 100864 41870
rect 100812 41806 100864 41812
rect 100810 40608 100866 40617
rect 100810 40543 100866 40552
rect 100824 39014 100852 40543
rect 100916 40510 100944 42039
rect 101008 41938 101036 42447
rect 100996 41932 101048 41938
rect 100996 41874 101048 41880
rect 100994 41288 101050 41297
rect 100994 41223 101050 41232
rect 101008 40578 101036 41223
rect 134588 40714 134616 46498
rect 134760 46488 134812 46494
rect 134758 46456 134760 46465
rect 134812 46456 134814 46465
rect 134758 46391 134814 46400
rect 135220 46420 135272 46426
rect 135220 46362 135272 46368
rect 135036 46352 135088 46358
rect 135036 46294 135088 46300
rect 134944 46284 134996 46290
rect 134944 46226 134996 46232
rect 134850 45504 134906 45513
rect 134850 45439 134906 45448
rect 134760 44924 134812 44930
rect 134760 44866 134812 44872
rect 134772 44833 134800 44866
rect 134758 44824 134814 44833
rect 134864 44794 134892 45439
rect 134758 44759 134814 44768
rect 134852 44788 134904 44794
rect 134852 44730 134904 44736
rect 134758 43872 134814 43881
rect 134758 43807 134814 43816
rect 134772 43706 134800 43807
rect 134760 43700 134812 43706
rect 134760 43642 134812 43648
rect 134758 43464 134814 43473
rect 134956 43450 134984 46226
rect 134758 43399 134814 43408
rect 134864 43422 134984 43450
rect 134772 43366 134800 43399
rect 134760 43360 134812 43366
rect 134760 43302 134812 43308
rect 134758 42648 134814 42657
rect 134758 42583 134814 42592
rect 134772 42346 134800 42583
rect 134760 42340 134812 42346
rect 134760 42282 134812 42288
rect 134758 42104 134814 42113
rect 134758 42039 134814 42048
rect 134772 42006 134800 42039
rect 134760 42000 134812 42006
rect 134760 41942 134812 41948
rect 134666 41288 134722 41297
rect 134666 41223 134722 41232
rect 134576 40708 134628 40714
rect 134576 40650 134628 40656
rect 134680 40646 134708 41223
rect 134758 41016 134814 41025
rect 134758 40951 134814 40960
rect 134772 40850 134800 40951
rect 134760 40844 134812 40850
rect 134760 40786 134812 40792
rect 134760 40708 134812 40714
rect 134760 40650 134812 40656
rect 134668 40640 134720 40646
rect 134668 40582 134720 40588
rect 100996 40572 101048 40578
rect 100996 40514 101048 40520
rect 100904 40504 100956 40510
rect 100904 40446 100956 40452
rect 101086 40064 101142 40073
rect 101086 39999 101142 40008
rect 134574 40064 134630 40073
rect 134574 39999 134630 40008
rect 100994 39384 101050 39393
rect 100994 39319 101050 39328
rect 101008 39150 101036 39319
rect 100996 39144 101048 39150
rect 100996 39086 101048 39092
rect 101100 39082 101128 39999
rect 134588 39286 134616 39999
rect 134666 39520 134722 39529
rect 134666 39455 134722 39464
rect 134576 39280 134628 39286
rect 134576 39222 134628 39228
rect 134680 39218 134708 39455
rect 134668 39212 134720 39218
rect 134668 39154 134720 39160
rect 101088 39076 101140 39082
rect 101088 39018 101140 39024
rect 100812 39008 100864 39014
rect 100812 38950 100864 38956
rect 101086 38840 101142 38849
rect 101086 38775 101142 38784
rect 134114 38840 134170 38849
rect 134114 38775 134170 38784
rect 100994 38296 101050 38305
rect 100994 38231 101050 38240
rect 98236 37920 98288 37926
rect 98236 37862 98288 37868
rect 100810 37888 100866 37897
rect 98248 37654 98276 37862
rect 98328 37852 98380 37858
rect 101008 37858 101036 38231
rect 101100 37926 101128 38775
rect 101088 37920 101140 37926
rect 101088 37862 101140 37868
rect 134128 37858 134156 38775
rect 134298 38296 134354 38305
rect 134298 38231 134354 38240
rect 134312 37926 134340 38231
rect 134666 38024 134722 38033
rect 134666 37959 134668 37968
rect 134720 37959 134722 37968
rect 134668 37930 134720 37936
rect 134300 37920 134352 37926
rect 134300 37862 134352 37868
rect 100810 37823 100866 37832
rect 100996 37852 101048 37858
rect 98328 37794 98380 37800
rect 98236 37648 98288 37654
rect 98236 37590 98288 37596
rect 98340 37110 98368 37794
rect 98328 37104 98380 37110
rect 98328 37046 98380 37052
rect 100824 36362 100852 37823
rect 100996 37794 101048 37800
rect 134116 37852 134168 37858
rect 134116 37794 134168 37800
rect 100994 36936 101050 36945
rect 100994 36871 101050 36880
rect 134666 36936 134722 36945
rect 134666 36871 134722 36880
rect 100902 36528 100958 36537
rect 100902 36463 100958 36472
rect 100812 36356 100864 36362
rect 100812 36298 100864 36304
rect 100718 35168 100774 35177
rect 100718 35103 100774 35112
rect 100732 33506 100760 35103
rect 100916 35002 100944 36463
rect 101008 36430 101036 36871
rect 134390 36664 134446 36673
rect 134390 36599 134392 36608
rect 134444 36599 134446 36608
rect 134392 36570 134444 36576
rect 134680 36498 134708 36871
rect 134668 36492 134720 36498
rect 134668 36434 134720 36440
rect 100996 36424 101048 36430
rect 100996 36366 101048 36372
rect 134666 35984 134722 35993
rect 134666 35919 134722 35928
rect 100994 35712 101050 35721
rect 134680 35682 134708 35919
rect 100994 35647 101050 35656
rect 134668 35676 134720 35682
rect 101008 35070 101036 35647
rect 134668 35618 134720 35624
rect 134114 35304 134170 35313
rect 134114 35239 134170 35248
rect 134128 35138 134156 35239
rect 134116 35132 134168 35138
rect 134116 35074 134168 35080
rect 100996 35064 101048 35070
rect 100996 35006 101048 35012
rect 100904 34996 100956 35002
rect 100904 34938 100956 34944
rect 101086 34488 101142 34497
rect 101086 34423 101142 34432
rect 134574 34488 134630 34497
rect 134574 34423 134630 34432
rect 100994 33944 101050 33953
rect 100994 33879 101050 33888
rect 100810 33808 100866 33817
rect 100810 33743 100866 33752
rect 100720 33500 100772 33506
rect 100720 33442 100772 33448
rect 100824 32214 100852 33743
rect 101008 33642 101036 33879
rect 100996 33636 101048 33642
rect 100996 33578 101048 33584
rect 101100 33574 101128 34423
rect 134588 33710 134616 34423
rect 134666 34216 134722 34225
rect 134666 34151 134722 34160
rect 134680 34050 134708 34151
rect 134668 34044 134720 34050
rect 134668 33986 134720 33992
rect 134666 33808 134722 33817
rect 134666 33743 134668 33752
rect 134720 33743 134722 33752
rect 134668 33714 134720 33720
rect 134576 33704 134628 33710
rect 134576 33646 134628 33652
rect 101088 33568 101140 33574
rect 101088 33510 101140 33516
rect 100994 32720 101050 32729
rect 100994 32655 101050 32664
rect 134298 32720 134354 32729
rect 134298 32655 134354 32664
rect 100902 32312 100958 32321
rect 101008 32282 101036 32655
rect 134312 32350 134340 32655
rect 134390 32448 134446 32457
rect 134390 32383 134392 32392
rect 134444 32383 134446 32392
rect 134392 32354 134444 32360
rect 134300 32344 134352 32350
rect 134300 32286 134352 32292
rect 100902 32247 100958 32256
rect 100996 32276 101048 32282
rect 100812 32208 100864 32214
rect 100812 32150 100864 32156
rect 100810 30952 100866 30961
rect 100810 30887 100866 30896
rect 100824 29358 100852 30887
rect 100916 30854 100944 32247
rect 100996 32218 101048 32224
rect 134666 31632 134722 31641
rect 134666 31567 134722 31576
rect 100994 31496 101050 31505
rect 100994 31431 101050 31440
rect 101008 30922 101036 31431
rect 134680 31330 134708 31567
rect 134668 31324 134720 31330
rect 134668 31266 134720 31272
rect 134666 31088 134722 31097
rect 134666 31023 134722 31032
rect 134680 30990 134708 31023
rect 134668 30984 134720 30990
rect 134668 30926 134720 30932
rect 100996 30916 101048 30922
rect 100996 30858 101048 30864
rect 134392 30916 134444 30922
rect 134392 30858 134444 30864
rect 100904 30848 100956 30854
rect 100904 30790 100956 30796
rect 101086 30272 101142 30281
rect 101086 30207 101142 30216
rect 100994 29728 101050 29737
rect 100994 29663 101050 29672
rect 101008 29426 101036 29663
rect 101100 29494 101128 30207
rect 134206 29864 134262 29873
rect 134206 29799 134262 29808
rect 134220 29562 134248 29799
rect 134208 29556 134260 29562
rect 134208 29498 134260 29504
rect 101088 29488 101140 29494
rect 101088 29430 101140 29436
rect 100996 29420 101048 29426
rect 100996 29362 101048 29368
rect 100812 29352 100864 29358
rect 100812 29294 100864 29300
rect 101178 29048 101234 29057
rect 101178 28983 101234 28992
rect 101086 28504 101142 28513
rect 101086 28439 101142 28448
rect 100994 28232 101050 28241
rect 100994 28167 100996 28176
rect 101048 28167 101050 28176
rect 100996 28138 101048 28144
rect 101100 28066 101128 28439
rect 101192 28134 101220 28983
rect 101180 28128 101232 28134
rect 101180 28070 101232 28076
rect 101088 28060 101140 28066
rect 101088 28002 101140 28008
rect 100994 27280 101050 27289
rect 100994 27215 101050 27224
rect 101008 26842 101036 27215
rect 101178 26872 101234 26881
rect 98236 26836 98288 26842
rect 98236 26778 98288 26784
rect 100996 26836 101048 26842
rect 101178 26807 101234 26816
rect 100996 26778 101048 26784
rect 98248 26366 98276 26778
rect 98236 26360 98288 26366
rect 98236 26302 98288 26308
rect 101086 26056 101142 26065
rect 101086 25991 101142 26000
rect 100994 25648 101050 25657
rect 100994 25583 101050 25592
rect 101008 25414 101036 25583
rect 100996 25408 101048 25414
rect 100996 25350 101048 25356
rect 101100 25346 101128 25991
rect 101088 25340 101140 25346
rect 101088 25282 101140 25288
rect 101192 25278 101220 26807
rect 101180 25272 101232 25278
rect 101180 25214 101232 25220
rect 101086 24832 101142 24841
rect 101086 24767 101142 24776
rect 100994 24152 101050 24161
rect 100994 24087 101050 24096
rect 101008 23986 101036 24087
rect 100996 23980 101048 23986
rect 100996 23922 101048 23928
rect 101100 23918 101128 24767
rect 101088 23912 101140 23918
rect 101088 23854 101140 23860
rect 100994 23608 101050 23617
rect 100994 23543 101050 23552
rect 101008 22762 101036 23543
rect 101086 22928 101142 22937
rect 101086 22863 101142 22872
rect 100996 22756 101048 22762
rect 100996 22698 101048 22704
rect 101100 22694 101128 22863
rect 101088 22688 101140 22694
rect 101088 22630 101140 22636
rect 101178 22656 101234 22665
rect 100996 22620 101048 22626
rect 134404 22626 134432 30858
rect 134772 30394 134800 40650
rect 134864 30922 134892 43422
rect 134944 43292 134996 43298
rect 134944 43234 134996 43240
rect 134852 30916 134904 30922
rect 134852 30858 134904 30864
rect 134496 30366 134800 30394
rect 101178 22591 101234 22600
rect 134392 22620 134444 22626
rect 100996 22562 101048 22568
rect 101008 22393 101036 22562
rect 101088 22552 101140 22558
rect 101088 22494 101140 22500
rect 100994 22384 101050 22393
rect 96120 22348 96172 22354
rect 100994 22319 101050 22328
rect 96120 22290 96172 22296
rect 101100 21985 101128 22494
rect 101086 21976 101142 21985
rect 101086 21911 101142 21920
rect 101192 21266 101220 22591
rect 134392 22562 134444 22568
rect 101180 21260 101232 21266
rect 101180 21202 101232 21208
rect 101824 19832 101876 19838
rect 101546 19800 101602 19809
rect 94740 19764 94792 19770
rect 101824 19774 101876 19780
rect 101546 19735 101548 19744
rect 94740 19706 94792 19712
rect 101600 19735 101602 19744
rect 101548 19706 101600 19712
rect 101836 19537 101864 19774
rect 134496 19537 134524 30366
rect 134758 30272 134814 30281
rect 134758 30207 134814 30216
rect 134772 29630 134800 30207
rect 134760 29624 134812 29630
rect 134760 29566 134812 29572
rect 134574 29048 134630 29057
rect 134574 28983 134630 28992
rect 134588 28202 134616 28983
rect 134758 28640 134814 28649
rect 134758 28575 134814 28584
rect 134772 28474 134800 28575
rect 134760 28468 134812 28474
rect 134760 28410 134812 28416
rect 134760 28264 134812 28270
rect 134758 28232 134760 28241
rect 134812 28232 134814 28241
rect 134576 28196 134628 28202
rect 134758 28167 134814 28176
rect 134576 28138 134628 28144
rect 134574 27280 134630 27289
rect 134574 27215 134630 27224
rect 134588 26842 134616 27215
rect 134758 27008 134814 27017
rect 134758 26943 134814 26952
rect 134772 26910 134800 26943
rect 134760 26904 134812 26910
rect 134760 26846 134812 26852
rect 134576 26836 134628 26842
rect 134576 26778 134628 26784
rect 134574 26056 134630 26065
rect 134574 25991 134630 26000
rect 134588 25482 134616 25991
rect 134758 25648 134814 25657
rect 134758 25583 134814 25592
rect 134772 25550 134800 25583
rect 134760 25544 134812 25550
rect 134760 25486 134812 25492
rect 134576 25476 134628 25482
rect 134576 25418 134628 25424
rect 134574 24832 134630 24841
rect 134574 24767 134630 24776
rect 134588 24122 134616 24767
rect 134758 24288 134814 24297
rect 134758 24223 134814 24232
rect 134576 24116 134628 24122
rect 134576 24058 134628 24064
rect 134772 24054 134800 24223
rect 134760 24048 134812 24054
rect 134760 23990 134812 23996
rect 134574 23608 134630 23617
rect 134574 23543 134630 23552
rect 134588 22694 134616 23543
rect 134758 23200 134814 23209
rect 134758 23135 134814 23144
rect 134772 23034 134800 23135
rect 134760 23028 134812 23034
rect 134760 22970 134812 22976
rect 134758 22792 134814 22801
rect 134758 22727 134760 22736
rect 134812 22727 134814 22736
rect 134760 22698 134812 22704
rect 134576 22688 134628 22694
rect 134576 22630 134628 22636
rect 134760 22620 134812 22626
rect 134760 22562 134812 22568
rect 134772 21169 134800 22562
rect 134758 21160 134814 21169
rect 134758 21095 134814 21104
rect 134956 19809 134984 43234
rect 135048 20761 135076 46294
rect 135128 46216 135180 46222
rect 135128 46158 135180 46164
rect 135140 21985 135168 46158
rect 135232 43298 135260 46362
rect 138360 46193 138388 55678
rect 145340 46556 145392 46562
rect 145340 46498 145392 46504
rect 142580 46488 142632 46494
rect 142580 46430 142632 46436
rect 138346 46184 138402 46193
rect 135312 46148 135364 46154
rect 135312 46090 135364 46096
rect 138070 46150 138126 46159
rect 138346 46119 138402 46128
rect 135220 43292 135272 43298
rect 135220 43234 135272 43240
rect 135324 22529 135352 46090
rect 138070 46085 138126 46094
rect 138084 40714 138112 46085
rect 142488 44856 142540 44862
rect 142488 44798 142540 44804
rect 142396 44720 142448 44726
rect 142396 44662 142448 44668
rect 142408 44289 142436 44662
rect 142394 44280 142450 44289
rect 142394 44215 142450 44224
rect 139636 43700 139688 43706
rect 139636 43642 139688 43648
rect 139648 43298 139676 43642
rect 139636 43292 139688 43298
rect 139636 43234 139688 43240
rect 142500 43201 142528 44798
rect 142592 44425 142620 46430
rect 142672 44924 142724 44930
rect 142672 44866 142724 44872
rect 142578 44416 142634 44425
rect 142578 44351 142634 44360
rect 142486 43192 142542 43201
rect 142486 43127 142542 43136
rect 142684 43065 142712 44866
rect 145352 44810 145380 46498
rect 146812 46420 146864 46426
rect 146812 46362 146864 46368
rect 146824 44810 146852 46362
rect 148284 46352 148336 46358
rect 148284 46294 148336 46300
rect 148296 44810 148324 46294
rect 149756 46284 149808 46290
rect 149756 46226 149808 46232
rect 149768 44810 149796 46226
rect 151320 46216 151372 46222
rect 151320 46158 151372 46164
rect 154262 46184 154318 46193
rect 151332 44810 151360 46158
rect 152792 46148 152844 46154
rect 154262 46119 154318 46128
rect 152792 46090 152844 46096
rect 152804 44810 152832 46090
rect 154276 44810 154304 46119
rect 156116 44810 156144 57786
rect 183072 49622 183100 68831
rect 183808 68186 183836 72526
rect 188500 69546 188528 73698
rect 190800 70809 190828 73698
rect 191984 73688 192036 73694
rect 191984 73630 192036 73636
rect 191996 72849 192024 73630
rect 191982 72840 192038 72849
rect 191982 72775 192038 72784
rect 191524 70968 191576 70974
rect 191524 70910 191576 70916
rect 190786 70800 190842 70809
rect 190786 70735 190842 70744
rect 189960 69948 190012 69954
rect 189960 69890 190012 69896
rect 188488 69540 188540 69546
rect 188488 69482 188540 69488
rect 183796 68180 183848 68186
rect 183796 68122 183848 68128
rect 183150 67672 183206 67681
rect 183150 67607 183206 67616
rect 183060 49616 183112 49622
rect 183060 49558 183112 49564
rect 183164 49554 183192 67607
rect 183242 66448 183298 66457
rect 183242 66383 183298 66392
rect 183256 49690 183284 66383
rect 183334 65224 183390 65233
rect 183334 65159 183390 65168
rect 183244 49684 183296 49690
rect 183244 49626 183296 49632
rect 183152 49548 183204 49554
rect 183152 49490 183204 49496
rect 183348 49146 183376 65159
rect 183610 64000 183666 64009
rect 183610 63935 183666 63944
rect 183426 62776 183482 62785
rect 183426 62711 183482 62720
rect 183440 49350 183468 62711
rect 183428 49344 183480 49350
rect 183428 49286 183480 49292
rect 183624 49282 183652 63935
rect 189972 62785 190000 69890
rect 190972 69540 191024 69546
rect 190972 69482 191024 69488
rect 190984 68769 191012 69482
rect 190970 68760 191026 68769
rect 190970 68695 191026 68704
rect 191340 68180 191392 68186
rect 191340 68122 191392 68128
rect 191352 66865 191380 68122
rect 191338 66856 191394 66865
rect 191338 66791 191394 66800
rect 191536 64825 191564 70910
rect 191522 64816 191578 64825
rect 191522 64751 191578 64760
rect 189958 62776 190014 62785
rect 189958 62711 190014 62720
rect 183702 61552 183758 61561
rect 183702 61487 183704 61496
rect 183756 61487 183758 61496
rect 188028 61516 188080 61522
rect 183704 61458 183756 61464
rect 188028 61458 188080 61464
rect 184440 60428 184492 60434
rect 184440 60370 184492 60376
rect 184452 50234 184480 60370
rect 188040 50522 188068 61458
rect 191982 60872 192038 60881
rect 191982 60807 192038 60816
rect 188040 50494 188344 50522
rect 184440 50228 184492 50234
rect 184440 50170 184492 50176
rect 188212 50228 188264 50234
rect 188212 50170 188264 50176
rect 183612 49276 183664 49282
rect 183612 49218 183664 49224
rect 183336 49140 183388 49146
rect 183336 49082 183388 49088
rect 164750 46864 164806 46873
rect 164750 46799 164806 46808
rect 161898 46728 161954 46737
rect 161898 46663 161954 46672
rect 158954 46592 159010 46601
rect 158954 46527 159010 46536
rect 157574 46320 157630 46329
rect 157574 46255 157630 46264
rect 157588 44810 157616 46255
rect 158968 44810 158996 46527
rect 160334 46456 160390 46465
rect 160334 46391 160390 46400
rect 160348 44810 160376 46391
rect 161912 44810 161940 46663
rect 163278 46320 163334 46329
rect 163278 46255 163334 46264
rect 163292 44810 163320 46255
rect 164764 44810 164792 46799
rect 188224 46700 188252 50170
rect 188316 46714 188344 50494
rect 191064 49684 191116 49690
rect 191064 49626 191116 49632
rect 189316 49344 189368 49350
rect 189316 49286 189368 49292
rect 188316 46686 188790 46714
rect 189328 46700 189356 49286
rect 189868 49276 189920 49282
rect 189868 49218 189920 49224
rect 189880 46700 189908 49218
rect 190420 49140 190472 49146
rect 190420 49082 190472 49088
rect 190432 46700 190460 49082
rect 191076 46700 191104 49626
rect 191996 49554 192024 60807
rect 193364 57232 193416 57238
rect 193364 57174 193416 57180
rect 193272 57164 193324 57170
rect 193272 57106 193324 57112
rect 192168 49616 192220 49622
rect 192168 49558 192220 49564
rect 191616 49548 191668 49554
rect 191616 49490 191668 49496
rect 191984 49548 192036 49554
rect 191984 49490 192036 49496
rect 191628 46700 191656 49490
rect 192180 46700 192208 49558
rect 193284 47122 193312 57106
rect 193192 47094 193312 47122
rect 193192 46714 193220 47094
rect 193376 46714 193404 57174
rect 194112 57170 194140 59892
rect 194480 57238 194508 59892
rect 194652 57300 194704 57306
rect 194652 57242 194704 57248
rect 194468 57232 194520 57238
rect 194468 57174 194520 57180
rect 194100 57164 194152 57170
rect 194100 57106 194152 57112
rect 194192 54376 194244 54382
rect 194192 54318 194244 54324
rect 194204 46714 194232 54318
rect 194664 46714 194692 57242
rect 194848 57186 194876 59892
rect 195308 57306 195336 59892
rect 195296 57300 195348 57306
rect 195296 57242 195348 57248
rect 194756 57158 194876 57186
rect 195112 57232 195164 57238
rect 195112 57174 195164 57180
rect 194928 57164 194980 57170
rect 194756 54382 194784 57158
rect 194928 57106 194980 57112
rect 194744 54376 194796 54382
rect 194744 54318 194796 54324
rect 192746 46686 193220 46714
rect 193298 46686 193404 46714
rect 193942 46686 194232 46714
rect 194494 46686 194692 46714
rect 194940 46714 194968 57106
rect 195124 46714 195152 57174
rect 195676 57170 195704 59892
rect 196044 57238 196072 59892
rect 196228 59878 196518 59906
rect 196032 57232 196084 57238
rect 196228 57186 196256 59878
rect 196872 57238 196900 59892
rect 196032 57174 196084 57180
rect 195664 57164 195716 57170
rect 195664 57106 195716 57112
rect 196136 57158 196256 57186
rect 196400 57232 196452 57238
rect 196400 57174 196452 57180
rect 196860 57232 196912 57238
rect 196860 57174 196912 57180
rect 196308 57164 196360 57170
rect 194940 46686 195046 46714
rect 195124 46686 195598 46714
rect 196136 46700 196164 57158
rect 196308 57106 196360 57112
rect 196320 57050 196348 57106
rect 196228 57022 196348 57050
rect 196228 50438 196256 57022
rect 196412 56914 196440 57174
rect 197240 57170 197268 59892
rect 197608 59878 197714 59906
rect 197792 59878 198082 59906
rect 198450 59878 198832 59906
rect 197228 57164 197280 57170
rect 197228 57106 197280 57112
rect 196320 56886 196440 56914
rect 196216 50432 196268 50438
rect 196216 50374 196268 50380
rect 196320 46850 196348 56886
rect 197044 50432 197096 50438
rect 197044 50374 197096 50380
rect 196320 46822 196624 46850
rect 196596 46714 196624 46822
rect 197056 46714 197084 50374
rect 197608 46714 197636 59878
rect 197792 57186 197820 59878
rect 197700 57158 197820 57186
rect 198804 57186 198832 59878
rect 198896 57306 198924 59892
rect 199080 59878 199278 59906
rect 198884 57300 198936 57306
rect 198884 57242 198936 57248
rect 198804 57158 199016 57186
rect 197700 50438 197728 57158
rect 198988 54382 199016 57158
rect 198976 54376 199028 54382
rect 198976 54318 199028 54324
rect 199080 50438 199108 59878
rect 199632 58530 199660 59892
rect 200106 59878 200304 59906
rect 200474 59878 200764 59906
rect 200276 58682 200304 59878
rect 200276 58654 200488 58682
rect 199620 58524 199672 58530
rect 199620 58466 199672 58472
rect 200356 58524 200408 58530
rect 200356 58466 200408 58472
rect 199160 57300 199212 57306
rect 199160 57242 199212 57248
rect 197688 50432 197740 50438
rect 197688 50374 197740 50380
rect 198148 50432 198200 50438
rect 198148 50374 198200 50380
rect 199068 50432 199120 50438
rect 199068 50374 199120 50380
rect 198160 46714 198188 50374
rect 199068 50296 199120 50302
rect 199068 50238 199120 50244
rect 199080 46714 199108 50238
rect 196596 46686 196794 46714
rect 197056 46686 197346 46714
rect 197608 46686 197898 46714
rect 198160 46686 198450 46714
rect 199002 46686 199108 46714
rect 199172 46714 199200 57242
rect 199252 54376 199304 54382
rect 199252 54318 199304 54324
rect 199264 50302 199292 54318
rect 199804 50432 199856 50438
rect 199804 50374 199856 50380
rect 199252 50296 199304 50302
rect 199252 50238 199304 50244
rect 199816 46714 199844 50374
rect 200368 46714 200396 58466
rect 200460 46986 200488 58654
rect 200736 57374 200764 59878
rect 200724 57368 200776 57374
rect 200724 57310 200776 57316
rect 200828 57170 200856 59892
rect 201288 57306 201316 59892
rect 201276 57300 201328 57306
rect 201276 57242 201328 57248
rect 201656 57238 201684 59892
rect 201828 57368 201880 57374
rect 201828 57310 201880 57316
rect 201644 57232 201696 57238
rect 201644 57174 201696 57180
rect 200816 57164 200868 57170
rect 200816 57106 200868 57112
rect 200460 46958 201040 46986
rect 201012 46714 201040 46958
rect 199172 46686 199646 46714
rect 199816 46686 200198 46714
rect 200368 46686 200750 46714
rect 201012 46686 201302 46714
rect 201840 46700 201868 57310
rect 202116 57170 202144 59892
rect 202484 57374 202512 59892
rect 202472 57368 202524 57374
rect 202472 57310 202524 57316
rect 202196 57300 202248 57306
rect 202196 57242 202248 57248
rect 201920 57164 201972 57170
rect 201920 57106 201972 57112
rect 202104 57164 202156 57170
rect 202104 57106 202156 57112
rect 201932 46850 201960 57106
rect 202208 46952 202236 57242
rect 202852 57238 202880 59892
rect 203312 57442 203340 59892
rect 203300 57436 203352 57442
rect 203300 57378 203352 57384
rect 203680 57306 203708 59892
rect 203668 57300 203720 57306
rect 203668 57242 203720 57248
rect 202380 57232 202432 57238
rect 202380 57174 202432 57180
rect 202840 57232 202892 57238
rect 202840 57174 202892 57180
rect 202392 50098 202420 57174
rect 204048 57170 204076 59892
rect 204508 57578 204536 59892
rect 204496 57572 204548 57578
rect 204496 57514 204548 57520
rect 204876 57374 204904 59892
rect 205244 57510 205272 59892
rect 205232 57504 205284 57510
rect 205232 57446 205284 57452
rect 205324 57436 205376 57442
rect 205324 57378 205376 57384
rect 204588 57368 204640 57374
rect 204588 57310 204640 57316
rect 204864 57368 204916 57374
rect 204864 57310 204916 57316
rect 204496 57232 204548 57238
rect 204496 57174 204548 57180
rect 203024 57164 203076 57170
rect 203024 57106 203076 57112
rect 204036 57164 204088 57170
rect 204036 57106 204088 57112
rect 202380 50092 202432 50098
rect 202380 50034 202432 50040
rect 203036 49146 203064 57106
rect 204508 50438 204536 57174
rect 204496 50432 204548 50438
rect 204496 50374 204548 50380
rect 203576 50092 203628 50098
rect 203576 50034 203628 50040
rect 203024 49140 203076 49146
rect 203024 49082 203076 49088
rect 202208 46924 202696 46952
rect 201932 46822 202328 46850
rect 202300 46714 202328 46822
rect 202668 46714 202696 46924
rect 202300 46686 202498 46714
rect 202668 46686 203050 46714
rect 203588 46700 203616 50034
rect 204128 49140 204180 49146
rect 204128 49082 204180 49088
rect 204140 46700 204168 49082
rect 204600 46714 204628 57310
rect 205232 57300 205284 57306
rect 205232 57242 205284 57248
rect 205140 57164 205192 57170
rect 205140 57106 205192 57112
rect 204956 50432 205008 50438
rect 204956 50374 205008 50380
rect 204968 46714 204996 50374
rect 205152 50098 205180 57106
rect 205244 50166 205272 57242
rect 205336 50234 205364 57378
rect 205704 57238 205732 59892
rect 205692 57232 205744 57238
rect 205692 57174 205744 57180
rect 206072 57170 206100 59892
rect 206440 57646 206468 59892
rect 206428 57640 206480 57646
rect 206428 57582 206480 57588
rect 206900 57442 206928 59892
rect 207268 58258 207296 59892
rect 207636 58394 207664 59892
rect 208096 58530 208124 59892
rect 208084 58524 208136 58530
rect 208084 58466 208136 58472
rect 207624 58388 207676 58394
rect 207624 58330 207676 58336
rect 207256 58252 207308 58258
rect 207256 58194 207308 58200
rect 208464 57850 208492 59892
rect 208832 58326 208860 59892
rect 208820 58320 208872 58326
rect 208820 58262 208872 58268
rect 209292 58122 209320 59892
rect 209660 58462 209688 59892
rect 210660 58524 210712 58530
rect 210660 58466 210712 58472
rect 209648 58456 209700 58462
rect 209648 58398 209700 58404
rect 209280 58116 209332 58122
rect 209280 58058 209332 58064
rect 208452 57844 208504 57850
rect 208452 57786 208504 57792
rect 210108 57640 210160 57646
rect 210108 57582 210160 57588
rect 207256 57572 207308 57578
rect 207256 57514 207308 57520
rect 206888 57436 206940 57442
rect 206888 57378 206940 57384
rect 206060 57164 206112 57170
rect 206060 57106 206112 57112
rect 207164 57164 207216 57170
rect 207164 57106 207216 57112
rect 205324 50228 205376 50234
rect 205324 50170 205376 50176
rect 205876 50228 205928 50234
rect 205876 50170 205928 50176
rect 205232 50160 205284 50166
rect 205232 50102 205284 50108
rect 205140 50092 205192 50098
rect 205140 50034 205192 50040
rect 204600 46686 204706 46714
rect 204968 46686 205350 46714
rect 205888 46700 205916 50170
rect 206428 50160 206480 50166
rect 206428 50102 206480 50108
rect 206440 46700 206468 50102
rect 206980 50092 207032 50098
rect 206980 50034 207032 50040
rect 206992 46700 207020 50034
rect 207176 49214 207204 57106
rect 207164 49208 207216 49214
rect 207164 49150 207216 49156
rect 207268 46714 207296 57514
rect 207992 57504 208044 57510
rect 207992 57446 208044 57452
rect 207348 57368 207400 57374
rect 207348 57310 207400 57316
rect 207360 46952 207388 57310
rect 207900 57232 207952 57238
rect 207900 57174 207952 57180
rect 207912 50166 207940 57174
rect 208004 50234 208032 57446
rect 210016 57436 210068 57442
rect 210016 57378 210068 57384
rect 210028 50438 210056 57378
rect 210016 50432 210068 50438
rect 210016 50374 210068 50380
rect 207992 50228 208044 50234
rect 207992 50170 208044 50176
rect 208728 50228 208780 50234
rect 208728 50170 208780 50176
rect 207900 50160 207952 50166
rect 207900 50102 207952 50108
rect 207360 46924 207664 46952
rect 207636 46714 207664 46924
rect 207268 46686 207558 46714
rect 207636 46686 208202 46714
rect 208740 46700 208768 50170
rect 209280 50160 209332 50166
rect 209280 50102 209332 50108
rect 209292 46700 209320 50102
rect 209832 49208 209884 49214
rect 209832 49150 209884 49156
rect 209844 46700 209872 49150
rect 210120 46714 210148 57582
rect 210672 50574 210700 58466
rect 210752 58388 210804 58394
rect 210752 58330 210804 58336
rect 210660 50568 210712 50574
rect 210660 50510 210712 50516
rect 210660 50432 210712 50438
rect 210660 50374 210712 50380
rect 210672 46714 210700 50374
rect 210764 50234 210792 58330
rect 210844 58252 210896 58258
rect 210844 58194 210896 58200
rect 210752 50228 210804 50234
rect 210752 50170 210804 50176
rect 210856 49554 210884 58194
rect 210936 50568 210988 50574
rect 210936 50510 210988 50516
rect 210948 50166 210976 50510
rect 210936 50160 210988 50166
rect 210936 50102 210988 50108
rect 210844 49548 210896 49554
rect 210844 49490 210896 49496
rect 211580 49548 211632 49554
rect 211580 49490 211632 49496
rect 210120 46686 210410 46714
rect 210672 46686 211054 46714
rect 211592 46700 211620 49490
rect 212052 48874 212080 83111
rect 212144 75054 212172 89775
rect 212132 75048 212184 75054
rect 212132 74990 212184 74996
rect 222344 75048 222396 75054
rect 222344 74990 222396 74996
rect 222356 74345 222384 74990
rect 222342 74336 222398 74345
rect 222342 74271 222398 74280
rect 212682 69848 212738 69857
rect 212682 69783 212684 69792
rect 212736 69783 212738 69792
rect 215628 69812 215680 69818
rect 212684 69754 212736 69760
rect 215628 69754 215680 69760
rect 212316 58456 212368 58462
rect 212316 58398 212368 58404
rect 212224 58320 212276 58326
rect 212224 58262 212276 58268
rect 212132 58116 212184 58122
rect 212132 58058 212184 58064
rect 212144 50370 212172 58058
rect 212132 50364 212184 50370
rect 212132 50306 212184 50312
rect 212132 50228 212184 50234
rect 212132 50170 212184 50176
rect 212040 48868 212092 48874
rect 212040 48810 212092 48816
rect 212144 46700 212172 50170
rect 212236 49690 212264 58262
rect 212224 49684 212276 49690
rect 212224 49626 212276 49632
rect 212328 49554 212356 58398
rect 212868 57844 212920 57850
rect 212868 57786 212920 57792
rect 212684 50160 212736 50166
rect 212684 50102 212736 50108
rect 212316 49548 212368 49554
rect 212316 49490 212368 49496
rect 212696 46700 212724 50102
rect 212880 46714 212908 57786
rect 214432 50228 214484 50234
rect 214432 50170 214484 50176
rect 213880 49684 213932 49690
rect 213880 49626 213932 49632
rect 212880 46686 213262 46714
rect 213892 46700 213920 49626
rect 214444 46700 214472 50170
rect 215536 49616 215588 49622
rect 215536 49558 215588 49564
rect 214984 49548 215036 49554
rect 214984 49490 215036 49496
rect 214996 46700 215024 49490
rect 215548 46700 215576 49558
rect 169902 46320 169958 46329
rect 169902 46255 169958 46264
rect 168432 46216 168484 46222
rect 168432 46158 168484 46164
rect 166960 46148 167012 46154
rect 166960 46090 167012 46096
rect 166972 44810 167000 46090
rect 168444 44810 168472 46158
rect 169916 44810 169944 46255
rect 177540 46216 177592 46222
rect 171098 46184 171154 46193
rect 177540 46158 177592 46164
rect 185818 46184 185874 46193
rect 171098 46119 171154 46128
rect 176160 46148 176212 46154
rect 145352 44782 145688 44810
rect 146824 44782 147160 44810
rect 148296 44782 148632 44810
rect 149768 44782 150104 44810
rect 151332 44782 151668 44810
rect 152804 44782 153140 44810
rect 154276 44782 154612 44810
rect 156116 44782 156176 44810
rect 157588 44782 157648 44810
rect 158968 44782 159120 44810
rect 160348 44782 160684 44810
rect 161912 44782 162156 44810
rect 163292 44782 163628 44810
rect 164764 44782 165100 44810
rect 166664 44782 167000 44810
rect 168136 44782 168472 44810
rect 169608 44782 169944 44810
rect 171112 44810 171140 46119
rect 176160 46090 176212 46096
rect 171112 44782 171172 44810
rect 172938 44688 172994 44697
rect 172644 44646 172938 44674
rect 172938 44623 172994 44632
rect 174116 44510 174452 44538
rect 143500 43360 143552 43366
rect 143500 43302 143552 43308
rect 143132 43292 143184 43298
rect 143132 43234 143184 43240
rect 142670 43056 142726 43065
rect 142670 42991 142726 43000
rect 143144 42521 143172 43234
rect 143130 42512 143186 42521
rect 143130 42447 143186 42456
rect 139636 42340 139688 42346
rect 139636 42282 139688 42288
rect 139648 41802 139676 42282
rect 143512 41977 143540 43302
rect 143684 42000 143736 42006
rect 143498 41968 143554 41977
rect 143684 41942 143736 41948
rect 143498 41903 143554 41912
rect 139636 41796 139688 41802
rect 139636 41738 139688 41744
rect 142764 41796 142816 41802
rect 142764 41738 142816 41744
rect 142776 41297 142804 41738
rect 142762 41288 142818 41297
rect 142762 41223 142818 41232
rect 139636 40844 139688 40850
rect 139636 40786 139688 40792
rect 138072 40708 138124 40714
rect 138072 40650 138124 40656
rect 137980 40572 138032 40578
rect 137980 40514 138032 40520
rect 135310 22520 135366 22529
rect 135310 22455 135366 22464
rect 135126 21976 135182 21985
rect 135126 21911 135182 21920
rect 137992 21266 138020 40514
rect 139648 39082 139676 40786
rect 142396 40572 142448 40578
rect 142396 40514 142448 40520
rect 142408 40073 142436 40514
rect 143696 40209 143724 41942
rect 143682 40200 143738 40209
rect 143682 40135 143738 40144
rect 142394 40064 142450 40073
rect 142394 39999 142450 40008
rect 142396 39144 142448 39150
rect 142396 39086 142448 39092
rect 142486 39112 142542 39121
rect 139636 39076 139688 39082
rect 139636 39018 139688 39024
rect 142408 38985 142436 39086
rect 142486 39047 142488 39056
rect 142540 39047 142542 39056
rect 142488 39018 142540 39024
rect 142580 39008 142632 39014
rect 142394 38976 142450 38985
rect 142580 38950 142632 38956
rect 142394 38911 142450 38920
rect 142592 38305 142620 38950
rect 142578 38296 142634 38305
rect 142578 38231 142634 38240
rect 142580 37988 142632 37994
rect 142580 37930 142632 37936
rect 142488 37920 142540 37926
rect 142488 37862 142540 37868
rect 142396 37852 142448 37858
rect 142396 37794 142448 37800
rect 142408 37761 142436 37794
rect 142394 37752 142450 37761
rect 142394 37687 142450 37696
rect 142500 37081 142528 37862
rect 142486 37072 142542 37081
rect 142486 37007 142542 37016
rect 140924 36628 140976 36634
rect 140924 36570 140976 36576
rect 140188 35676 140240 35682
rect 140188 35618 140240 35624
rect 140200 34934 140228 35618
rect 140936 35070 140964 36570
rect 142396 36492 142448 36498
rect 142396 36434 142448 36440
rect 142408 35993 142436 36434
rect 142592 36401 142620 37930
rect 142578 36392 142634 36401
rect 142578 36327 142634 36336
rect 142394 35984 142450 35993
rect 142394 35919 142450 35928
rect 142488 35132 142540 35138
rect 142488 35074 142540 35080
rect 140924 35064 140976 35070
rect 140924 35006 140976 35012
rect 140188 34928 140240 34934
rect 140188 34870 140240 34876
rect 142396 34928 142448 34934
rect 142396 34870 142448 34876
rect 142408 34769 142436 34870
rect 142394 34760 142450 34769
rect 142394 34695 142450 34704
rect 140188 34044 140240 34050
rect 140188 33986 140240 33992
rect 140200 33234 140228 33986
rect 140924 33772 140976 33778
rect 140924 33714 140976 33720
rect 140188 33228 140240 33234
rect 140188 33170 140240 33176
rect 139728 32412 139780 32418
rect 139728 32354 139780 32360
rect 139636 31324 139688 31330
rect 139636 31266 139688 31272
rect 139648 30582 139676 31266
rect 139740 30786 139768 32354
rect 140936 32214 140964 33714
rect 142500 33681 142528 35074
rect 142580 35064 142632 35070
rect 142580 35006 142632 35012
rect 142592 34905 142620 35006
rect 142578 34896 142634 34905
rect 142578 34831 142634 34840
rect 142486 33672 142542 33681
rect 142396 33636 142448 33642
rect 142486 33607 142542 33616
rect 142396 33578 142448 33584
rect 142408 33409 142436 33578
rect 142394 33400 142450 33409
rect 142394 33335 142450 33344
rect 142396 33228 142448 33234
rect 142396 33170 142448 33176
rect 142408 33001 142436 33170
rect 142394 32992 142450 33001
rect 142394 32927 142450 32936
rect 142396 32276 142448 32282
rect 142396 32218 142448 32224
rect 140924 32208 140976 32214
rect 140924 32150 140976 32156
rect 142408 31777 142436 32218
rect 142488 32208 142540 32214
rect 142486 32176 142488 32185
rect 142540 32176 142542 32185
rect 142486 32111 142542 32120
rect 142394 31768 142450 31777
rect 142394 31703 142450 31712
rect 143592 30984 143644 30990
rect 143592 30926 143644 30932
rect 139728 30780 139780 30786
rect 139728 30722 139780 30728
rect 142396 30780 142448 30786
rect 142396 30722 142448 30728
rect 142408 30689 142436 30722
rect 142394 30680 142450 30689
rect 142394 30615 142450 30624
rect 139636 30576 139688 30582
rect 142396 30576 142448 30582
rect 139636 30518 139688 30524
rect 142394 30544 142396 30553
rect 142448 30544 142450 30553
rect 142394 30479 142450 30488
rect 142396 29488 142448 29494
rect 143604 29465 143632 30926
rect 142396 29430 142448 29436
rect 143590 29456 143646 29465
rect 142408 29329 142436 29430
rect 142488 29420 142540 29426
rect 143590 29391 143646 29400
rect 142488 29362 142540 29368
rect 142394 29320 142450 29329
rect 142394 29255 142450 29264
rect 142500 28785 142528 29362
rect 142486 28776 142542 28785
rect 142486 28711 142542 28720
rect 140280 28468 140332 28474
rect 140280 28410 140332 28416
rect 140292 27794 140320 28410
rect 140924 28264 140976 28270
rect 140924 28206 140976 28212
rect 140280 27788 140332 27794
rect 140280 27730 140332 27736
rect 140936 26774 140964 28206
rect 142396 28128 142448 28134
rect 142396 28070 142448 28076
rect 142408 27969 142436 28070
rect 142394 27960 142450 27969
rect 142394 27895 142450 27904
rect 142396 27788 142448 27794
rect 142396 27730 142448 27736
rect 142408 27561 142436 27730
rect 142394 27552 142450 27561
rect 142394 27487 142450 27496
rect 142580 26904 142632 26910
rect 142580 26846 142632 26852
rect 142396 26836 142448 26842
rect 142396 26778 142448 26784
rect 140924 26768 140976 26774
rect 140924 26710 140976 26716
rect 142408 26337 142436 26778
rect 142488 26768 142540 26774
rect 142486 26736 142488 26745
rect 142540 26736 142542 26745
rect 142486 26671 142542 26680
rect 142394 26328 142450 26337
rect 142394 26263 142450 26272
rect 142488 25544 142540 25550
rect 142488 25486 142540 25492
rect 142396 25476 142448 25482
rect 142396 25418 142448 25424
rect 142408 25113 142436 25418
rect 142394 25104 142450 25113
rect 142394 25039 142450 25048
rect 142500 24569 142528 25486
rect 142592 25249 142620 26846
rect 142578 25240 142634 25249
rect 142578 25175 142634 25184
rect 142486 24560 142542 24569
rect 142486 24495 142542 24504
rect 142396 23980 142448 23986
rect 142396 23922 142448 23928
rect 142408 23889 142436 23922
rect 142488 23912 142540 23918
rect 142394 23880 142450 23889
rect 142488 23854 142540 23860
rect 142394 23815 142450 23824
rect 142500 23345 142528 23854
rect 142486 23336 142542 23345
rect 142486 23271 142542 23280
rect 140740 23028 140792 23034
rect 140740 22970 140792 22976
rect 139728 22756 139780 22762
rect 139728 22698 139780 22704
rect 139740 21266 139768 22698
rect 140752 22558 140780 22970
rect 142396 22620 142448 22626
rect 142396 22562 142448 22568
rect 140740 22552 140792 22558
rect 142408 22529 142436 22562
rect 142488 22552 142540 22558
rect 140740 22494 140792 22500
rect 142394 22520 142450 22529
rect 142488 22494 142540 22500
rect 142394 22455 142450 22464
rect 142500 22121 142528 22494
rect 174424 22490 174452 44510
rect 174412 22484 174464 22490
rect 174412 22426 174464 22432
rect 142486 22112 142542 22121
rect 142486 22047 142542 22056
rect 137980 21260 138032 21266
rect 137980 21202 138032 21208
rect 138164 21260 138216 21266
rect 138164 21202 138216 21208
rect 139728 21260 139780 21266
rect 139728 21202 139780 21208
rect 143684 21260 143736 21266
rect 143684 21202 143736 21208
rect 135034 20752 135090 20761
rect 135034 20687 135090 20696
rect 134942 19800 134998 19809
rect 134942 19735 134998 19744
rect 101822 19528 101878 19537
rect 101822 19463 101878 19472
rect 134482 19528 134538 19537
rect 134482 19463 134538 19472
rect 106712 18478 106740 18956
rect 112232 18478 112260 18956
rect 106700 18472 106752 18478
rect 106700 18414 106752 18420
rect 112220 18472 112272 18478
rect 112220 18414 112272 18420
rect 96856 17792 96908 17798
rect 96856 17734 96908 17740
rect 88944 17248 88996 17254
rect 88944 17190 88996 17196
rect 87932 17180 87984 17186
rect 87932 17122 87984 17128
rect 85448 12556 85500 12562
rect 85448 12498 85500 12504
rect 88956 12426 88984 17190
rect 88944 12420 88996 12426
rect 88944 12362 88996 12368
rect 90784 12420 90836 12426
rect 90784 12362 90836 12368
rect 90796 9304 90824 12362
rect 96868 9304 96896 17734
rect 117844 17118 117872 18956
rect 126848 17860 126900 17866
rect 126848 17802 126900 17808
rect 120868 17792 120920 17798
rect 120868 17734 120920 17740
rect 117832 17112 117884 17118
rect 117832 17054 117884 17060
rect 102836 12420 102888 12426
rect 102836 12362 102888 12368
rect 102848 9304 102876 12362
rect 108816 12352 108868 12358
rect 108816 12294 108868 12300
rect 108828 9304 108856 12294
rect 114796 12284 114848 12290
rect 114796 12226 114848 12232
rect 114808 9304 114836 12226
rect 120880 9304 120908 17734
rect 126860 9304 126888 17802
rect 129068 17089 129096 18956
rect 138176 18410 138204 21202
rect 143696 21169 143724 21202
rect 143682 21160 143738 21169
rect 143682 21095 143738 21104
rect 146258 21024 146314 21033
rect 147730 21024 147786 21033
rect 146314 20982 146424 21010
rect 147436 20982 147730 21010
rect 146258 20959 146314 20968
rect 148742 21024 148798 21033
rect 148448 20982 148742 21010
rect 147730 20959 147786 20968
rect 150858 21024 150914 21033
rect 150564 20982 150858 21010
rect 148742 20959 148798 20968
rect 150858 20959 150914 20968
rect 145706 20888 145762 20897
rect 145412 20846 145706 20874
rect 149460 20846 149796 20874
rect 151576 20846 151912 20874
rect 145706 20823 145762 20832
rect 138164 18404 138216 18410
rect 138164 18346 138216 18352
rect 138176 18206 138204 18346
rect 149768 18313 149796 20846
rect 149754 18304 149810 18313
rect 149754 18239 149810 18248
rect 138164 18200 138216 18206
rect 138164 18142 138216 18148
rect 132828 17996 132880 18002
rect 132828 17938 132880 17944
rect 129054 17080 129110 17089
rect 129054 17015 129110 17024
rect 132840 9304 132868 17938
rect 138808 17928 138860 17934
rect 138808 17870 138860 17876
rect 138820 9304 138848 17870
rect 150860 17180 150912 17186
rect 150860 17122 150912 17128
rect 144788 12284 144840 12290
rect 144788 12226 144840 12232
rect 144800 9304 144828 12226
rect 150872 9304 150900 17122
rect 151884 17118 151912 20846
rect 152252 20846 152588 20874
rect 153448 20846 153600 20874
rect 154368 20846 154704 20874
rect 155380 20846 155716 20874
rect 156392 20846 156728 20874
rect 157588 20846 157740 20874
rect 158508 20846 158844 20874
rect 159520 20846 159856 20874
rect 160348 20846 160868 20874
rect 161820 20846 161880 20874
rect 162924 20846 162984 20874
rect 163996 20846 164332 20874
rect 152252 18478 152280 20846
rect 153448 18478 153476 20846
rect 152240 18472 152292 18478
rect 152240 18414 152292 18420
rect 153436 18472 153488 18478
rect 153436 18414 153488 18420
rect 153448 18274 153476 18414
rect 153436 18268 153488 18274
rect 153436 18210 153488 18216
rect 154368 17186 154396 20846
rect 154356 17180 154408 17186
rect 154356 17122 154408 17128
rect 151872 17112 151924 17118
rect 151872 17054 151924 17060
rect 155380 12290 155408 20846
rect 156392 17934 156420 20846
rect 157588 18002 157616 20846
rect 157576 17996 157628 18002
rect 157576 17938 157628 17944
rect 156380 17928 156432 17934
rect 156380 17870 156432 17876
rect 158508 17866 158536 20846
rect 158496 17860 158548 17866
rect 158496 17802 158548 17808
rect 159520 17798 159548 20846
rect 159508 17792 159560 17798
rect 159508 17734 159560 17740
rect 160348 12630 160376 20846
rect 161820 12766 161848 20846
rect 162924 17594 162952 20846
rect 164304 18274 164332 20846
rect 164672 20846 165008 20874
rect 165868 20846 166020 20874
rect 166788 20846 167124 20874
rect 167800 20846 168136 20874
rect 168628 20846 169148 20874
rect 170100 20846 170160 20874
rect 170928 20846 171264 20874
rect 171940 20846 172276 20874
rect 164292 18268 164344 18274
rect 164292 18210 164344 18216
rect 162912 17588 162964 17594
rect 162912 17530 162964 17536
rect 164672 17458 164700 20846
rect 162820 17452 162872 17458
rect 162820 17394 162872 17400
rect 164660 17452 164712 17458
rect 164660 17394 164712 17400
rect 161808 12760 161860 12766
rect 161808 12702 161860 12708
rect 160336 12624 160388 12630
rect 160336 12566 160388 12572
rect 155368 12284 155420 12290
rect 155368 12226 155420 12232
rect 156840 12284 156892 12290
rect 156840 12226 156892 12232
rect 156852 9304 156880 12226
rect 162832 9304 162860 17394
rect 165868 12290 165896 20846
rect 166788 18342 166816 20846
rect 165948 18336 166000 18342
rect 165948 18278 166000 18284
rect 166776 18336 166828 18342
rect 166776 18278 166828 18284
rect 165960 15706 165988 18278
rect 167800 18002 167828 20846
rect 168524 18268 168576 18274
rect 168524 18210 168576 18216
rect 167236 17996 167288 18002
rect 167236 17938 167288 17944
rect 167788 17996 167840 18002
rect 167788 17938 167840 17944
rect 167144 17588 167196 17594
rect 167144 17530 167196 17536
rect 165960 15678 166172 15706
rect 166144 12290 166172 15678
rect 167156 12834 167184 17530
rect 167144 12828 167196 12834
rect 167144 12770 167196 12776
rect 167248 12358 167276 17938
rect 167236 12352 167288 12358
rect 167236 12294 167288 12300
rect 168536 12306 168564 18210
rect 168628 12426 168656 20846
rect 169996 17588 170048 17594
rect 169996 17530 170048 17536
rect 170008 12562 170036 17530
rect 169996 12556 170048 12562
rect 169996 12498 170048 12504
rect 170100 12494 170128 20846
rect 170928 17594 170956 20846
rect 171940 18342 171968 20846
rect 176172 19838 176200 46090
rect 177264 40572 177316 40578
rect 177264 40514 177316 40520
rect 177276 39665 177304 40514
rect 177262 39656 177318 39665
rect 177262 39591 177318 39600
rect 177356 39144 177408 39150
rect 177356 39086 177408 39092
rect 177368 37897 177396 39086
rect 177448 39076 177500 39082
rect 177448 39018 177500 39024
rect 177460 38441 177488 39018
rect 177446 38432 177502 38441
rect 177446 38367 177502 38376
rect 177354 37888 177410 37897
rect 177354 37823 177410 37832
rect 177448 37376 177500 37382
rect 177448 37318 177500 37324
rect 177460 37217 177488 37318
rect 177446 37208 177502 37217
rect 177446 37143 177502 37152
rect 177356 36424 177408 36430
rect 177356 36366 177408 36372
rect 177368 35449 177396 36366
rect 177354 35440 177410 35449
rect 177354 35375 177410 35384
rect 176988 32208 177040 32214
rect 176988 32150 177040 32156
rect 177000 31913 177028 32150
rect 176986 31904 177042 31913
rect 176986 31839 177042 31848
rect 177172 30916 177224 30922
rect 177172 30858 177224 30864
rect 177184 30145 177212 30858
rect 177448 30848 177500 30854
rect 177448 30790 177500 30796
rect 177460 30689 177488 30790
rect 177446 30680 177502 30689
rect 177446 30615 177502 30624
rect 177170 30136 177226 30145
rect 177170 30071 177226 30080
rect 177448 28196 177500 28202
rect 177448 28138 177500 28144
rect 177264 28060 177316 28066
rect 177264 28002 177316 28008
rect 177276 27153 177304 28002
rect 177262 27144 177318 27153
rect 177262 27079 177318 27088
rect 177460 26473 177488 28138
rect 177446 26464 177502 26473
rect 177446 26399 177502 26408
rect 177356 25408 177408 25414
rect 177356 25350 177408 25356
rect 177368 24161 177396 25350
rect 177354 24152 177410 24161
rect 177552 24138 177580 46158
rect 185818 46119 185874 46128
rect 185174 45504 185230 45513
rect 185174 45439 185230 45448
rect 185188 45338 185216 45439
rect 181036 45332 181088 45338
rect 181036 45274 181088 45280
rect 185176 45332 185228 45338
rect 185176 45274 185228 45280
rect 177724 44720 177776 44726
rect 177724 44662 177776 44668
rect 177736 44425 177764 44662
rect 177722 44416 177778 44425
rect 177722 44351 177778 44360
rect 181048 43910 181076 45274
rect 185450 44960 185506 44969
rect 185450 44895 185506 44904
rect 177724 43904 177776 43910
rect 177722 43872 177724 43881
rect 181036 43904 181088 43910
rect 177776 43872 177778 43881
rect 181036 43846 181088 43852
rect 177722 43807 177778 43816
rect 185174 43736 185230 43745
rect 185174 43671 185230 43680
rect 184990 43464 185046 43473
rect 184990 43399 185046 43408
rect 181772 43360 181824 43366
rect 181772 43302 181824 43308
rect 177724 43292 177776 43298
rect 177724 43234 177776 43240
rect 177632 43224 177684 43230
rect 177736 43201 177764 43234
rect 177632 43166 177684 43172
rect 177722 43192 177778 43201
rect 177644 42657 177672 43166
rect 177722 43127 177778 43136
rect 177630 42648 177686 42657
rect 177630 42583 177686 42592
rect 181784 42482 181812 43302
rect 177724 42476 177776 42482
rect 177724 42418 177776 42424
rect 181772 42476 181824 42482
rect 181772 42418 181824 42424
rect 177736 42113 177764 42418
rect 177722 42104 177778 42113
rect 177722 42039 177778 42048
rect 177632 41932 177684 41938
rect 177632 41874 177684 41880
rect 177644 40889 177672 41874
rect 185004 41870 185032 43399
rect 185188 43366 185216 43671
rect 185176 43360 185228 43366
rect 185176 43302 185228 43308
rect 185464 43298 185492 44895
rect 185542 44824 185598 44833
rect 185542 44759 185598 44768
rect 185452 43292 185504 43298
rect 185452 43234 185504 43240
rect 185556 43230 185584 44759
rect 185832 44726 185860 46119
rect 185820 44720 185872 44726
rect 185820 44662 185872 44668
rect 185544 43224 185596 43230
rect 185544 43166 185596 43172
rect 185174 42512 185230 42521
rect 185174 42447 185230 42456
rect 185082 42104 185138 42113
rect 185082 42039 185138 42048
rect 177724 41864 177776 41870
rect 177724 41806 177776 41812
rect 184992 41864 185044 41870
rect 184992 41806 185044 41812
rect 177736 41433 177764 41806
rect 177722 41424 177778 41433
rect 177722 41359 177778 41368
rect 177630 40880 177686 40889
rect 177630 40815 177686 40824
rect 184990 40608 185046 40617
rect 184990 40543 185046 40552
rect 177724 40504 177776 40510
rect 177724 40446 177776 40452
rect 177736 40209 177764 40446
rect 177722 40200 177778 40209
rect 177722 40135 177778 40144
rect 177722 39112 177778 39121
rect 177722 39047 177778 39056
rect 177736 39014 177764 39047
rect 185004 39014 185032 40543
rect 185096 40510 185124 42039
rect 185188 41938 185216 42447
rect 185176 41932 185228 41938
rect 185176 41874 185228 41880
rect 185174 41288 185230 41297
rect 185174 41223 185230 41232
rect 185188 40578 185216 41223
rect 185176 40572 185228 40578
rect 185176 40514 185228 40520
rect 185084 40504 185136 40510
rect 185084 40446 185136 40452
rect 185266 40064 185322 40073
rect 185266 39999 185322 40008
rect 185174 39384 185230 39393
rect 185174 39319 185230 39328
rect 185188 39150 185216 39319
rect 185176 39144 185228 39150
rect 185176 39086 185228 39092
rect 185280 39082 185308 39999
rect 185268 39076 185320 39082
rect 185268 39018 185320 39024
rect 177724 39008 177776 39014
rect 177724 38950 177776 38956
rect 184992 39008 185044 39014
rect 184992 38950 185044 38956
rect 185266 38840 185322 38849
rect 185266 38775 185322 38784
rect 185280 38198 185308 38775
rect 183704 38192 183756 38198
rect 185268 38192 185320 38198
rect 183704 38134 183756 38140
rect 185174 38160 185230 38169
rect 183244 37852 183296 37858
rect 183244 37794 183296 37800
rect 183256 36906 183284 37794
rect 183716 37382 183744 38134
rect 185268 38134 185320 38140
rect 185174 38095 185230 38104
rect 184990 37888 185046 37897
rect 185188 37858 185216 38095
rect 184990 37823 185046 37832
rect 185176 37852 185228 37858
rect 183704 37376 183756 37382
rect 183704 37318 183756 37324
rect 177724 36900 177776 36906
rect 177724 36842 177776 36848
rect 183244 36900 183296 36906
rect 183244 36842 183296 36848
rect 177736 36673 177764 36842
rect 177722 36664 177778 36673
rect 177722 36599 177778 36608
rect 185004 36362 185032 37823
rect 185176 37794 185228 37800
rect 185174 36936 185230 36945
rect 185174 36871 185230 36880
rect 185082 36528 185138 36537
rect 185082 36463 185138 36472
rect 177724 36356 177776 36362
rect 177724 36298 177776 36304
rect 184992 36356 185044 36362
rect 184992 36298 185044 36304
rect 177736 36129 177764 36298
rect 177722 36120 177778 36129
rect 177722 36055 177778 36064
rect 184898 35304 184954 35313
rect 184898 35239 184954 35248
rect 177632 35064 177684 35070
rect 177632 35006 177684 35012
rect 177644 34225 177672 35006
rect 177724 34996 177776 35002
rect 177724 34938 177776 34944
rect 177736 34905 177764 34938
rect 177722 34896 177778 34905
rect 177722 34831 177778 34840
rect 177630 34216 177686 34225
rect 177630 34151 177686 34160
rect 177630 33672 177686 33681
rect 177630 33607 177686 33616
rect 177816 33636 177868 33642
rect 177644 33506 177672 33607
rect 177816 33578 177868 33584
rect 177724 33568 177776 33574
rect 177724 33510 177776 33516
rect 177632 33500 177684 33506
rect 177632 33442 177684 33448
rect 177736 33137 177764 33510
rect 177722 33128 177778 33137
rect 177722 33063 177778 33072
rect 177828 32457 177856 33578
rect 184912 33506 184940 35239
rect 185096 35002 185124 36463
rect 185188 36430 185216 36871
rect 185176 36424 185228 36430
rect 185176 36366 185228 36372
rect 185450 35712 185506 35721
rect 185450 35647 185506 35656
rect 185464 35070 185492 35647
rect 185452 35064 185504 35070
rect 185452 35006 185504 35012
rect 185084 34996 185136 35002
rect 185084 34938 185136 34944
rect 185266 34488 185322 34497
rect 185266 34423 185322 34432
rect 185174 33944 185230 33953
rect 185174 33879 185230 33888
rect 184990 33808 185046 33817
rect 184990 33743 185046 33752
rect 184900 33500 184952 33506
rect 184900 33442 184952 33448
rect 177814 32448 177870 32457
rect 177814 32383 177870 32392
rect 177724 32276 177776 32282
rect 177724 32218 177776 32224
rect 177736 31233 177764 32218
rect 185004 32214 185032 33743
rect 185188 33642 185216 33879
rect 185176 33636 185228 33642
rect 185176 33578 185228 33584
rect 185280 33574 185308 34423
rect 185268 33568 185320 33574
rect 185268 33510 185320 33516
rect 215640 33386 215668 69754
rect 222252 48868 222304 48874
rect 222252 48810 222304 48816
rect 222264 48097 222292 48810
rect 222250 48088 222306 48097
rect 222250 48023 222306 48032
rect 215718 33400 215774 33409
rect 215640 33358 215718 33386
rect 215718 33335 215774 33344
rect 185174 32720 185230 32729
rect 185174 32655 185230 32664
rect 185082 32312 185138 32321
rect 185188 32282 185216 32655
rect 185082 32247 185138 32256
rect 185176 32276 185228 32282
rect 184992 32208 185044 32214
rect 184992 32150 185044 32156
rect 177722 31224 177778 31233
rect 177722 31159 177778 31168
rect 184990 30952 185046 30961
rect 184990 30887 185046 30896
rect 177816 29488 177868 29494
rect 177722 29456 177778 29465
rect 177632 29420 177684 29426
rect 177816 29430 177868 29436
rect 177722 29391 177778 29400
rect 177632 29362 177684 29368
rect 177644 28241 177672 29362
rect 177736 29358 177764 29391
rect 177724 29352 177776 29358
rect 177724 29294 177776 29300
rect 177828 28921 177856 29430
rect 185004 29358 185032 30887
rect 185096 30854 185124 32247
rect 185176 32218 185228 32224
rect 185174 31496 185230 31505
rect 185174 31431 185230 31440
rect 185188 30922 185216 31431
rect 185176 30916 185228 30922
rect 185176 30858 185228 30864
rect 185084 30848 185136 30854
rect 185084 30790 185136 30796
rect 185266 30272 185322 30281
rect 185266 30207 185322 30216
rect 185174 29728 185230 29737
rect 185174 29663 185230 29672
rect 185188 29426 185216 29663
rect 185280 29494 185308 30207
rect 185268 29488 185320 29494
rect 185268 29430 185320 29436
rect 185176 29420 185228 29426
rect 185176 29362 185228 29368
rect 184992 29352 185044 29358
rect 184992 29294 185044 29300
rect 185358 29048 185414 29057
rect 185358 28983 185414 28992
rect 177814 28912 177870 28921
rect 177814 28847 177870 28856
rect 185266 28504 185322 28513
rect 185266 28439 185322 28448
rect 177630 28232 177686 28241
rect 177630 28167 177686 28176
rect 185174 28232 185230 28241
rect 185174 28167 185176 28176
rect 185228 28167 185230 28176
rect 185176 28138 185228 28144
rect 177724 28128 177776 28134
rect 177724 28070 177776 28076
rect 177736 27697 177764 28070
rect 185280 28066 185308 28439
rect 185372 28134 185400 28983
rect 185360 28128 185412 28134
rect 185360 28070 185412 28076
rect 185268 28060 185320 28066
rect 185268 28002 185320 28008
rect 177722 27688 177778 27697
rect 177722 27623 177778 27632
rect 185174 27280 185230 27289
rect 185174 27215 185230 27224
rect 185188 26842 185216 27215
rect 185358 26872 185414 26881
rect 185176 26836 185228 26842
rect 185358 26807 185414 26816
rect 185176 26778 185228 26784
rect 177724 26768 177776 26774
rect 177724 26710 177776 26716
rect 177736 25929 177764 26710
rect 177722 25920 177778 25929
rect 177722 25855 177778 25864
rect 185372 25346 185400 26807
rect 185542 26056 185598 26065
rect 185542 25991 185598 26000
rect 185450 25648 185506 25657
rect 185450 25583 185506 25592
rect 185464 25414 185492 25583
rect 185452 25408 185504 25414
rect 185452 25350 185504 25356
rect 177724 25340 177776 25346
rect 177724 25282 177776 25288
rect 185360 25340 185412 25346
rect 185360 25282 185412 25288
rect 177632 25272 177684 25278
rect 177736 25249 177764 25282
rect 185556 25278 185584 25991
rect 185544 25272 185596 25278
rect 177632 25214 177684 25220
rect 177722 25240 177778 25249
rect 177644 24705 177672 25214
rect 185544 25214 185596 25220
rect 177722 25175 177778 25184
rect 185266 24832 185322 24841
rect 185266 24767 185322 24776
rect 177630 24696 177686 24705
rect 177630 24631 177686 24640
rect 185174 24152 185230 24161
rect 177552 24110 177856 24138
rect 177354 24087 177410 24096
rect 177540 23980 177592 23986
rect 177540 23922 177592 23928
rect 177552 22937 177580 23922
rect 177724 23912 177776 23918
rect 177724 23854 177776 23860
rect 177736 23481 177764 23854
rect 177722 23472 177778 23481
rect 177722 23407 177778 23416
rect 177538 22928 177594 22937
rect 177538 22863 177594 22872
rect 177632 22620 177684 22626
rect 177632 22562 177684 22568
rect 177644 22257 177672 22562
rect 177724 22552 177776 22558
rect 177724 22494 177776 22500
rect 177630 22248 177686 22257
rect 177630 22183 177686 22192
rect 177736 21713 177764 22494
rect 177722 21704 177778 21713
rect 177722 21639 177778 21648
rect 177724 21260 177776 21266
rect 177724 21202 177776 21208
rect 177736 21169 177764 21202
rect 177722 21160 177778 21169
rect 177722 21095 177778 21104
rect 176160 19832 176212 19838
rect 176160 19774 176212 19780
rect 177828 19770 177856 24110
rect 185174 24087 185230 24096
rect 185188 23986 185216 24087
rect 185176 23980 185228 23986
rect 185176 23922 185228 23928
rect 185280 23918 185308 24767
rect 185268 23912 185320 23918
rect 185268 23854 185320 23860
rect 185266 23608 185322 23617
rect 185266 23543 185322 23552
rect 185174 22928 185230 22937
rect 185174 22863 185230 22872
rect 185188 22694 185216 22863
rect 185280 22830 185308 23543
rect 185268 22824 185320 22830
rect 185268 22766 185320 22772
rect 185176 22688 185228 22694
rect 185176 22630 185228 22636
rect 185266 22656 185322 22665
rect 185266 22591 185322 22600
rect 185176 22484 185228 22490
rect 185176 22426 185228 22432
rect 185188 22393 185216 22426
rect 185174 22384 185230 22393
rect 185174 22319 185230 22328
rect 185280 21266 185308 22591
rect 185268 21260 185320 21266
rect 185268 21202 185320 21208
rect 185268 19832 185320 19838
rect 185174 19800 185230 19809
rect 177816 19764 177868 19770
rect 185268 19774 185320 19780
rect 185174 19735 185176 19744
rect 177816 19706 177868 19712
rect 185228 19735 185230 19744
rect 185176 19706 185228 19712
rect 185280 19537 185308 19774
rect 185266 19528 185322 19537
rect 185266 19463 185322 19472
rect 194940 18478 194968 18956
rect 194928 18472 194980 18478
rect 194928 18414 194980 18420
rect 171376 18336 171428 18342
rect 171376 18278 171428 18284
rect 171928 18336 171980 18342
rect 171928 18278 171980 18284
rect 170916 17588 170968 17594
rect 170916 17530 170968 17536
rect 171388 12698 171416 18278
rect 208924 17118 208952 18956
rect 212500 18472 212552 18478
rect 212498 18440 212500 18449
rect 212552 18440 212554 18449
rect 212498 18375 212554 18384
rect 208912 17112 208964 17118
rect 208912 17054 208964 17060
rect 174872 12828 174924 12834
rect 174872 12770 174924 12776
rect 171376 12692 171428 12698
rect 171376 12634 171428 12640
rect 170088 12488 170140 12494
rect 170088 12430 170140 12436
rect 168616 12420 168668 12426
rect 168616 12362 168668 12368
rect 165856 12284 165908 12290
rect 165856 12226 165908 12232
rect 166132 12284 166184 12290
rect 168536 12278 168840 12306
rect 166132 12226 166184 12232
rect 168812 9304 168840 12278
rect 174884 9304 174912 12770
rect 180852 12760 180904 12766
rect 180852 12702 180904 12708
rect 180864 9304 180892 12702
rect 192812 12692 192864 12698
rect 192812 12634 192864 12640
rect 186832 12624 186884 12630
rect 186832 12566 186884 12572
rect 186844 9304 186872 12566
rect 192824 9304 192852 12634
rect 198792 12556 198844 12562
rect 198792 12498 198844 12504
rect 198804 9304 198832 12498
rect 204864 12488 204916 12494
rect 204864 12430 204916 12436
rect 204876 9304 204904 12430
rect 210844 12420 210896 12426
rect 210844 12362 210896 12368
rect 210856 9304 210884 12362
rect 216824 12352 216876 12358
rect 216824 12294 216876 12300
rect 216836 9304 216864 12294
rect 222804 12284 222856 12290
rect 222804 12226 222856 12232
rect 222816 9304 222844 12226
rect 12858 8824 12914 9304
rect 18838 8824 18894 9304
rect 24818 8824 24874 9304
rect 30798 8824 30854 9304
rect 36778 8824 36834 9304
rect 42850 8824 42906 9304
rect 48830 8824 48886 9304
rect 54810 8824 54866 9304
rect 60790 8824 60846 9304
rect 66862 8824 66918 9304
rect 72842 8824 72898 9304
rect 78822 8824 78878 9304
rect 84802 8824 84858 9304
rect 90782 8824 90838 9304
rect 96854 8824 96910 9304
rect 102834 8824 102890 9304
rect 108814 8824 108870 9304
rect 114794 8824 114850 9304
rect 120866 8824 120922 9304
rect 126846 8824 126902 9304
rect 132826 8824 132882 9304
rect 138806 8824 138862 9304
rect 144786 8824 144842 9304
rect 150858 8824 150914 9304
rect 156838 8824 156894 9304
rect 162818 8824 162874 9304
rect 168798 8824 168854 9304
rect 174870 8824 174926 9304
rect 180850 8824 180906 9304
rect 186830 8824 186886 9304
rect 192810 8824 192866 9304
rect 198790 8824 198846 9304
rect 204862 8824 204918 9304
rect 210842 8824 210898 9304
rect 216822 8824 216878 9304
rect 222802 8824 222858 9304
<< via2 >>
rect 12766 232856 12822 232912
rect 18102 220888 18158 220944
rect 13318 209328 13374 209384
rect 50670 234488 50726 234544
rect 49934 233944 49990 234000
rect 50578 233400 50634 233456
rect 58122 232992 58178 233048
rect 51222 232856 51278 232912
rect 79558 235168 79614 235224
rect 134758 234488 134814 234544
rect 101638 234080 101694 234136
rect 100994 233128 101050 233184
rect 100994 232584 101050 232640
rect 51130 232176 51186 232232
rect 51222 231632 51278 231688
rect 51222 231108 51278 231144
rect 51222 231088 51224 231108
rect 51224 231088 51276 231108
rect 51276 231088 51278 231108
rect 51130 230544 51186 230600
rect 51222 230000 51278 230056
rect 92714 232448 92770 232504
rect 100994 232040 101050 232096
rect 58122 231904 58178 231960
rect 94002 231904 94058 231960
rect 100994 231496 101050 231552
rect 58030 231224 58086 231280
rect 92714 231224 92770 231280
rect 58214 230680 58270 230736
rect 92714 230680 92770 230736
rect 101086 231088 101142 231144
rect 58306 230136 58362 230192
rect 94094 230136 94150 230192
rect 101086 230136 101142 230192
rect 51130 229320 51186 229376
rect 50762 228776 50818 228832
rect 100994 229728 101050 229784
rect 58214 229456 58270 229512
rect 92714 229456 92770 229512
rect 58214 228912 58270 228968
rect 51222 228268 51224 228288
rect 51224 228268 51276 228288
rect 51276 228268 51278 228288
rect 50486 225920 50542 225976
rect 50210 220208 50266 220264
rect 50210 219120 50266 219176
rect 50394 215040 50450 215096
rect 50210 213428 50266 213464
rect 50210 213408 50212 213428
rect 50212 213408 50264 213428
rect 50264 213408 50266 213428
rect 51222 228232 51278 228268
rect 50946 227688 51002 227744
rect 51222 227144 51278 227200
rect 50762 226464 50818 226520
rect 100994 229184 101050 229240
rect 93174 228912 93230 228968
rect 101086 228640 101142 228696
rect 58306 228232 58362 228288
rect 92714 228232 92770 228288
rect 100994 228232 101050 228288
rect 58214 227688 58270 227744
rect 93174 227688 93230 227744
rect 101086 227416 101142 227472
rect 58306 227144 58362 227200
rect 92714 227144 92770 227200
rect 100994 227008 101050 227064
rect 58214 226464 58270 226520
rect 92714 226464 92770 226520
rect 101086 226328 101142 226384
rect 58306 225920 58362 225976
rect 93634 225920 93690 225976
rect 51130 225376 51186 225432
rect 51038 224308 51094 224344
rect 51038 224288 51040 224308
rect 51040 224288 51092 224308
rect 51092 224288 51094 224308
rect 58214 225240 58270 225296
rect 51222 224832 51278 224888
rect 58306 224696 58362 224752
rect 50946 223608 51002 223664
rect 51222 223084 51278 223120
rect 51222 223064 51224 223084
rect 51224 223064 51276 223084
rect 51276 223064 51278 223084
rect 100994 225512 101050 225568
rect 101178 225648 101234 225704
rect 92806 225240 92862 225296
rect 92714 224696 92770 224752
rect 101086 224560 101142 224616
rect 58398 224152 58454 224208
rect 92898 224152 92954 224208
rect 100994 224152 101050 224208
rect 58214 223472 58270 223528
rect 51130 222520 51186 222576
rect 51222 221976 51278 222032
rect 51222 221452 51278 221488
rect 51222 221432 51224 221452
rect 51224 221432 51276 221452
rect 51276 221432 51278 221452
rect 50946 220752 51002 220808
rect 93726 223472 93782 223528
rect 101454 223472 101510 223528
rect 58306 222928 58362 222984
rect 93910 222928 93966 222984
rect 101270 222792 101326 222848
rect 58214 222248 58270 222304
rect 92714 222248 92770 222304
rect 58306 221704 58362 221760
rect 92990 221704 93046 221760
rect 58214 221160 58270 221216
rect 92714 221180 92770 221216
rect 92714 221160 92716 221180
rect 92716 221160 92768 221180
rect 92768 221160 92770 221180
rect 58214 220480 58270 220536
rect 50854 219664 50910 219720
rect 51222 218576 51278 218632
rect 51222 217896 51278 217952
rect 51222 217372 51278 217408
rect 51222 217352 51224 217372
rect 51224 217352 51276 217372
rect 51276 217352 51278 217372
rect 101546 223064 101602 223120
rect 101546 221840 101602 221896
rect 93726 220480 93782 220536
rect 58306 219936 58362 219992
rect 93174 219936 93230 219992
rect 58214 219256 58270 219312
rect 51130 216808 51186 216864
rect 51222 216264 51278 216320
rect 51222 215720 51278 215776
rect 51130 214532 51132 214552
rect 51132 214532 51184 214552
rect 51184 214532 51186 214552
rect 51130 214496 51186 214532
rect 92806 219256 92862 219312
rect 58306 218712 58362 218768
rect 92714 218712 92770 218768
rect 58214 218168 58270 218224
rect 92806 218168 92862 218224
rect 58214 217488 58270 217544
rect 93726 217488 93782 217544
rect 58214 216944 58270 217000
rect 93910 216944 93966 217000
rect 58306 216264 58362 216320
rect 92714 216264 92770 216320
rect 58214 215740 58270 215776
rect 58214 215720 58216 215740
rect 58216 215720 58268 215740
rect 58268 215720 58270 215740
rect 92714 215740 92770 215776
rect 92714 215720 92716 215740
rect 92716 215720 92768 215740
rect 92768 215720 92770 215740
rect 58306 215176 58362 215232
rect 92806 215176 92862 215232
rect 50946 213952 51002 214008
rect 58214 214496 58270 214552
rect 93542 214496 93598 214552
rect 58214 213952 58270 214008
rect 50762 212864 50818 212920
rect 51222 212184 51278 212240
rect 51130 211640 51186 211696
rect 50670 211096 50726 211152
rect 22334 190424 22390 190480
rect 50854 210552 50910 210608
rect 50762 210008 50818 210064
rect 92806 213952 92862 214008
rect 58306 213272 58362 213328
rect 92714 213272 92770 213328
rect 58214 212728 58270 212784
rect 92714 212728 92770 212784
rect 58306 212184 58362 212240
rect 93634 212184 93690 212240
rect 58214 211504 58270 211560
rect 92714 211524 92770 211560
rect 92714 211504 92716 211524
rect 92716 211504 92768 211524
rect 92768 211504 92770 211524
rect 58306 210960 58362 211016
rect 92806 210960 92862 211016
rect 58398 210280 58454 210336
rect 100994 215040 101050 215096
rect 100994 213952 101050 214008
rect 58214 209736 58270 209792
rect 50946 209328 51002 209384
rect 58306 209192 58362 209248
rect 51130 208784 51186 208840
rect 51038 208240 51094 208296
rect 51222 207716 51278 207752
rect 51222 207696 51224 207716
rect 51224 207696 51276 207716
rect 51276 207696 51278 207716
rect 51130 207152 51186 207208
rect 85722 207424 85778 207480
rect 93542 210280 93598 210336
rect 92714 209736 92770 209792
rect 101178 213408 101234 213464
rect 101086 213156 101142 213192
rect 101086 213136 101088 213156
rect 101088 213136 101140 213156
rect 101140 213136 101142 213156
rect 100994 212320 101050 212376
rect 101086 211912 101142 211968
rect 101178 211096 101234 211152
rect 101086 210688 101142 210744
rect 100994 210416 101050 210472
rect 101086 209464 101142 209520
rect 94094 209192 94150 209248
rect 100994 209056 101050 209112
rect 134298 233400 134354 233456
rect 134574 225920 134630 225976
rect 134482 221976 134538 222032
rect 101730 221432 101786 221488
rect 101730 220616 101786 220672
rect 101822 220208 101878 220264
rect 101914 219936 101970 219992
rect 101730 218984 101786 219040
rect 102006 218576 102062 218632
rect 101914 217896 101970 217952
rect 101822 217488 101878 217544
rect 101730 217236 101786 217272
rect 101730 217216 101732 217236
rect 101732 217216 101784 217236
rect 101784 217216 101786 217236
rect 101822 216128 101878 216184
rect 101730 215992 101786 216048
rect 101822 214904 101878 214960
rect 134666 213952 134722 214008
rect 102098 208376 102154 208432
rect 101914 207832 101970 207888
rect 101730 207560 101786 207616
rect 100994 206472 101050 206528
rect 41838 189200 41894 189256
rect 13410 185664 13466 185720
rect 99246 190696 99302 190752
rect 99154 189472 99210 189528
rect 135402 233964 135458 234000
rect 135402 233944 135404 233964
rect 135404 233944 135456 233964
rect 135456 233944 135458 233964
rect 142302 232992 142358 233048
rect 135402 232856 135458 232912
rect 194926 236528 194982 236584
rect 186002 234488 186058 234544
rect 185082 233944 185138 234000
rect 185174 233400 185230 233456
rect 177170 232992 177226 233048
rect 135402 232176 135458 232232
rect 134850 231632 134906 231688
rect 135310 231108 135366 231144
rect 135310 231088 135312 231108
rect 135312 231088 135364 231108
rect 135364 231088 135366 231108
rect 135402 230544 135458 230600
rect 135310 230020 135366 230056
rect 135310 230000 135312 230020
rect 135312 230000 135364 230020
rect 135364 230000 135366 230020
rect 163554 232584 163610 232640
rect 177722 232176 177778 232232
rect 142302 231904 142358 231960
rect 185266 232856 185322 232912
rect 185266 232176 185322 232232
rect 185174 231632 185230 231688
rect 177722 231496 177778 231552
rect 142210 231224 142266 231280
rect 143682 230680 143738 230736
rect 178182 230816 178238 230872
rect 185358 231088 185414 231144
rect 185266 230544 185322 230600
rect 177722 230408 177778 230464
rect 142946 230136 143002 230192
rect 185174 230000 185230 230056
rect 135402 229320 135458 229376
rect 135310 228776 135366 228832
rect 135402 228268 135404 228288
rect 135404 228268 135456 228288
rect 135456 228268 135458 228288
rect 135402 228232 135458 228268
rect 143682 229492 143684 229512
rect 143684 229492 143736 229512
rect 143736 229492 143738 229512
rect 143682 229456 143738 229492
rect 177722 229320 177778 229376
rect 177630 229184 177686 229240
rect 143590 228912 143646 228968
rect 185634 229320 185690 229376
rect 177814 228640 177870 228696
rect 135402 227688 135458 227744
rect 135310 227144 135366 227200
rect 143498 228232 143554 228288
rect 185174 228268 185176 228288
rect 185176 228268 185228 228288
rect 185228 228268 185230 228288
rect 143682 227688 143738 227744
rect 177722 227960 177778 228016
rect 177630 227416 177686 227472
rect 143314 227144 143370 227200
rect 135218 226464 135274 226520
rect 143682 226464 143738 226520
rect 185174 228232 185230 228268
rect 185910 228776 185966 228832
rect 185174 227688 185230 227744
rect 177722 226636 177724 226656
rect 177724 226636 177776 226656
rect 177776 226636 177778 226656
rect 177722 226600 177778 226636
rect 177630 226192 177686 226248
rect 143314 225920 143370 225976
rect 135310 225376 135366 225432
rect 135218 224308 135274 224344
rect 135218 224288 135220 224308
rect 135220 224288 135272 224308
rect 135272 224288 135274 224308
rect 135402 224832 135458 224888
rect 135402 223608 135458 223664
rect 135310 223084 135366 223120
rect 135310 223064 135312 223084
rect 135312 223064 135364 223084
rect 135364 223064 135366 223084
rect 143682 225240 143738 225296
rect 177722 225376 177778 225432
rect 177630 224968 177686 225024
rect 143590 224696 143646 224752
rect 185266 227144 185322 227200
rect 185174 226464 185230 226520
rect 185266 225920 185322 225976
rect 185358 225376 185414 225432
rect 185174 224832 185230 224888
rect 177814 224424 177870 224480
rect 143498 224152 143554 224208
rect 134850 222520 134906 222576
rect 135310 221452 135366 221488
rect 135310 221432 135312 221452
rect 135312 221432 135364 221452
rect 135364 221432 135366 221452
rect 135402 220752 135458 220808
rect 135310 220208 135366 220264
rect 143682 223472 143738 223528
rect 185266 224288 185322 224344
rect 177722 223744 177778 223800
rect 185174 223608 185230 223664
rect 177354 223200 177410 223256
rect 143314 222928 143370 222984
rect 143682 222248 143738 222304
rect 185450 223064 185506 223120
rect 185266 222520 185322 222576
rect 177722 222384 177778 222440
rect 177630 221976 177686 222032
rect 185174 221976 185230 222032
rect 143314 221704 143370 221760
rect 143682 221160 143738 221216
rect 185358 221432 185414 221488
rect 177722 221024 177778 221080
rect 177630 220888 177686 220944
rect 143590 220480 143646 220536
rect 135402 219664 135458 219720
rect 135034 219120 135090 219176
rect 135310 218612 135312 218632
rect 135312 218612 135364 218632
rect 135364 218612 135366 218632
rect 135310 218576 135366 218612
rect 135402 217896 135458 217952
rect 135402 217372 135458 217408
rect 135402 217352 135404 217372
rect 135404 217352 135456 217372
rect 135456 217352 135458 217372
rect 135402 216808 135458 216864
rect 135494 216264 135550 216320
rect 135402 215720 135458 215776
rect 134850 215040 134906 215096
rect 135310 214532 135312 214552
rect 135312 214532 135364 214552
rect 135364 214532 135366 214552
rect 135310 214496 135366 214532
rect 185174 220752 185230 220808
rect 177814 220208 177870 220264
rect 143682 219936 143738 219992
rect 143682 219256 143738 219312
rect 185542 220208 185598 220264
rect 177722 219528 177778 219584
rect 177630 218984 177686 219040
rect 143130 218712 143186 218768
rect 185726 219664 185782 219720
rect 185634 219120 185690 219176
rect 143682 218168 143738 218224
rect 177722 218304 177778 218360
rect 177630 217896 177686 217952
rect 143498 217488 143554 217544
rect 185542 217352 185598 217408
rect 177722 217116 177724 217136
rect 177724 217116 177776 217136
rect 177776 217116 177778 217136
rect 177722 217080 177778 217116
rect 143682 216944 143738 217000
rect 177630 216672 177686 216728
rect 143130 216264 143186 216320
rect 143130 215740 143186 215776
rect 143130 215720 143132 215740
rect 143132 215720 143184 215740
rect 143184 215720 143186 215740
rect 142946 215176 143002 215232
rect 135402 213428 135458 213464
rect 135402 213408 135404 213428
rect 135404 213408 135456 213428
rect 135456 213408 135458 213428
rect 134850 212864 134906 212920
rect 135402 212184 135458 212240
rect 135402 211640 135458 211696
rect 135034 211096 135090 211152
rect 134850 210552 134906 210608
rect 99522 193688 99578 193744
rect 134942 209328 134998 209384
rect 177722 215620 177724 215640
rect 177724 215620 177776 215640
rect 177776 215620 177778 215640
rect 177722 215584 177778 215620
rect 177722 215312 177778 215368
rect 177630 214904 177686 214960
rect 143498 214496 143554 214552
rect 142946 213952 143002 214008
rect 177722 214088 177778 214144
rect 177630 213680 177686 213736
rect 143682 213272 143738 213328
rect 215718 230680 215774 230736
rect 185726 217896 185782 217952
rect 185726 216264 185782 216320
rect 185634 215720 185690 215776
rect 185266 214532 185268 214552
rect 185268 214532 185320 214552
rect 185320 214532 185322 214552
rect 177722 212864 177778 212920
rect 143682 212728 143738 212784
rect 185266 214496 185322 214532
rect 185726 215040 185782 215096
rect 185726 213952 185782 214008
rect 185174 213408 185230 213464
rect 177722 212320 177778 212376
rect 143498 212184 143554 212240
rect 177722 211660 177778 211696
rect 177722 211640 177724 211660
rect 177724 211640 177776 211660
rect 177776 211640 177778 211660
rect 143682 211504 143738 211560
rect 177722 211096 177778 211152
rect 143682 210960 143738 211016
rect 177722 210688 177778 210744
rect 143590 210280 143646 210336
rect 135126 210008 135182 210064
rect 142946 209736 143002 209792
rect 143682 209192 143738 209248
rect 135310 208784 135366 208840
rect 135218 208240 135274 208296
rect 135402 207696 135458 207752
rect 135310 207152 135366 207208
rect 169902 208920 169958 208976
rect 167142 195184 167198 195240
rect 177722 209872 177778 209928
rect 178182 209464 178238 209520
rect 185726 212864 185782 212920
rect 185726 211640 185782 211696
rect 185910 218576 185966 218632
rect 185910 216808 185966 216864
rect 185910 212184 185966 212240
rect 222342 231632 222398 231688
rect 220318 220752 220374 220808
rect 216914 211504 216970 211560
rect 185818 211096 185874 211152
rect 185726 210008 185782 210064
rect 185818 209328 185874 209384
rect 186002 210552 186058 210608
rect 186094 208784 186150 208840
rect 186002 207696 186058 207752
rect 185174 207152 185230 207208
rect 182874 193180 182876 193200
rect 182876 193180 182928 193200
rect 182928 193180 182930 193200
rect 182874 193144 182930 193180
rect 105778 192464 105834 192520
rect 99430 192328 99486 192384
rect 99338 188928 99394 188984
rect 99062 187704 99118 187760
rect 98970 186480 99026 186536
rect 98878 185256 98934 185312
rect 22334 183760 22390 183816
rect 98602 182400 98658 182456
rect 99522 183624 99578 183680
rect 99430 181040 99486 181096
rect 99522 179816 99578 179872
rect 107158 190152 107214 190208
rect 106790 187840 106846 187896
rect 106790 185392 106846 185448
rect 183426 190696 183482 190752
rect 183334 189472 183390 189528
rect 186278 208240 186334 208296
rect 187934 206880 187990 206936
rect 191982 192736 192038 192792
rect 183610 191920 183666 191976
rect 191982 188656 192038 188712
rect 183518 188248 183574 188304
rect 183242 187024 183298 187080
rect 183150 185800 183206 185856
rect 183058 184576 183114 184632
rect 191154 186752 191210 186808
rect 128502 183760 128558 183816
rect 107158 183080 107214 183136
rect 182874 183352 182930 183408
rect 106974 180768 107030 180824
rect 98418 179272 98474 179328
rect 44414 178728 44470 178784
rect 22334 177132 22336 177152
rect 22336 177132 22388 177152
rect 22388 177132 22390 177152
rect 22334 177096 22390 177132
rect 99522 177388 99578 177424
rect 106790 178320 106846 178376
rect 99522 177368 99524 177388
rect 99524 177368 99576 177388
rect 99576 177368 99578 177388
rect 98602 176688 98658 176744
rect 106606 176008 106662 176064
rect 98234 175328 98290 175384
rect 190602 182672 190658 182728
rect 191982 184712 192038 184768
rect 183150 182128 183206 182184
rect 183702 181040 183758 181096
rect 183702 179836 183758 179872
rect 190694 180768 190750 180824
rect 183702 179816 183704 179836
rect 183704 179816 183756 179836
rect 183756 179816 183758 179836
rect 191982 178728 192038 178784
rect 182506 178592 182562 178648
rect 182506 177368 182562 177424
rect 191982 176688 192038 176744
rect 183242 176144 183298 176200
rect 183702 174920 183758 174976
rect 191522 174784 191578 174840
rect 137518 174376 137574 174432
rect 52694 173832 52750 173888
rect 99522 173716 99578 173752
rect 99522 173696 99524 173716
rect 99524 173696 99576 173716
rect 99576 173696 99578 173716
rect 106790 173716 106846 173752
rect 106790 173696 106792 173716
rect 106792 173696 106844 173716
rect 106844 173696 106846 173716
rect 183334 173696 183390 173752
rect 191982 172744 192038 172800
rect 99522 172472 99578 172528
rect 183518 172472 183574 172528
rect 106790 171384 106846 171440
rect 99246 171248 99302 171304
rect 182690 171268 182746 171304
rect 182690 171248 182692 171268
rect 182692 171248 182744 171268
rect 182744 171248 182746 171268
rect 22978 170432 23034 170488
rect 99522 170024 99578 170080
rect 182506 170024 182562 170080
rect 106790 168936 106846 168992
rect 99430 168800 99486 168856
rect 44414 168664 44470 168720
rect 99522 167712 99578 167768
rect 23622 163768 23678 163824
rect 13134 162136 13190 162192
rect 209922 190696 209978 190752
rect 212130 190424 212186 190480
rect 212038 183760 212094 183816
rect 211578 177096 211634 177152
rect 209830 170976 209886 171032
rect 191154 170704 191210 170760
rect 183702 168800 183758 168856
rect 106698 166624 106754 166680
rect 99522 166488 99578 166544
rect 99522 165264 99578 165320
rect 106790 164312 106846 164368
rect 99522 164040 99578 164096
rect 98970 162816 99026 162872
rect 53338 160504 53394 160560
rect 44506 158736 44562 158792
rect 23622 157104 23678 157160
rect 98786 154384 98842 154440
rect 49934 140412 49936 140432
rect 49936 140412 49988 140432
rect 49988 140412 49990 140432
rect 49934 140376 49990 140412
rect 49934 140104 49990 140160
rect 49658 139016 49714 139072
rect 13318 138472 13374 138528
rect 49934 138744 49990 138800
rect 50026 137792 50082 137848
rect 49934 137384 49990 137440
rect 51038 136704 51094 136760
rect 51130 136160 51186 136216
rect 51222 135924 51224 135944
rect 51224 135924 51276 135944
rect 51276 135924 51278 135944
rect 51222 135888 51278 135924
rect 51130 134936 51186 134992
rect 51222 134664 51278 134720
rect 50394 133848 50450 133904
rect 18102 133304 18158 133360
rect 18010 119296 18066 119352
rect 13410 114944 13466 115000
rect 51130 133304 51186 133360
rect 51222 133068 51224 133088
rect 51224 133068 51276 133088
rect 51276 133068 51278 133088
rect 51222 133032 51278 133068
rect 51130 132080 51186 132136
rect 51222 131808 51278 131864
rect 50210 130992 50266 131048
rect 51130 130584 51186 130640
rect 51222 130448 51278 130504
rect 51130 129224 51186 129280
rect 51222 128988 51224 129008
rect 51224 128988 51276 129008
rect 51276 128988 51278 129008
rect 51222 128952 51278 128988
rect 50762 128136 50818 128192
rect 51222 127728 51278 127784
rect 50210 126912 50266 126968
rect 50394 126504 50450 126560
rect 51222 126096 51278 126152
rect 51130 125280 51186 125336
rect 51222 125008 51278 125064
rect 50210 124056 50266 124112
rect 51222 123784 51278 123840
rect 51222 123532 51278 123568
rect 51222 123512 51224 123532
rect 51224 123512 51276 123532
rect 51276 123512 51278 123532
rect 51130 122424 51186 122480
rect 51222 122172 51278 122208
rect 51222 122152 51224 122172
rect 51224 122152 51276 122172
rect 51276 122152 51278 122172
rect 51130 121200 51186 121256
rect 51222 120928 51278 120984
rect 50210 120112 50266 120168
rect 51222 119704 51278 119760
rect 51222 119296 51278 119352
rect 50578 118344 50634 118400
rect 51222 118092 51278 118128
rect 51222 118072 51224 118092
rect 51224 118072 51276 118092
rect 51276 118072 51278 118092
rect 50026 117256 50082 117312
rect 50578 116712 50634 116768
rect 50486 113856 50542 113912
rect 22334 96448 22390 96504
rect 50762 116440 50818 116496
rect 50670 115488 50726 115544
rect 50854 115080 50910 115136
rect 51130 114400 51186 114456
rect 50946 113720 51002 113776
rect 51222 112788 51278 112824
rect 51222 112768 51224 112788
rect 51224 112768 51276 112788
rect 51276 112768 51278 112788
rect 58490 138880 58546 138936
rect 58214 136568 58270 136624
rect 92714 138508 92716 138528
rect 92716 138508 92768 138528
rect 92768 138508 92770 138528
rect 92714 138472 92770 138508
rect 58950 138200 59006 138256
rect 92806 138064 92862 138120
rect 58398 137112 58454 137168
rect 92714 137132 92770 137168
rect 92714 137112 92716 137132
rect 92716 137112 92768 137132
rect 92768 137112 92770 137132
rect 92806 136840 92862 136896
rect 92714 136432 92770 136488
rect 58306 136024 58362 136080
rect 92714 135480 92770 135536
rect 58214 135344 58270 135400
rect 92806 135208 92862 135264
rect 58306 134800 58362 134856
rect 58398 134120 58454 134176
rect 58214 133576 58270 133632
rect 58306 133032 58362 133088
rect 92714 134120 92770 134176
rect 92806 133984 92862 134040
rect 92898 133440 92954 133496
rect 92714 132624 92770 132680
rect 58306 132352 58362 132408
rect 92806 132216 92862 132272
rect 58214 131808 58270 131864
rect 58214 131128 58270 131184
rect 58306 130584 58362 130640
rect 92714 131264 92770 131320
rect 92806 130992 92862 131048
rect 58490 130040 58546 130096
rect 92714 130040 92770 130096
rect 92806 129768 92862 129824
rect 58214 129360 58270 129416
rect 58214 128836 58270 128872
rect 58214 128816 58216 128836
rect 58216 128816 58268 128836
rect 58268 128816 58270 128836
rect 92714 128816 92770 128872
rect 92806 128408 92862 128464
rect 58398 128136 58454 128192
rect 92898 128000 92954 128056
rect 58306 127592 58362 127648
rect 58214 126368 58270 126424
rect 92714 127184 92770 127240
rect 58398 127048 58454 127104
rect 92806 126912 92862 126968
rect 92714 125960 92770 126016
rect 58306 125824 58362 125880
rect 92806 125552 92862 125608
rect 58214 125144 58270 125200
rect 58306 124636 58308 124656
rect 58308 124636 58360 124656
rect 58360 124636 58362 124656
rect 58306 124600 58362 124636
rect 58214 123376 58270 123432
rect 92714 124636 92716 124656
rect 92716 124636 92768 124656
rect 92768 124636 92770 124656
rect 92714 124600 92770 124636
rect 92806 124328 92862 124384
rect 58490 124056 58546 124112
rect 92898 123920 92954 123976
rect 92714 122968 92770 123024
rect 58398 122832 58454 122888
rect 92806 122696 92862 122752
rect 58214 122152 58270 122208
rect 92714 121744 92770 121800
rect 58214 121608 58270 121664
rect 92806 121472 92862 121528
rect 58214 121064 58270 121120
rect 58214 120384 58270 120440
rect 58398 119840 58454 119896
rect 58306 119160 58362 119216
rect 92714 120384 92770 120440
rect 92806 119976 92862 120032
rect 92714 119160 92770 119216
rect 92806 118888 92862 118944
rect 58490 118616 58546 118672
rect 92898 118480 92954 118536
rect 58214 118072 58270 118128
rect 58214 117392 58270 117448
rect 92714 117528 92770 117584
rect 92806 117120 92862 117176
rect 58306 116848 58362 116904
rect 58306 116168 58362 116224
rect 58398 115624 58454 115680
rect 58214 115080 58270 115136
rect 41838 95224 41894 95280
rect 13502 91280 13558 91336
rect 22334 89784 22390 89840
rect 44414 84772 44470 84808
rect 44414 84752 44416 84772
rect 44416 84752 44468 84772
rect 44468 84752 44470 84772
rect 22334 83120 22390 83176
rect 52694 79856 52750 79912
rect 22334 76456 22390 76512
rect 44414 74688 44470 74744
rect 92714 116168 92770 116224
rect 92806 115760 92862 115816
rect 92898 115488 92954 115544
rect 23622 69792 23678 69848
rect 53338 66528 53394 66584
rect 44414 64760 44470 64816
rect 23622 63128 23678 63184
rect 59226 58368 59282 58424
rect 50394 46808 50450 46864
rect 13318 44088 13374 44144
rect 50026 43680 50082 43736
rect 50210 42864 50266 42920
rect 18102 39328 18158 39384
rect 50026 35656 50082 35712
rect 50210 34432 50266 34488
rect 50026 32664 50082 32720
rect 50486 26136 50542 26192
rect 18102 25456 18158 25512
rect 13318 20560 13374 20616
rect 50210 23144 50266 23200
rect 50670 21104 50726 21160
rect 50946 21784 51002 21840
rect 51314 45176 51370 45232
rect 51222 44788 51278 44824
rect 51222 44768 51224 44788
rect 51224 44768 51276 44788
rect 51276 44768 51278 44788
rect 79190 58232 79246 58288
rect 98786 99712 98842 99768
rect 98786 89920 98842 89976
rect 98694 87336 98750 87392
rect 98234 75504 98290 75560
rect 99062 161592 99118 161648
rect 99154 160368 99210 160424
rect 99430 159144 99486 159200
rect 99246 157920 99302 157976
rect 99338 156696 99394 156752
rect 99522 155472 99578 155528
rect 183794 167712 183850 167768
rect 182874 166508 182930 166544
rect 182874 166488 182876 166508
rect 182876 166488 182928 166508
rect 182928 166488 182930 166508
rect 106882 161864 106938 161920
rect 183702 165264 183758 165320
rect 183058 164040 183114 164096
rect 128502 163768 128558 163824
rect 183058 162816 183114 162872
rect 137518 160504 137574 160560
rect 107250 159552 107306 159608
rect 107158 157240 107214 157296
rect 137518 156696 137574 156752
rect 106514 154928 106570 154984
rect 134850 140512 134906 140568
rect 100810 140104 100866 140160
rect 100902 139968 100958 140024
rect 135402 139988 135458 140024
rect 135402 139968 135404 139988
rect 135404 139968 135456 139988
rect 135456 139968 135458 139988
rect 134666 139424 134722 139480
rect 101178 138880 101234 138936
rect 101086 138744 101142 138800
rect 135402 138764 135458 138800
rect 135402 138744 135404 138764
rect 135404 138744 135456 138764
rect 135456 138744 135458 138764
rect 134666 138200 134722 138256
rect 101822 137792 101878 137848
rect 101270 137656 101326 137712
rect 135402 137656 135458 137712
rect 135034 136976 135090 137032
rect 101178 136568 101234 136624
rect 101270 136024 101326 136080
rect 135310 136432 135366 136488
rect 101730 135888 101786 135944
rect 135402 135888 135458 135944
rect 134850 135344 134906 135400
rect 101822 134800 101878 134856
rect 100902 134392 100958 134448
rect 134482 134684 134538 134720
rect 134482 134664 134484 134684
rect 134484 134664 134536 134684
rect 134536 134664 134538 134684
rect 135402 134120 135458 134176
rect 101362 133712 101418 133768
rect 135034 133576 135090 133632
rect 101730 133032 101786 133088
rect 101454 131944 101510 132000
rect 101638 131808 101694 131864
rect 135310 132896 135366 132952
rect 101822 132488 101878 132544
rect 135034 131828 135090 131864
rect 135034 131808 135036 131828
rect 135036 131808 135088 131828
rect 135088 131808 135090 131828
rect 135402 132352 135458 132408
rect 135034 131264 135090 131320
rect 101730 130720 101786 130776
rect 101362 129632 101418 129688
rect 101270 128952 101326 129008
rect 100994 128408 101050 128464
rect 101178 127864 101234 127920
rect 101086 127728 101142 127784
rect 100994 126232 101050 126288
rect 101822 130312 101878 130368
rect 135402 130604 135458 130640
rect 135402 130584 135404 130604
rect 135404 130584 135456 130604
rect 135456 130584 135458 130604
rect 135402 130040 135458 130096
rect 135310 129496 135366 129552
rect 135402 128816 135458 128872
rect 134666 128272 134722 128328
rect 135310 127748 135366 127784
rect 135310 127728 135312 127748
rect 135312 127728 135364 127748
rect 135364 127728 135366 127748
rect 135402 127184 135458 127240
rect 101270 126640 101326 126696
rect 135402 126504 135458 126560
rect 135218 125960 135274 126016
rect 100994 125552 101050 125608
rect 101270 125008 101326 125064
rect 101086 124736 101142 124792
rect 100994 123376 101050 123432
rect 101178 123784 101234 123840
rect 101086 122016 101142 122072
rect 100994 121472 101050 121528
rect 100994 120676 101050 120712
rect 100994 120656 100996 120676
rect 100996 120656 101048 120676
rect 101048 120656 101050 120676
rect 135402 125436 135458 125472
rect 135402 125416 135404 125436
rect 135404 125416 135456 125436
rect 135456 125416 135458 125436
rect 135402 124736 135458 124792
rect 134114 124192 134170 124248
rect 135034 123668 135090 123704
rect 135034 123648 135036 123668
rect 135036 123648 135088 123668
rect 135088 123648 135090 123668
rect 135218 122968 135274 123024
rect 101270 122560 101326 122616
rect 101178 120792 101234 120848
rect 135218 122424 135274 122480
rect 134850 121880 134906 121936
rect 134666 121336 134722 121392
rect 135402 120676 135458 120712
rect 135402 120656 135404 120676
rect 135404 120656 135456 120676
rect 135456 120656 135458 120676
rect 134298 120132 134354 120168
rect 134298 120112 134300 120132
rect 134300 120112 134352 120132
rect 134352 120112 134354 120132
rect 101086 119704 101142 119760
rect 135402 119588 135458 119624
rect 135402 119568 135404 119588
rect 135404 119568 135456 119588
rect 135456 119568 135458 119588
rect 100994 119316 101050 119352
rect 100994 119296 100996 119316
rect 100996 119296 101048 119316
rect 101048 119296 101050 119316
rect 134850 118888 134906 118944
rect 101086 118480 101142 118536
rect 100994 117936 101050 117992
rect 134482 118344 134538 118400
rect 134850 117800 134906 117856
rect 101178 117392 101234 117448
rect 101086 116712 101142 116768
rect 100994 116576 101050 116632
rect 134758 116576 134814 116632
rect 101086 115624 101142 115680
rect 100994 115216 101050 115272
rect 102006 114400 102062 114456
rect 101638 113856 101694 113912
rect 100994 112496 101050 112552
rect 99246 95496 99302 95552
rect 99154 94272 99210 94328
rect 101822 113720 101878 113776
rect 99522 98488 99578 98544
rect 106790 98488 106846 98544
rect 99430 96992 99486 97048
rect 106790 96176 106846 96232
rect 99338 93592 99394 93648
rect 99062 92368 99118 92424
rect 98970 91144 99026 91200
rect 106514 93864 106570 93920
rect 106790 91416 106846 91472
rect 99522 88696 99578 88752
rect 99522 85296 99578 85352
rect 99522 84636 99578 84672
rect 128502 89784 128558 89840
rect 106790 89104 106846 89160
rect 106790 86792 106846 86848
rect 99522 84616 99524 84636
rect 99524 84616 99576 84636
rect 99576 84616 99578 84636
rect 107802 84344 107858 84400
rect 99430 83936 99486 83992
rect 99522 82712 99578 82768
rect 106790 82068 106792 82088
rect 106792 82068 106844 82088
rect 106844 82068 106846 82088
rect 106790 82032 106846 82068
rect 99522 81488 99578 81544
rect 99522 79720 99578 79776
rect 106790 79720 106846 79776
rect 99522 77952 99578 78008
rect 106514 77408 106570 77464
rect 99522 76728 99578 76784
rect 106790 74996 106792 75016
rect 106792 74996 106844 75016
rect 106844 74996 106846 75016
rect 106790 74960 106846 74996
rect 99430 74280 99486 74336
rect 99522 73736 99578 73792
rect 99522 72512 99578 72568
rect 99522 71036 99578 71072
rect 99522 71016 99524 71036
rect 99524 71016 99576 71036
rect 99576 71016 99578 71036
rect 99522 69792 99578 69848
rect 98970 68296 99026 68352
rect 99062 67072 99118 67128
rect 99154 65848 99210 65904
rect 99246 64624 99302 64680
rect 99522 63400 99578 63456
rect 99338 62720 99394 62776
rect 99522 61496 99578 61552
rect 106790 72648 106846 72704
rect 106698 70336 106754 70392
rect 134942 117256 134998 117312
rect 134850 116032 134906 116088
rect 135034 115488 135090 115544
rect 135126 114808 135182 114864
rect 135310 114264 135366 114320
rect 135218 113176 135274 113232
rect 135402 113740 135458 113776
rect 135402 113720 135404 113740
rect 135404 113720 135456 113740
rect 135456 113720 135458 113740
rect 182782 155492 182838 155528
rect 182782 155472 182784 155492
rect 182784 155472 182836 155492
rect 182836 155472 182838 155492
rect 143590 138472 143646 138528
rect 143314 138200 143370 138256
rect 143130 136840 143186 136896
rect 143590 137112 143646 137168
rect 143498 136296 143554 136352
rect 143406 135752 143462 135808
rect 143314 135208 143370 135264
rect 143590 134256 143646 134312
rect 143222 133984 143278 134040
rect 142946 133304 143002 133360
rect 143590 132796 143592 132816
rect 143592 132796 143644 132816
rect 143644 132796 143646 132816
rect 143590 132760 143646 132796
rect 143222 132216 143278 132272
rect 143590 131400 143646 131456
rect 142486 130992 142542 131048
rect 143590 130212 143592 130232
rect 143592 130212 143644 130232
rect 143644 130212 143646 130232
rect 143590 130176 143646 130212
rect 143038 129904 143094 129960
rect 142762 128836 142818 128872
rect 142762 128816 142764 128836
rect 142764 128816 142816 128836
rect 142816 128816 142818 128836
rect 143590 128716 143592 128736
rect 143592 128716 143644 128736
rect 143644 128716 143646 128736
rect 143590 128680 143646 128716
rect 143130 128000 143186 128056
rect 142486 127356 142488 127376
rect 142488 127356 142540 127376
rect 142540 127356 142542 127376
rect 142486 127320 142542 127356
rect 143314 126912 143370 126968
rect 143590 125996 143592 126016
rect 143592 125996 143644 126016
rect 143644 125996 143646 126016
rect 143590 125960 143646 125996
rect 143498 125552 143554 125608
rect 142486 124364 142488 124384
rect 142488 124364 142540 124384
rect 142540 124364 142542 124384
rect 142486 124328 142542 124364
rect 143590 124600 143646 124656
rect 142762 123920 142818 123976
rect 143590 123276 143592 123296
rect 143592 123276 143644 123296
rect 143644 123276 143646 123296
rect 143590 123240 143646 123276
rect 143590 122424 143646 122480
rect 143038 121744 143094 121800
rect 142762 121472 142818 121528
rect 142946 120556 142948 120576
rect 142948 120556 143000 120576
rect 143000 120556 143002 120576
rect 142946 120520 143002 120556
rect 143590 120248 143646 120304
rect 143590 119196 143592 119216
rect 143592 119196 143644 119216
rect 143644 119196 143646 119216
rect 143590 119160 143646 119196
rect 143038 118888 143094 118944
rect 143314 118480 143370 118536
rect 142578 117664 142634 117720
rect 143222 117256 143278 117312
rect 142946 116340 142948 116360
rect 142948 116340 143000 116360
rect 143000 116340 143002 116360
rect 142946 116304 143002 116340
rect 143590 116032 143646 116088
rect 142762 115488 142818 115544
rect 183150 161592 183206 161648
rect 183242 160368 183298 160424
rect 183518 159144 183574 159200
rect 183334 157920 183390 157976
rect 183426 156696 183482 156752
rect 191982 168664 192038 168720
rect 191890 166760 191946 166816
rect 191338 164720 191394 164776
rect 211762 163768 211818 163824
rect 191522 162680 191578 162736
rect 191982 160776 192038 160832
rect 190050 158736 190106 158792
rect 189958 156696 190014 156752
rect 183610 154384 183666 154440
rect 191982 154792 192038 154848
rect 212682 157124 212738 157160
rect 212682 157104 212684 157124
rect 212684 157104 212736 157124
rect 212736 157104 212738 157124
rect 184990 140104 185046 140160
rect 177722 138492 177778 138528
rect 185082 139968 185138 140024
rect 185358 138880 185414 138936
rect 185266 138608 185322 138664
rect 177722 138472 177724 138492
rect 177724 138472 177776 138492
rect 177776 138472 177778 138492
rect 177630 138200 177686 138256
rect 185174 137792 185230 137848
rect 177722 136976 177778 137032
rect 177630 136840 177686 136896
rect 177722 136296 177778 136352
rect 177722 135480 177778 135536
rect 177630 135208 177686 135264
rect 185450 137248 185506 137304
rect 185174 136568 185230 136624
rect 177722 134292 177724 134312
rect 177724 134292 177776 134312
rect 177776 134292 177778 134312
rect 177722 134256 177778 134292
rect 185266 136024 185322 136080
rect 185358 135908 185414 135944
rect 185358 135888 185360 135908
rect 185360 135888 185412 135908
rect 185412 135888 185414 135908
rect 185174 134800 185230 134856
rect 185082 134392 185138 134448
rect 177722 133848 177778 133904
rect 177630 133440 177686 133496
rect 185174 133712 185230 133768
rect 185818 133032 185874 133088
rect 177722 132624 177778 132680
rect 185450 132488 185506 132544
rect 177630 132216 177686 132272
rect 185726 131944 185782 132000
rect 185542 131672 185598 131728
rect 177722 131264 177778 131320
rect 177630 130992 177686 131048
rect 185266 130720 185322 130776
rect 177722 130196 177778 130232
rect 177722 130176 177724 130196
rect 177724 130176 177776 130196
rect 177776 130176 177778 130196
rect 177630 129768 177686 129824
rect 185174 129632 185230 129688
rect 185358 130312 185414 130368
rect 177722 128680 177778 128736
rect 177630 128408 177686 128464
rect 185450 128952 185506 129008
rect 185174 128408 185230 128464
rect 177814 128000 177870 128056
rect 185358 127864 185414 127920
rect 185266 127592 185322 127648
rect 177170 127184 177226 127240
rect 177722 126912 177778 126968
rect 185174 126232 185230 126288
rect 177722 125960 177778 126016
rect 177630 125552 177686 125608
rect 177170 124192 177226 124248
rect 177722 124464 177778 124520
rect 220318 205384 220374 205440
rect 222342 179136 222398 179192
rect 217006 127320 217062 127376
rect 185450 126640 185506 126696
rect 185174 125552 185230 125608
rect 185450 124872 185506 124928
rect 185358 124736 185414 124792
rect 177630 123920 177686 123976
rect 185266 123376 185322 123432
rect 177722 122968 177778 123024
rect 177630 122696 177686 122752
rect 185818 123784 185874 123840
rect 185634 122560 185690 122616
rect 177722 121744 177778 121800
rect 177354 121472 177410 121528
rect 185358 121472 185414 121528
rect 185174 120792 185230 120848
rect 177722 120540 177778 120576
rect 177722 120520 177724 120540
rect 177724 120520 177776 120540
rect 177776 120520 177778 120540
rect 177630 120248 177686 120304
rect 177722 119060 177724 119080
rect 177724 119060 177776 119080
rect 177776 119060 177778 119080
rect 177722 119024 177778 119060
rect 177722 118752 177778 118808
rect 177630 118480 177686 118536
rect 177722 117528 177778 117584
rect 177170 117120 177226 117176
rect 177722 116340 177724 116360
rect 177724 116340 177776 116360
rect 177776 116340 177778 116360
rect 177722 116304 177778 116340
rect 177722 115896 177778 115952
rect 177078 115488 177134 115544
rect 185266 120692 185268 120712
rect 185268 120692 185320 120712
rect 185320 120692 185322 120712
rect 185266 120656 185322 120692
rect 185910 122152 185966 122208
rect 185266 119704 185322 119760
rect 185174 119316 185230 119352
rect 185174 119296 185176 119316
rect 185176 119296 185228 119316
rect 185228 119296 185230 119316
rect 185266 118480 185322 118536
rect 185174 117936 185230 117992
rect 222250 152888 222306 152944
rect 218386 135888 218442 135944
rect 218294 117800 218350 117856
rect 185358 117392 185414 117448
rect 185266 116712 185322 116768
rect 185174 116476 185176 116496
rect 185176 116476 185228 116496
rect 185228 116476 185230 116496
rect 185174 116440 185230 116476
rect 185266 115624 185322 115680
rect 185174 115216 185230 115272
rect 186002 114400 186058 114456
rect 185818 113856 185874 113912
rect 185174 112632 185230 112688
rect 183334 95496 183390 95552
rect 183242 94272 183298 94328
rect 186186 113720 186242 113776
rect 222342 126776 222398 126832
rect 183702 99168 183758 99224
rect 220962 100528 221018 100584
rect 191982 98760 192038 98816
rect 183610 97944 183666 98000
rect 183518 96720 183574 96776
rect 191982 94680 192038 94736
rect 183426 93048 183482 93104
rect 183150 91824 183206 91880
rect 183058 90600 183114 90656
rect 191154 92776 191210 92832
rect 190786 90736 190842 90792
rect 182874 89376 182930 89432
rect 183518 88152 183574 88208
rect 191706 88696 191762 88752
rect 183702 87064 183758 87120
rect 191614 86792 191670 86848
rect 183702 85840 183758 85896
rect 183702 84636 183758 84672
rect 191982 84752 192038 84808
rect 183702 84616 183704 84636
rect 183704 84616 183756 84636
rect 183756 84616 183758 84636
rect 182506 83392 182562 83448
rect 191982 82712 192038 82768
rect 183702 82168 183758 82224
rect 183242 80944 183298 81000
rect 191890 80808 191946 80864
rect 136874 80400 136930 80456
rect 183702 79720 183758 79776
rect 191982 78768 192038 78824
rect 183518 78496 183574 78552
rect 183058 77272 183114 77328
rect 209830 96856 209886 96912
rect 212314 96448 212370 96504
rect 212130 89784 212186 89840
rect 212038 83120 212094 83176
rect 209830 76864 209886 76920
rect 191982 76728 192038 76784
rect 183242 76048 183298 76104
rect 183702 74824 183758 74880
rect 183702 73756 183758 73792
rect 183702 73736 183704 73756
rect 183704 73736 183756 73756
rect 183756 73736 183758 73756
rect 191522 74688 191578 74744
rect 183702 72512 183758 72568
rect 183702 71288 183758 71344
rect 128502 69792 128558 69848
rect 106606 67888 106662 67944
rect 182874 70064 182930 70120
rect 183058 68840 183114 68896
rect 136874 66528 136930 66584
rect 137978 66528 138034 66584
rect 106514 65576 106570 65632
rect 106606 63264 106662 63320
rect 100258 59864 100314 59920
rect 79282 46808 79338 46864
rect 73394 46536 73450 46592
rect 76338 46400 76394 46456
rect 74866 46264 74922 46320
rect 77810 46128 77866 46184
rect 80754 46672 80810 46728
rect 85722 46264 85778 46320
rect 87102 46128 87158 46184
rect 58214 44360 58270 44416
rect 51222 44088 51278 44144
rect 107158 60952 107214 61008
rect 182690 60428 182746 60464
rect 182690 60408 182692 60428
rect 182692 60408 182744 60428
rect 182744 60408 182746 60428
rect 58306 43816 58362 43872
rect 58214 43172 58216 43192
rect 58216 43172 58268 43192
rect 58268 43172 58270 43192
rect 58214 43136 58270 43172
rect 58306 42592 58362 42648
rect 51130 42320 51186 42376
rect 51222 42048 51278 42104
rect 58214 42048 58270 42104
rect 58214 41368 58270 41424
rect 51130 41096 51186 41152
rect 51222 40824 51278 40880
rect 58306 40824 58362 40880
rect 58214 40144 58270 40200
rect 51130 39872 51186 39928
rect 58306 39600 58362 39656
rect 51222 39464 51278 39520
rect 58214 39092 58216 39112
rect 58216 39092 58268 39112
rect 58268 39092 58270 39112
rect 58214 39056 58270 39092
rect 51222 38784 51278 38840
rect 51130 38104 51186 38160
rect 58398 38376 58454 38432
rect 51222 37852 51278 37888
rect 51222 37832 51224 37852
rect 51224 37832 51276 37852
rect 51276 37832 51278 37852
rect 58306 37832 58362 37888
rect 51130 36880 51186 36936
rect 58398 37152 58454 37208
rect 51222 36608 51278 36664
rect 58214 36608 58270 36664
rect 58214 36064 58270 36120
rect 58306 35384 58362 35440
rect 51222 35248 51278 35304
rect 58214 34840 58270 34896
rect 51222 34160 51278 34216
rect 58306 34160 58362 34216
rect 51222 33752 51278 33808
rect 58214 33636 58270 33672
rect 58214 33616 58216 33636
rect 58216 33616 58268 33636
rect 58268 33616 58270 33636
rect 58214 33072 58270 33128
rect 51222 32412 51278 32448
rect 51222 32392 51224 32412
rect 51224 32392 51276 32412
rect 51276 32392 51278 32412
rect 58214 32392 58270 32448
rect 58214 31848 58270 31904
rect 51130 31576 51186 31632
rect 51222 31168 51278 31224
rect 58306 31168 58362 31224
rect 58214 30624 58270 30680
rect 51130 30352 51186 30408
rect 58306 30080 58362 30136
rect 51222 29808 51278 29864
rect 58214 29436 58216 29456
rect 58216 29436 58268 29456
rect 58268 29436 58270 29456
rect 58214 29400 58270 29436
rect 51130 29128 51186 29184
rect 58214 28856 58270 28912
rect 51222 28720 51278 28776
rect 51222 28332 51278 28368
rect 51222 28312 51224 28332
rect 51224 28312 51276 28332
rect 51276 28312 51278 28332
rect 58214 28176 58270 28232
rect 58214 27632 58270 27688
rect 51130 27360 51186 27416
rect 58306 27088 58362 27144
rect 51222 26952 51278 27008
rect 58214 26408 58270 26464
rect 58306 25864 58362 25920
rect 51222 25728 51278 25784
rect 51130 25456 51186 25512
rect 51130 24368 51186 24424
rect 59502 25184 59558 25240
rect 59410 24640 59466 24696
rect 51222 24096 51278 24152
rect 59318 24096 59374 24152
rect 58214 23416 58270 23472
rect 51222 22872 51278 22928
rect 58306 22872 58362 22928
rect 58214 22192 58270 22248
rect 51222 21920 51278 21976
rect 58306 21648 58362 21704
rect 92714 41232 92770 41288
rect 92714 40008 92770 40064
rect 92898 38240 92954 38296
rect 92898 35928 92954 35984
rect 92714 30488 92770 30544
rect 92714 28720 92770 28776
rect 92714 27496 92770 27552
rect 92898 23280 92954 23336
rect 58214 21104 58270 21160
rect 51038 20968 51094 21024
rect 61710 20968 61766 21024
rect 63182 20968 63238 21024
rect 64746 20968 64802 21024
rect 65114 20968 65170 21024
rect 62722 20832 62778 20888
rect 50854 20424 50910 20480
rect 50762 19744 50818 19800
rect 50578 19200 50634 19256
rect 66494 18248 66550 18304
rect 94002 44360 94058 44416
rect 93910 44224 93966 44280
rect 94002 43172 94004 43192
rect 94004 43172 94056 43192
rect 94056 43172 94058 43192
rect 94002 43136 94058 43172
rect 93910 42864 93966 42920
rect 94002 42456 94058 42512
rect 94002 41640 94058 41696
rect 94002 40144 94058 40200
rect 94002 39056 94058 39112
rect 93910 38648 93966 38704
rect 94002 37596 94004 37616
rect 94004 37596 94056 37616
rect 94056 37596 94058 37616
rect 94002 37560 94058 37596
rect 94002 37052 94004 37072
rect 94004 37052 94056 37072
rect 94056 37052 94058 37072
rect 94002 37016 94058 37052
rect 94002 36064 94058 36120
rect 94002 34840 94058 34896
rect 93450 34568 93506 34624
rect 93910 33616 93966 33672
rect 94002 33344 94058 33400
rect 93818 32936 93874 32992
rect 94002 31848 94058 31904
rect 93910 31712 93966 31768
rect 94002 30624 94058 30680
rect 94002 29400 94058 29456
rect 93910 29128 93966 29184
rect 94002 27904 94058 27960
rect 93910 26680 93966 26736
rect 94002 26308 94004 26328
rect 94004 26308 94056 26328
rect 94056 26308 94058 26328
rect 94002 26272 94058 26308
rect 94002 25220 94004 25240
rect 94004 25220 94056 25240
rect 94056 25220 94058 25240
rect 94002 25184 94058 25220
rect 93910 24912 93966 24968
rect 93818 24504 93874 24560
rect 94002 23688 94058 23744
rect 94002 22464 94058 22520
rect 93910 22056 93966 22112
rect 94002 21104 94058 21160
rect 101178 46128 101234 46184
rect 100994 45448 101050 45504
rect 101086 44768 101142 44824
rect 100994 43680 101050 43736
rect 100810 43408 100866 43464
rect 134298 45040 134354 45096
rect 101270 44904 101326 44960
rect 100994 42456 101050 42512
rect 100902 42048 100958 42104
rect 100810 40552 100866 40608
rect 100994 41232 101050 41288
rect 134758 46436 134760 46456
rect 134760 46436 134812 46456
rect 134812 46436 134814 46456
rect 134758 46400 134814 46436
rect 134850 45448 134906 45504
rect 134758 44768 134814 44824
rect 134758 43816 134814 43872
rect 134758 43408 134814 43464
rect 134758 42592 134814 42648
rect 134758 42048 134814 42104
rect 134666 41232 134722 41288
rect 134758 40960 134814 41016
rect 101086 40008 101142 40064
rect 134574 40008 134630 40064
rect 100994 39328 101050 39384
rect 134666 39464 134722 39520
rect 101086 38784 101142 38840
rect 134114 38784 134170 38840
rect 100994 38240 101050 38296
rect 100810 37832 100866 37888
rect 134298 38240 134354 38296
rect 134666 37988 134722 38024
rect 134666 37968 134668 37988
rect 134668 37968 134720 37988
rect 134720 37968 134722 37988
rect 100994 36880 101050 36936
rect 134666 36880 134722 36936
rect 100902 36472 100958 36528
rect 100718 35112 100774 35168
rect 134390 36628 134446 36664
rect 134390 36608 134392 36628
rect 134392 36608 134444 36628
rect 134444 36608 134446 36628
rect 134666 35928 134722 35984
rect 100994 35656 101050 35712
rect 134114 35248 134170 35304
rect 101086 34432 101142 34488
rect 134574 34432 134630 34488
rect 100994 33888 101050 33944
rect 100810 33752 100866 33808
rect 134666 34160 134722 34216
rect 134666 33772 134722 33808
rect 134666 33752 134668 33772
rect 134668 33752 134720 33772
rect 134720 33752 134722 33772
rect 100994 32664 101050 32720
rect 134298 32664 134354 32720
rect 100902 32256 100958 32312
rect 134390 32412 134446 32448
rect 134390 32392 134392 32412
rect 134392 32392 134444 32412
rect 134444 32392 134446 32412
rect 100810 30896 100866 30952
rect 134666 31576 134722 31632
rect 100994 31440 101050 31496
rect 134666 31032 134722 31088
rect 101086 30216 101142 30272
rect 100994 29672 101050 29728
rect 134206 29808 134262 29864
rect 101178 28992 101234 29048
rect 101086 28448 101142 28504
rect 100994 28196 101050 28232
rect 100994 28176 100996 28196
rect 100996 28176 101048 28196
rect 101048 28176 101050 28196
rect 100994 27224 101050 27280
rect 101178 26816 101234 26872
rect 101086 26000 101142 26056
rect 100994 25592 101050 25648
rect 101086 24776 101142 24832
rect 100994 24096 101050 24152
rect 100994 23552 101050 23608
rect 101086 22872 101142 22928
rect 101178 22600 101234 22656
rect 100994 22328 101050 22384
rect 101086 21920 101142 21976
rect 101546 19764 101602 19800
rect 101546 19744 101548 19764
rect 101548 19744 101600 19764
rect 101600 19744 101602 19764
rect 134758 30216 134814 30272
rect 134574 28992 134630 29048
rect 134758 28584 134814 28640
rect 134758 28212 134760 28232
rect 134760 28212 134812 28232
rect 134812 28212 134814 28232
rect 134758 28176 134814 28212
rect 134574 27224 134630 27280
rect 134758 26952 134814 27008
rect 134574 26000 134630 26056
rect 134758 25592 134814 25648
rect 134574 24776 134630 24832
rect 134758 24232 134814 24288
rect 134574 23552 134630 23608
rect 134758 23144 134814 23200
rect 134758 22756 134814 22792
rect 134758 22736 134760 22756
rect 134760 22736 134812 22756
rect 134812 22736 134814 22756
rect 134758 21104 134814 21160
rect 138070 46094 138126 46150
rect 138346 46128 138402 46184
rect 142394 44224 142450 44280
rect 142578 44360 142634 44416
rect 142486 43136 142542 43192
rect 154262 46128 154318 46184
rect 191982 72784 192038 72840
rect 190786 70744 190842 70800
rect 183150 67616 183206 67672
rect 183242 66392 183298 66448
rect 183334 65168 183390 65224
rect 183610 63944 183666 64000
rect 183426 62720 183482 62776
rect 190970 68704 191026 68760
rect 191338 66800 191394 66856
rect 191522 64760 191578 64816
rect 189958 62720 190014 62776
rect 183702 61516 183758 61552
rect 183702 61496 183704 61516
rect 183704 61496 183756 61516
rect 183756 61496 183758 61516
rect 191982 60816 192038 60872
rect 164750 46808 164806 46864
rect 161898 46672 161954 46728
rect 158954 46536 159010 46592
rect 157574 46264 157630 46320
rect 160334 46400 160390 46456
rect 163278 46264 163334 46320
rect 222342 74280 222398 74336
rect 212682 69812 212738 69848
rect 212682 69792 212684 69812
rect 212684 69792 212736 69812
rect 212736 69792 212738 69812
rect 169902 46264 169958 46320
rect 171098 46128 171154 46184
rect 172938 44632 172994 44688
rect 142670 43000 142726 43056
rect 143130 42456 143186 42512
rect 143498 41912 143554 41968
rect 142762 41232 142818 41288
rect 135310 22464 135366 22520
rect 135126 21920 135182 21976
rect 143682 40144 143738 40200
rect 142394 40008 142450 40064
rect 142486 39076 142542 39112
rect 142486 39056 142488 39076
rect 142488 39056 142540 39076
rect 142540 39056 142542 39076
rect 142394 38920 142450 38976
rect 142578 38240 142634 38296
rect 142394 37696 142450 37752
rect 142486 37016 142542 37072
rect 142578 36336 142634 36392
rect 142394 35928 142450 35984
rect 142394 34704 142450 34760
rect 142578 34840 142634 34896
rect 142486 33616 142542 33672
rect 142394 33344 142450 33400
rect 142394 32936 142450 32992
rect 142486 32156 142488 32176
rect 142488 32156 142540 32176
rect 142540 32156 142542 32176
rect 142486 32120 142542 32156
rect 142394 31712 142450 31768
rect 142394 30624 142450 30680
rect 142394 30524 142396 30544
rect 142396 30524 142448 30544
rect 142448 30524 142450 30544
rect 142394 30488 142450 30524
rect 143590 29400 143646 29456
rect 142394 29264 142450 29320
rect 142486 28720 142542 28776
rect 142394 27904 142450 27960
rect 142394 27496 142450 27552
rect 142486 26716 142488 26736
rect 142488 26716 142540 26736
rect 142540 26716 142542 26736
rect 142486 26680 142542 26716
rect 142394 26272 142450 26328
rect 142394 25048 142450 25104
rect 142578 25184 142634 25240
rect 142486 24504 142542 24560
rect 142394 23824 142450 23880
rect 142486 23280 142542 23336
rect 142394 22464 142450 22520
rect 142486 22056 142542 22112
rect 135034 20696 135090 20752
rect 134942 19744 134998 19800
rect 101822 19472 101878 19528
rect 134482 19472 134538 19528
rect 143682 21104 143738 21160
rect 146258 20968 146314 21024
rect 147730 20968 147786 21024
rect 148742 20968 148798 21024
rect 150858 20968 150914 21024
rect 145706 20832 145762 20888
rect 149754 18248 149810 18304
rect 129054 17024 129110 17080
rect 177262 39600 177318 39656
rect 177446 38376 177502 38432
rect 177354 37832 177410 37888
rect 177446 37152 177502 37208
rect 177354 35384 177410 35440
rect 176986 31848 177042 31904
rect 177446 30624 177502 30680
rect 177170 30080 177226 30136
rect 177262 27088 177318 27144
rect 177446 26408 177502 26464
rect 177354 24096 177410 24152
rect 185818 46128 185874 46184
rect 185174 45448 185230 45504
rect 177722 44360 177778 44416
rect 185450 44904 185506 44960
rect 177722 43852 177724 43872
rect 177724 43852 177776 43872
rect 177776 43852 177778 43872
rect 177722 43816 177778 43852
rect 185174 43680 185230 43736
rect 184990 43408 185046 43464
rect 177722 43136 177778 43192
rect 177630 42592 177686 42648
rect 177722 42048 177778 42104
rect 185542 44768 185598 44824
rect 185174 42456 185230 42512
rect 185082 42048 185138 42104
rect 177722 41368 177778 41424
rect 177630 40824 177686 40880
rect 184990 40552 185046 40608
rect 177722 40144 177778 40200
rect 177722 39056 177778 39112
rect 185174 41232 185230 41288
rect 185266 40008 185322 40064
rect 185174 39328 185230 39384
rect 185266 38784 185322 38840
rect 185174 38104 185230 38160
rect 184990 37832 185046 37888
rect 177722 36608 177778 36664
rect 185174 36880 185230 36936
rect 185082 36472 185138 36528
rect 177722 36064 177778 36120
rect 184898 35248 184954 35304
rect 177722 34840 177778 34896
rect 177630 34160 177686 34216
rect 177630 33616 177686 33672
rect 177722 33072 177778 33128
rect 185450 35656 185506 35712
rect 185266 34432 185322 34488
rect 185174 33888 185230 33944
rect 184990 33752 185046 33808
rect 177814 32392 177870 32448
rect 222250 48032 222306 48088
rect 215718 33344 215774 33400
rect 185174 32664 185230 32720
rect 185082 32256 185138 32312
rect 177722 31168 177778 31224
rect 184990 30896 185046 30952
rect 177722 29400 177778 29456
rect 185174 31440 185230 31496
rect 185266 30216 185322 30272
rect 185174 29672 185230 29728
rect 185358 28992 185414 29048
rect 177814 28856 177870 28912
rect 185266 28448 185322 28504
rect 177630 28176 177686 28232
rect 185174 28196 185230 28232
rect 185174 28176 185176 28196
rect 185176 28176 185228 28196
rect 185228 28176 185230 28196
rect 177722 27632 177778 27688
rect 185174 27224 185230 27280
rect 185358 26816 185414 26872
rect 177722 25864 177778 25920
rect 185542 26000 185598 26056
rect 185450 25592 185506 25648
rect 177722 25184 177778 25240
rect 185266 24776 185322 24832
rect 177630 24640 177686 24696
rect 177722 23416 177778 23472
rect 177538 22872 177594 22928
rect 177630 22192 177686 22248
rect 177722 21648 177778 21704
rect 177722 21104 177778 21160
rect 185174 24096 185230 24152
rect 185266 23552 185322 23608
rect 185174 22872 185230 22928
rect 185266 22600 185322 22656
rect 185174 22328 185230 22384
rect 185174 19764 185230 19800
rect 185174 19744 185176 19764
rect 185176 19744 185228 19764
rect 185228 19744 185230 19764
rect 185266 19472 185322 19528
rect 212498 18420 212500 18440
rect 212500 18420 212552 18440
rect 212552 18420 212554 18440
rect 212498 18384 212554 18420
<< metal3 >>
rect 189166 236524 189172 236588
rect 189236 236586 189242 236588
rect 194921 236586 194987 236589
rect 189236 236584 194987 236586
rect 189236 236528 194926 236584
rect 194982 236528 194987 236584
rect 189236 236526 194987 236528
rect 189236 236524 189242 236526
rect 194921 236523 194987 236526
rect 79553 235226 79619 235229
rect 88518 235226 88524 235228
rect 79553 235224 88524 235226
rect 79553 235168 79558 235224
rect 79614 235168 88524 235224
rect 79553 235166 88524 235168
rect 79553 235163 79619 235166
rect 88518 235164 88524 235166
rect 88588 235164 88594 235228
rect 50665 234546 50731 234549
rect 134753 234546 134819 234549
rect 47892 234544 50731 234546
rect 47892 234488 50670 234544
rect 50726 234488 50731 234544
rect 47892 234486 50731 234488
rect 131796 234544 134819 234546
rect 131796 234488 134758 234544
rect 134814 234488 134819 234544
rect 131796 234486 134819 234488
rect 50665 234483 50731 234486
rect 134753 234483 134819 234486
rect 185997 234546 186063 234549
rect 185997 234544 187916 234546
rect 185997 234488 186002 234544
rect 186058 234488 187916 234544
rect 185997 234486 187916 234488
rect 185997 234483 186063 234486
rect 101633 234138 101699 234141
rect 101633 234136 103674 234138
rect 101633 234080 101638 234136
rect 101694 234080 103674 234136
rect 101633 234078 103674 234080
rect 101633 234075 101699 234078
rect 49929 234002 49995 234005
rect 47892 234000 49995 234002
rect 47892 233944 49934 234000
rect 49990 233944 49995 234000
rect 47892 233942 49995 233944
rect 49929 233939 49995 233942
rect 103614 233934 103674 234078
rect 135397 234002 135463 234005
rect 131796 234000 135463 234002
rect 131796 233944 135402 234000
rect 135458 233944 135463 234000
rect 131796 233942 135463 233944
rect 135397 233939 135463 233942
rect 185077 234002 185143 234005
rect 185077 234000 187916 234002
rect 185077 233944 185082 234000
rect 185138 233944 187916 234000
rect 185077 233942 187916 233944
rect 185077 233939 185143 233942
rect 103614 233874 104012 233934
rect 50573 233458 50639 233461
rect 134293 233458 134359 233461
rect 47892 233456 50639 233458
rect 47892 233400 50578 233456
rect 50634 233400 50639 233456
rect 47892 233398 50639 233400
rect 131796 233456 134359 233458
rect 131796 233400 134298 233456
rect 134354 233400 134359 233456
rect 131796 233398 134359 233400
rect 50573 233395 50639 233398
rect 134293 233395 134359 233398
rect 185169 233458 185235 233461
rect 185169 233456 187916 233458
rect 185169 233400 185174 233456
rect 185230 233400 187916 233456
rect 185169 233398 187916 233400
rect 185169 233395 185235 233398
rect 100989 233186 101055 233189
rect 103982 233186 104042 233360
rect 100989 233184 104042 233186
rect 100989 233128 100994 233184
rect 101050 233128 104042 233184
rect 100989 233126 104042 233128
rect 100989 233123 101055 233126
rect 58117 233050 58183 233053
rect 142297 233050 142363 233053
rect 177165 233050 177231 233053
rect 58117 233048 60986 233050
rect 58117 232992 58122 233048
rect 58178 232992 60986 233048
rect 58117 232990 60986 232992
rect 58117 232987 58183 232990
rect 9896 232914 10376 232944
rect 12761 232914 12827 232917
rect 51217 232914 51283 232917
rect 9896 232912 12827 232914
rect 9896 232856 12766 232912
rect 12822 232856 12827 232912
rect 9896 232854 12827 232856
rect 47892 232912 51283 232914
rect 47892 232856 51222 232912
rect 51278 232856 51283 232912
rect 47892 232854 51283 232856
rect 9896 232824 10376 232854
rect 12761 232851 12827 232854
rect 51217 232851 51283 232854
rect 60926 232476 60986 232990
rect 142297 233048 145074 233050
rect 142297 232992 142302 233048
rect 142358 232992 145074 233048
rect 142297 232990 145074 232992
rect 142297 232987 142363 232990
rect 135397 232914 135463 232917
rect 131796 232912 135463 232914
rect 131796 232856 135402 232912
rect 135458 232856 135463 232912
rect 131796 232854 135463 232856
rect 135397 232851 135463 232854
rect 100989 232642 101055 232645
rect 103982 232642 104042 232816
rect 100989 232640 104042 232642
rect 100989 232584 100994 232640
rect 101050 232584 104042 232640
rect 100989 232582 104042 232584
rect 100989 232579 101055 232582
rect 92709 232506 92775 232509
rect 90764 232504 92775 232506
rect 90764 232448 92714 232504
rect 92770 232448 92775 232504
rect 145014 232476 145074 232990
rect 174822 233048 177231 233050
rect 174822 232992 177170 233048
rect 177226 232992 177231 233048
rect 174822 232990 177231 232992
rect 163549 232642 163615 232645
rect 171134 232642 171140 232644
rect 163549 232640 171140 232642
rect 163549 232584 163554 232640
rect 163610 232584 171140 232640
rect 163549 232582 171140 232584
rect 163549 232579 163615 232582
rect 171134 232580 171140 232582
rect 171204 232580 171210 232644
rect 174822 232476 174882 232990
rect 177165 232987 177231 232990
rect 185261 232914 185327 232917
rect 185261 232912 187916 232914
rect 185261 232856 185266 232912
rect 185322 232856 187916 232912
rect 185261 232854 187916 232856
rect 185261 232851 185327 232854
rect 90764 232446 92775 232448
rect 92709 232443 92775 232446
rect 51125 232234 51191 232237
rect 47892 232232 51191 232234
rect 47892 232176 51130 232232
rect 51186 232176 51191 232232
rect 47892 232174 51191 232176
rect 51125 232171 51191 232174
rect 100989 232098 101055 232101
rect 103982 232098 104042 232272
rect 135397 232234 135463 232237
rect 177717 232234 177783 232237
rect 131796 232232 135463 232234
rect 131796 232176 135402 232232
rect 135458 232176 135463 232232
rect 131796 232174 135463 232176
rect 135397 232171 135463 232174
rect 174822 232232 177783 232234
rect 174822 232176 177722 232232
rect 177778 232176 177783 232232
rect 174822 232174 177783 232176
rect 100989 232096 104042 232098
rect 100989 232040 100994 232096
rect 101050 232040 104042 232096
rect 100989 232038 104042 232040
rect 100989 232035 101055 232038
rect 58117 231962 58183 231965
rect 93997 231962 94063 231965
rect 58117 231960 60956 231962
rect 58117 231904 58122 231960
rect 58178 231904 60956 231960
rect 58117 231902 60956 231904
rect 90764 231960 94063 231962
rect 90764 231904 94002 231960
rect 94058 231904 94063 231960
rect 90764 231902 94063 231904
rect 58117 231899 58183 231902
rect 93997 231899 94063 231902
rect 142297 231962 142363 231965
rect 142297 231960 145044 231962
rect 142297 231904 142302 231960
rect 142358 231904 145044 231960
rect 174822 231932 174882 232174
rect 177717 232171 177783 232174
rect 185261 232234 185327 232237
rect 185261 232232 187916 232234
rect 185261 232176 185266 232232
rect 185322 232176 187916 232232
rect 185261 232174 187916 232176
rect 185261 232171 185327 232174
rect 142297 231902 145044 231904
rect 142297 231899 142363 231902
rect 51217 231690 51283 231693
rect 47892 231688 51283 231690
rect 47892 231632 51222 231688
rect 51278 231632 51283 231688
rect 47892 231630 51283 231632
rect 51217 231627 51283 231630
rect 100989 231554 101055 231557
rect 103982 231554 104042 231728
rect 134845 231690 134911 231693
rect 131796 231688 134911 231690
rect 131796 231632 134850 231688
rect 134906 231632 134911 231688
rect 131796 231630 134911 231632
rect 134845 231627 134911 231630
rect 185169 231690 185235 231693
rect 222337 231690 222403 231693
rect 225416 231690 225896 231720
rect 185169 231688 187916 231690
rect 185169 231632 185174 231688
rect 185230 231632 187916 231688
rect 185169 231630 187916 231632
rect 222337 231688 225896 231690
rect 222337 231632 222342 231688
rect 222398 231632 225896 231688
rect 222337 231630 225896 231632
rect 185169 231627 185235 231630
rect 222337 231627 222403 231630
rect 225416 231600 225896 231630
rect 177717 231554 177783 231557
rect 100989 231552 104042 231554
rect 100989 231496 100994 231552
rect 101050 231496 104042 231552
rect 100989 231494 104042 231496
rect 174822 231552 177783 231554
rect 174822 231496 177722 231552
rect 177778 231496 177783 231552
rect 174822 231494 177783 231496
rect 100989 231491 101055 231494
rect 58025 231282 58091 231285
rect 92709 231282 92775 231285
rect 58025 231280 60956 231282
rect 58025 231224 58030 231280
rect 58086 231224 60956 231280
rect 58025 231222 60956 231224
rect 90764 231280 92775 231282
rect 90764 231224 92714 231280
rect 92770 231224 92775 231280
rect 90764 231222 92775 231224
rect 58025 231219 58091 231222
rect 92709 231219 92775 231222
rect 142205 231282 142271 231285
rect 142205 231280 145044 231282
rect 142205 231224 142210 231280
rect 142266 231224 145044 231280
rect 174822 231252 174882 231494
rect 177717 231491 177783 231494
rect 142205 231222 145044 231224
rect 142205 231219 142271 231222
rect 103614 231154 104012 231214
rect 51217 231146 51283 231149
rect 47892 231144 51283 231146
rect 47892 231088 51222 231144
rect 51278 231088 51283 231144
rect 47892 231086 51283 231088
rect 51217 231083 51283 231086
rect 101081 231146 101147 231149
rect 103614 231146 103674 231154
rect 135305 231146 135371 231149
rect 101081 231144 103674 231146
rect 101081 231088 101086 231144
rect 101142 231088 103674 231144
rect 101081 231086 103674 231088
rect 131796 231144 135371 231146
rect 131796 231088 135310 231144
rect 135366 231088 135371 231144
rect 131796 231086 135371 231088
rect 101081 231083 101147 231086
rect 135305 231083 135371 231086
rect 185353 231146 185419 231149
rect 185353 231144 187916 231146
rect 185353 231088 185358 231144
rect 185414 231088 187916 231144
rect 185353 231086 187916 231088
rect 185353 231083 185419 231086
rect 178177 230874 178243 230877
rect 174822 230872 178243 230874
rect 174822 230816 178182 230872
rect 178238 230816 178243 230872
rect 174822 230814 178243 230816
rect 58209 230738 58275 230741
rect 92709 230738 92775 230741
rect 58209 230736 60956 230738
rect 58209 230680 58214 230736
rect 58270 230680 60956 230736
rect 58209 230678 60956 230680
rect 90764 230736 92775 230738
rect 90764 230680 92714 230736
rect 92770 230680 92775 230736
rect 90764 230678 92775 230680
rect 58209 230675 58275 230678
rect 92709 230675 92775 230678
rect 143677 230738 143743 230741
rect 143677 230736 145044 230738
rect 143677 230680 143682 230736
rect 143738 230680 145044 230736
rect 174822 230708 174882 230814
rect 178177 230811 178243 230814
rect 215713 230738 215779 230741
rect 215670 230736 215779 230738
rect 143677 230678 145044 230680
rect 215670 230680 215718 230736
rect 215774 230680 215779 230736
rect 143677 230675 143743 230678
rect 215670 230675 215779 230680
rect 51125 230602 51191 230605
rect 47892 230600 51191 230602
rect 47892 230544 51130 230600
rect 51186 230544 51191 230600
rect 47892 230542 51191 230544
rect 51125 230539 51191 230542
rect 58301 230194 58367 230197
rect 94089 230194 94155 230197
rect 58301 230192 60956 230194
rect 58301 230136 58306 230192
rect 58362 230136 60956 230192
rect 58301 230134 60956 230136
rect 90764 230192 94155 230194
rect 90764 230136 94094 230192
rect 94150 230136 94155 230192
rect 90764 230134 94155 230136
rect 58301 230131 58367 230134
rect 94089 230131 94155 230134
rect 101081 230194 101147 230197
rect 103982 230194 104042 230640
rect 135397 230602 135463 230605
rect 131796 230600 135463 230602
rect 131796 230544 135402 230600
rect 135458 230544 135463 230600
rect 131796 230542 135463 230544
rect 135397 230539 135463 230542
rect 185261 230602 185327 230605
rect 185261 230600 187916 230602
rect 185261 230544 185266 230600
rect 185322 230544 187916 230600
rect 185261 230542 187916 230544
rect 185261 230539 185327 230542
rect 177717 230466 177783 230469
rect 174822 230464 177783 230466
rect 174822 230408 177722 230464
rect 177778 230408 177783 230464
rect 174822 230406 177783 230408
rect 101081 230192 104042 230194
rect 101081 230136 101086 230192
rect 101142 230136 104042 230192
rect 101081 230134 104042 230136
rect 142941 230194 143007 230197
rect 142941 230192 145044 230194
rect 142941 230136 142946 230192
rect 143002 230136 145044 230192
rect 174822 230164 174882 230406
rect 177717 230403 177783 230406
rect 215670 230164 215730 230675
rect 142941 230134 145044 230136
rect 101081 230131 101147 230134
rect 142941 230131 143007 230134
rect 51217 230058 51283 230061
rect 135305 230058 135371 230061
rect 47892 230056 51283 230058
rect 47892 230000 51222 230056
rect 51278 230000 51283 230056
rect 47892 229998 51283 230000
rect 131796 230056 135371 230058
rect 131796 230000 135310 230056
rect 135366 230000 135371 230056
rect 131796 229998 135371 230000
rect 51217 229995 51283 229998
rect 135305 229995 135371 229998
rect 185169 230058 185235 230061
rect 185169 230056 187916 230058
rect 185169 230000 185174 230056
rect 185230 230000 187916 230056
rect 185169 229998 187916 230000
rect 185169 229995 185235 229998
rect 100989 229786 101055 229789
rect 103982 229786 104042 229960
rect 100989 229784 104042 229786
rect 100989 229728 100994 229784
rect 101050 229728 104042 229784
rect 100989 229726 104042 229728
rect 100989 229723 101055 229726
rect 58209 229514 58275 229517
rect 92709 229514 92775 229517
rect 58209 229512 60956 229514
rect 58209 229456 58214 229512
rect 58270 229456 60956 229512
rect 58209 229454 60956 229456
rect 90764 229512 92775 229514
rect 90764 229456 92714 229512
rect 92770 229456 92775 229512
rect 90764 229454 92775 229456
rect 58209 229451 58275 229454
rect 92709 229451 92775 229454
rect 143677 229514 143743 229517
rect 143677 229512 145044 229514
rect 143677 229456 143682 229512
rect 143738 229456 145044 229512
rect 143677 229454 145044 229456
rect 143677 229451 143743 229454
rect 51125 229378 51191 229381
rect 47892 229376 51191 229378
rect 47892 229320 51130 229376
rect 51186 229320 51191 229376
rect 47892 229318 51191 229320
rect 51125 229315 51191 229318
rect 100989 229242 101055 229245
rect 103982 229242 104042 229416
rect 135397 229378 135463 229381
rect 131796 229376 135463 229378
rect 131796 229320 135402 229376
rect 135458 229320 135463 229376
rect 131796 229318 135463 229320
rect 174822 229378 174882 229484
rect 177717 229378 177783 229381
rect 174822 229376 177783 229378
rect 174822 229320 177722 229376
rect 177778 229320 177783 229376
rect 174822 229318 177783 229320
rect 135397 229315 135463 229318
rect 177717 229315 177783 229318
rect 185629 229378 185695 229381
rect 185629 229376 187916 229378
rect 185629 229320 185634 229376
rect 185690 229320 187916 229376
rect 185629 229318 187916 229320
rect 185629 229315 185695 229318
rect 177625 229242 177691 229245
rect 100989 229240 104042 229242
rect 100989 229184 100994 229240
rect 101050 229184 104042 229240
rect 100989 229182 104042 229184
rect 174822 229240 177691 229242
rect 174822 229184 177630 229240
rect 177686 229184 177691 229240
rect 174822 229182 177691 229184
rect 100989 229179 101055 229182
rect 58209 228970 58275 228973
rect 93169 228970 93235 228973
rect 58209 228968 60956 228970
rect 58209 228912 58214 228968
rect 58270 228912 60956 228968
rect 58209 228910 60956 228912
rect 90764 228968 93235 228970
rect 90764 228912 93174 228968
rect 93230 228912 93235 228968
rect 90764 228910 93235 228912
rect 58209 228907 58275 228910
rect 93169 228907 93235 228910
rect 143585 228970 143651 228973
rect 143585 228968 145044 228970
rect 143585 228912 143590 228968
rect 143646 228912 145044 228968
rect 174822 228940 174882 229182
rect 177625 229179 177691 229182
rect 143585 228910 145044 228912
rect 143585 228907 143651 228910
rect 50757 228834 50823 228837
rect 47892 228832 50823 228834
rect 47892 228776 50762 228832
rect 50818 228776 50823 228832
rect 47892 228774 50823 228776
rect 50757 228771 50823 228774
rect 101081 228698 101147 228701
rect 103982 228698 104042 228872
rect 135305 228834 135371 228837
rect 131796 228832 135371 228834
rect 131796 228776 135310 228832
rect 135366 228776 135371 228832
rect 131796 228774 135371 228776
rect 135305 228771 135371 228774
rect 185905 228834 185971 228837
rect 185905 228832 187916 228834
rect 185905 228776 185910 228832
rect 185966 228776 187916 228832
rect 185905 228774 187916 228776
rect 185905 228771 185971 228774
rect 177809 228698 177875 228701
rect 101081 228696 104042 228698
rect 101081 228640 101086 228696
rect 101142 228640 104042 228696
rect 101081 228638 104042 228640
rect 174822 228696 177875 228698
rect 174822 228640 177814 228696
rect 177870 228640 177875 228696
rect 174822 228638 177875 228640
rect 101081 228635 101147 228638
rect 103614 228298 104012 228358
rect 51217 228290 51283 228293
rect 47892 228288 51283 228290
rect 47892 228232 51222 228288
rect 51278 228232 51283 228288
rect 47892 228230 51283 228232
rect 51217 228227 51283 228230
rect 58301 228290 58367 228293
rect 92709 228290 92775 228293
rect 58301 228288 60956 228290
rect 58301 228232 58306 228288
rect 58362 228232 60956 228288
rect 58301 228230 60956 228232
rect 90764 228288 92775 228290
rect 90764 228232 92714 228288
rect 92770 228232 92775 228288
rect 90764 228230 92775 228232
rect 58301 228227 58367 228230
rect 92709 228227 92775 228230
rect 100989 228290 101055 228293
rect 103614 228290 103674 228298
rect 135397 228290 135463 228293
rect 100989 228288 103674 228290
rect 100989 228232 100994 228288
rect 101050 228232 103674 228288
rect 100989 228230 103674 228232
rect 131796 228288 135463 228290
rect 131796 228232 135402 228288
rect 135458 228232 135463 228288
rect 131796 228230 135463 228232
rect 100989 228227 101055 228230
rect 135397 228227 135463 228230
rect 143493 228290 143559 228293
rect 143493 228288 145044 228290
rect 143493 228232 143498 228288
rect 143554 228232 145044 228288
rect 174822 228260 174882 228638
rect 177809 228635 177875 228638
rect 185169 228290 185235 228293
rect 185169 228288 187916 228290
rect 143493 228230 145044 228232
rect 185169 228232 185174 228288
rect 185230 228232 187916 228288
rect 185169 228230 187916 228232
rect 143493 228227 143559 228230
rect 185169 228227 185235 228230
rect 177717 228018 177783 228021
rect 174822 228016 177783 228018
rect 174822 227960 177722 228016
rect 177778 227960 177783 228016
rect 174822 227958 177783 227960
rect 50941 227746 51007 227749
rect 47892 227744 51007 227746
rect 47892 227688 50946 227744
rect 51002 227688 51007 227744
rect 47892 227686 51007 227688
rect 50941 227683 51007 227686
rect 58209 227746 58275 227749
rect 93169 227746 93235 227749
rect 58209 227744 60956 227746
rect 58209 227688 58214 227744
rect 58270 227688 60956 227744
rect 58209 227686 60956 227688
rect 90764 227744 93235 227746
rect 90764 227688 93174 227744
rect 93230 227688 93235 227744
rect 90764 227686 93235 227688
rect 58209 227683 58275 227686
rect 93169 227683 93235 227686
rect 101081 227474 101147 227477
rect 103982 227474 104042 227784
rect 135397 227746 135463 227749
rect 131796 227744 135463 227746
rect 131796 227688 135402 227744
rect 135458 227688 135463 227744
rect 131796 227686 135463 227688
rect 135397 227683 135463 227686
rect 143677 227746 143743 227749
rect 143677 227744 145044 227746
rect 143677 227688 143682 227744
rect 143738 227688 145044 227744
rect 174822 227716 174882 227958
rect 177717 227955 177783 227958
rect 185169 227746 185235 227749
rect 185169 227744 187916 227746
rect 143677 227686 145044 227688
rect 185169 227688 185174 227744
rect 185230 227688 187916 227744
rect 185169 227686 187916 227688
rect 143677 227683 143743 227686
rect 185169 227683 185235 227686
rect 177625 227474 177691 227477
rect 101081 227472 104042 227474
rect 101081 227416 101086 227472
rect 101142 227416 104042 227472
rect 101081 227414 104042 227416
rect 174822 227472 177691 227474
rect 174822 227416 177630 227472
rect 177686 227416 177691 227472
rect 174822 227414 177691 227416
rect 101081 227411 101147 227414
rect 51217 227202 51283 227205
rect 47892 227200 51283 227202
rect 47892 227144 51222 227200
rect 51278 227144 51283 227200
rect 47892 227142 51283 227144
rect 51217 227139 51283 227142
rect 58301 227202 58367 227205
rect 92709 227202 92775 227205
rect 58301 227200 60956 227202
rect 58301 227144 58306 227200
rect 58362 227144 60956 227200
rect 58301 227142 60956 227144
rect 90764 227200 92775 227202
rect 90764 227144 92714 227200
rect 92770 227144 92775 227200
rect 90764 227142 92775 227144
rect 58301 227139 58367 227142
rect 92709 227139 92775 227142
rect 100989 227066 101055 227069
rect 103982 227066 104042 227240
rect 135305 227202 135371 227205
rect 131796 227200 135371 227202
rect 131796 227144 135310 227200
rect 135366 227144 135371 227200
rect 131796 227142 135371 227144
rect 135305 227139 135371 227142
rect 143309 227202 143375 227205
rect 143309 227200 145044 227202
rect 143309 227144 143314 227200
rect 143370 227144 145044 227200
rect 174822 227172 174882 227414
rect 177625 227411 177691 227414
rect 185261 227202 185327 227205
rect 185261 227200 187916 227202
rect 143309 227142 145044 227144
rect 185261 227144 185266 227200
rect 185322 227144 187916 227200
rect 185261 227142 187916 227144
rect 143309 227139 143375 227142
rect 185261 227139 185327 227142
rect 100989 227064 104042 227066
rect 100989 227008 100994 227064
rect 101050 227008 104042 227064
rect 100989 227006 104042 227008
rect 100989 227003 101055 227006
rect 50757 226522 50823 226525
rect 47892 226520 50823 226522
rect 47892 226464 50762 226520
rect 50818 226464 50823 226520
rect 47892 226462 50823 226464
rect 50757 226459 50823 226462
rect 58209 226522 58275 226525
rect 92709 226522 92775 226525
rect 58209 226520 60956 226522
rect 58209 226464 58214 226520
rect 58270 226464 60956 226520
rect 58209 226462 60956 226464
rect 90764 226520 92775 226522
rect 90764 226464 92714 226520
rect 92770 226464 92775 226520
rect 90764 226462 92775 226464
rect 58209 226459 58275 226462
rect 92709 226459 92775 226462
rect 101081 226386 101147 226389
rect 103982 226386 104042 226696
rect 177717 226658 177783 226661
rect 174822 226656 177783 226658
rect 174822 226600 177722 226656
rect 177778 226600 177783 226656
rect 174822 226598 177783 226600
rect 135213 226522 135279 226525
rect 131796 226520 135279 226522
rect 131796 226464 135218 226520
rect 135274 226464 135279 226520
rect 131796 226462 135279 226464
rect 135213 226459 135279 226462
rect 143677 226522 143743 226525
rect 143677 226520 145044 226522
rect 143677 226464 143682 226520
rect 143738 226464 145044 226520
rect 174822 226492 174882 226598
rect 177717 226595 177783 226598
rect 185169 226522 185235 226525
rect 185169 226520 187916 226522
rect 143677 226462 145044 226464
rect 185169 226464 185174 226520
rect 185230 226464 187916 226520
rect 185169 226462 187916 226464
rect 143677 226459 143743 226462
rect 185169 226459 185235 226462
rect 101081 226384 104042 226386
rect 101081 226328 101086 226384
rect 101142 226328 104042 226384
rect 101081 226326 104042 226328
rect 101081 226323 101147 226326
rect 177625 226250 177691 226253
rect 174822 226248 177691 226250
rect 174822 226192 177630 226248
rect 177686 226192 177691 226248
rect 174822 226190 177691 226192
rect 50481 225978 50547 225981
rect 47892 225976 50547 225978
rect 47892 225920 50486 225976
rect 50542 225920 50547 225976
rect 47892 225918 50547 225920
rect 50481 225915 50547 225918
rect 58301 225978 58367 225981
rect 93629 225978 93695 225981
rect 58301 225976 60956 225978
rect 58301 225920 58306 225976
rect 58362 225920 60956 225976
rect 58301 225918 60956 225920
rect 90764 225976 93695 225978
rect 90764 225920 93634 225976
rect 93690 225920 93695 225976
rect 90764 225918 93695 225920
rect 58301 225915 58367 225918
rect 93629 225915 93695 225918
rect 101173 225706 101239 225709
rect 103982 225706 104042 226152
rect 134569 225978 134635 225981
rect 131796 225976 134635 225978
rect 131796 225920 134574 225976
rect 134630 225920 134635 225976
rect 131796 225918 134635 225920
rect 134569 225915 134635 225918
rect 143309 225978 143375 225981
rect 143309 225976 145044 225978
rect 143309 225920 143314 225976
rect 143370 225920 145044 225976
rect 174822 225948 174882 226190
rect 177625 226187 177691 226190
rect 185261 225978 185327 225981
rect 185261 225976 187916 225978
rect 143309 225918 145044 225920
rect 185261 225920 185266 225976
rect 185322 225920 187916 225976
rect 185261 225918 187916 225920
rect 143309 225915 143375 225918
rect 185261 225915 185327 225918
rect 101173 225704 104042 225706
rect 101173 225648 101178 225704
rect 101234 225648 104042 225704
rect 101173 225646 104042 225648
rect 101173 225643 101239 225646
rect 100989 225570 101055 225573
rect 100989 225568 104012 225570
rect 100989 225512 100994 225568
rect 101050 225512 104012 225568
rect 100989 225510 104012 225512
rect 100989 225507 101055 225510
rect 51125 225434 51191 225437
rect 135305 225434 135371 225437
rect 177717 225434 177783 225437
rect 47892 225432 51191 225434
rect 47892 225376 51130 225432
rect 51186 225376 51191 225432
rect 47892 225374 51191 225376
rect 131796 225432 135371 225434
rect 131796 225376 135310 225432
rect 135366 225376 135371 225432
rect 131796 225374 135371 225376
rect 51125 225371 51191 225374
rect 135305 225371 135371 225374
rect 174822 225432 177783 225434
rect 174822 225376 177722 225432
rect 177778 225376 177783 225432
rect 174822 225374 177783 225376
rect 58209 225298 58275 225301
rect 92801 225298 92867 225301
rect 58209 225296 60956 225298
rect 58209 225240 58214 225296
rect 58270 225240 60956 225296
rect 58209 225238 60956 225240
rect 90764 225296 92867 225298
rect 90764 225240 92806 225296
rect 92862 225240 92867 225296
rect 90764 225238 92867 225240
rect 58209 225235 58275 225238
rect 92801 225235 92867 225238
rect 143677 225298 143743 225301
rect 143677 225296 145044 225298
rect 143677 225240 143682 225296
rect 143738 225240 145044 225296
rect 174822 225268 174882 225374
rect 177717 225371 177783 225374
rect 185353 225434 185419 225437
rect 185353 225432 187916 225434
rect 185353 225376 185358 225432
rect 185414 225376 187916 225432
rect 185353 225374 187916 225376
rect 185353 225371 185419 225374
rect 143677 225238 145044 225240
rect 143677 225235 143743 225238
rect 177625 225026 177691 225029
rect 174822 225024 177691 225026
rect 174822 224968 177630 225024
rect 177686 224968 177691 225024
rect 174822 224966 177691 224968
rect 51217 224890 51283 224893
rect 47892 224888 51283 224890
rect 47892 224832 51222 224888
rect 51278 224832 51283 224888
rect 47892 224830 51283 224832
rect 51217 224827 51283 224830
rect 58301 224754 58367 224757
rect 92709 224754 92775 224757
rect 58301 224752 60956 224754
rect 58301 224696 58306 224752
rect 58362 224696 60956 224752
rect 58301 224694 60956 224696
rect 90764 224752 92775 224754
rect 90764 224696 92714 224752
rect 92770 224696 92775 224752
rect 90764 224694 92775 224696
rect 58301 224691 58367 224694
rect 92709 224691 92775 224694
rect 101081 224618 101147 224621
rect 103982 224618 104042 224928
rect 135397 224890 135463 224893
rect 131796 224888 135463 224890
rect 131796 224832 135402 224888
rect 135458 224832 135463 224888
rect 131796 224830 135463 224832
rect 135397 224827 135463 224830
rect 143585 224754 143651 224757
rect 143585 224752 145044 224754
rect 143585 224696 143590 224752
rect 143646 224696 145044 224752
rect 174822 224724 174882 224966
rect 177625 224963 177691 224966
rect 185169 224890 185235 224893
rect 185169 224888 187916 224890
rect 185169 224832 185174 224888
rect 185230 224832 187916 224888
rect 185169 224830 187916 224832
rect 185169 224827 185235 224830
rect 143585 224694 145044 224696
rect 143585 224691 143651 224694
rect 101081 224616 104042 224618
rect 101081 224560 101086 224616
rect 101142 224560 104042 224616
rect 101081 224558 104042 224560
rect 101081 224555 101147 224558
rect 177809 224482 177875 224485
rect 174822 224480 177875 224482
rect 174822 224424 177814 224480
rect 177870 224424 177875 224480
rect 174822 224422 177875 224424
rect 51033 224346 51099 224349
rect 47892 224344 51099 224346
rect 47892 224288 51038 224344
rect 51094 224288 51099 224344
rect 47892 224286 51099 224288
rect 51033 224283 51099 224286
rect 58393 224210 58459 224213
rect 92893 224210 92959 224213
rect 58393 224208 60956 224210
rect 58393 224152 58398 224208
rect 58454 224152 60956 224208
rect 58393 224150 60956 224152
rect 90764 224208 92959 224210
rect 90764 224152 92898 224208
rect 92954 224152 92959 224208
rect 90764 224150 92959 224152
rect 58393 224147 58459 224150
rect 92893 224147 92959 224150
rect 100989 224210 101055 224213
rect 103982 224210 104042 224384
rect 135213 224346 135279 224349
rect 131796 224344 135279 224346
rect 131796 224288 135218 224344
rect 135274 224288 135279 224344
rect 131796 224286 135279 224288
rect 135213 224283 135279 224286
rect 100989 224208 104042 224210
rect 100989 224152 100994 224208
rect 101050 224152 104042 224208
rect 100989 224150 104042 224152
rect 143493 224210 143559 224213
rect 143493 224208 145044 224210
rect 143493 224152 143498 224208
rect 143554 224152 145044 224208
rect 174822 224180 174882 224422
rect 177809 224419 177875 224422
rect 185261 224346 185327 224349
rect 185261 224344 187916 224346
rect 185261 224288 185266 224344
rect 185322 224288 187916 224344
rect 185261 224286 187916 224288
rect 185261 224283 185327 224286
rect 143493 224150 145044 224152
rect 100989 224147 101055 224150
rect 143493 224147 143559 224150
rect 50941 223666 51007 223669
rect 47892 223664 51007 223666
rect 47892 223608 50946 223664
rect 51002 223608 51007 223664
rect 47892 223606 51007 223608
rect 50941 223603 51007 223606
rect 58209 223530 58275 223533
rect 93721 223530 93787 223533
rect 58209 223528 60956 223530
rect 58209 223472 58214 223528
rect 58270 223472 60956 223528
rect 58209 223470 60956 223472
rect 90764 223528 93787 223530
rect 90764 223472 93726 223528
rect 93782 223472 93787 223528
rect 90764 223470 93787 223472
rect 58209 223467 58275 223470
rect 93721 223467 93787 223470
rect 101449 223530 101515 223533
rect 103982 223530 104042 223840
rect 177717 223802 177783 223805
rect 174822 223800 177783 223802
rect 174822 223744 177722 223800
rect 177778 223744 177783 223800
rect 174822 223742 177783 223744
rect 135397 223666 135463 223669
rect 131796 223664 135463 223666
rect 131796 223608 135402 223664
rect 135458 223608 135463 223664
rect 131796 223606 135463 223608
rect 135397 223603 135463 223606
rect 101449 223528 104042 223530
rect 101449 223472 101454 223528
rect 101510 223472 104042 223528
rect 101449 223470 104042 223472
rect 143677 223530 143743 223533
rect 143677 223528 145044 223530
rect 143677 223472 143682 223528
rect 143738 223472 145044 223528
rect 174822 223500 174882 223742
rect 177717 223739 177783 223742
rect 185169 223666 185235 223669
rect 185169 223664 187916 223666
rect 185169 223608 185174 223664
rect 185230 223608 187916 223664
rect 185169 223606 187916 223608
rect 185169 223603 185235 223606
rect 143677 223470 145044 223472
rect 101449 223467 101515 223470
rect 143677 223467 143743 223470
rect 51217 223122 51283 223125
rect 47892 223120 51283 223122
rect 47892 223064 51222 223120
rect 51278 223064 51283 223120
rect 47892 223062 51283 223064
rect 51217 223059 51283 223062
rect 101541 223122 101607 223125
rect 103982 223122 104042 223296
rect 177349 223258 177415 223261
rect 174822 223256 177415 223258
rect 174822 223200 177354 223256
rect 177410 223200 177415 223256
rect 174822 223198 177415 223200
rect 135305 223122 135371 223125
rect 101541 223120 104042 223122
rect 101541 223064 101546 223120
rect 101602 223064 104042 223120
rect 101541 223062 104042 223064
rect 131796 223120 135371 223122
rect 131796 223064 135310 223120
rect 135366 223064 135371 223120
rect 131796 223062 135371 223064
rect 101541 223059 101607 223062
rect 135305 223059 135371 223062
rect 58301 222986 58367 222989
rect 93905 222986 93971 222989
rect 58301 222984 60956 222986
rect 58301 222928 58306 222984
rect 58362 222928 60956 222984
rect 58301 222926 60956 222928
rect 90764 222984 93971 222986
rect 90764 222928 93910 222984
rect 93966 222928 93971 222984
rect 90764 222926 93971 222928
rect 58301 222923 58367 222926
rect 93905 222923 93971 222926
rect 143309 222986 143375 222989
rect 143309 222984 145044 222986
rect 143309 222928 143314 222984
rect 143370 222928 145044 222984
rect 174822 222956 174882 223198
rect 177349 223195 177415 223198
rect 185445 223122 185511 223125
rect 185445 223120 187916 223122
rect 185445 223064 185450 223120
rect 185506 223064 187916 223120
rect 185445 223062 187916 223064
rect 185445 223059 185511 223062
rect 143309 222926 145044 222928
rect 143309 222923 143375 222926
rect 101265 222850 101331 222853
rect 101265 222848 104012 222850
rect 101265 222792 101270 222848
rect 101326 222792 104012 222848
rect 101265 222790 104012 222792
rect 101265 222787 101331 222790
rect 51125 222578 51191 222581
rect 134845 222578 134911 222581
rect 47892 222576 51191 222578
rect 47892 222520 51130 222576
rect 51186 222520 51191 222576
rect 47892 222518 51191 222520
rect 131796 222576 134911 222578
rect 131796 222520 134850 222576
rect 134906 222520 134911 222576
rect 131796 222518 134911 222520
rect 51125 222515 51191 222518
rect 134845 222515 134911 222518
rect 185261 222578 185327 222581
rect 185261 222576 187916 222578
rect 185261 222520 185266 222576
rect 185322 222520 187916 222576
rect 185261 222518 187916 222520
rect 185261 222515 185327 222518
rect 177717 222442 177783 222445
rect 174822 222440 177783 222442
rect 174822 222384 177722 222440
rect 177778 222384 177783 222440
rect 174822 222382 177783 222384
rect 58209 222306 58275 222309
rect 92709 222306 92775 222309
rect 58209 222304 60956 222306
rect 58209 222248 58214 222304
rect 58270 222248 60956 222304
rect 58209 222246 60956 222248
rect 90764 222304 92775 222306
rect 90764 222248 92714 222304
rect 92770 222248 92775 222304
rect 90764 222246 92775 222248
rect 58209 222243 58275 222246
rect 92709 222243 92775 222246
rect 143677 222306 143743 222309
rect 143677 222304 145044 222306
rect 143677 222248 143682 222304
rect 143738 222248 145044 222304
rect 174822 222276 174882 222382
rect 177717 222379 177783 222382
rect 143677 222246 145044 222248
rect 143677 222243 143743 222246
rect 51217 222034 51283 222037
rect 47892 222032 51283 222034
rect 47892 221976 51222 222032
rect 51278 221976 51283 222032
rect 47892 221974 51283 221976
rect 51217 221971 51283 221974
rect 101541 221898 101607 221901
rect 103982 221898 104042 222208
rect 134477 222034 134543 222037
rect 177625 222034 177691 222037
rect 131796 222032 134543 222034
rect 131796 221976 134482 222032
rect 134538 221976 134543 222032
rect 131796 221974 134543 221976
rect 134477 221971 134543 221974
rect 174822 222032 177691 222034
rect 174822 221976 177630 222032
rect 177686 221976 177691 222032
rect 174822 221974 177691 221976
rect 101541 221896 104042 221898
rect 101541 221840 101546 221896
rect 101602 221840 104042 221896
rect 101541 221838 104042 221840
rect 101541 221835 101607 221838
rect 58301 221762 58367 221765
rect 92985 221762 93051 221765
rect 58301 221760 60956 221762
rect 58301 221704 58306 221760
rect 58362 221704 60956 221760
rect 58301 221702 60956 221704
rect 90764 221760 93051 221762
rect 90764 221704 92990 221760
rect 93046 221704 93051 221760
rect 90764 221702 93051 221704
rect 58301 221699 58367 221702
rect 92985 221699 93051 221702
rect 143309 221762 143375 221765
rect 143309 221760 145044 221762
rect 143309 221704 143314 221760
rect 143370 221704 145044 221760
rect 174822 221732 174882 221974
rect 177625 221971 177691 221974
rect 185169 222034 185235 222037
rect 185169 222032 187916 222034
rect 185169 221976 185174 222032
rect 185230 221976 187916 222032
rect 185169 221974 187916 221976
rect 185169 221971 185235 221974
rect 143309 221702 145044 221704
rect 143309 221699 143375 221702
rect 51217 221490 51283 221493
rect 47892 221488 51283 221490
rect 47892 221432 51222 221488
rect 51278 221432 51283 221488
rect 47892 221430 51283 221432
rect 51217 221427 51283 221430
rect 101725 221490 101791 221493
rect 103982 221490 104042 221664
rect 135305 221490 135371 221493
rect 101725 221488 104042 221490
rect 101725 221432 101730 221488
rect 101786 221432 104042 221488
rect 101725 221430 104042 221432
rect 131796 221488 135371 221490
rect 131796 221432 135310 221488
rect 135366 221432 135371 221488
rect 131796 221430 135371 221432
rect 101725 221427 101791 221430
rect 135305 221427 135371 221430
rect 185353 221490 185419 221493
rect 185353 221488 187916 221490
rect 185353 221432 185358 221488
rect 185414 221432 187916 221488
rect 185353 221430 187916 221432
rect 185353 221427 185419 221430
rect 58209 221218 58275 221221
rect 92709 221218 92775 221221
rect 58209 221216 60956 221218
rect 58209 221160 58214 221216
rect 58270 221160 60956 221216
rect 58209 221158 60956 221160
rect 90764 221216 92775 221218
rect 90764 221160 92714 221216
rect 92770 221160 92775 221216
rect 90764 221158 92775 221160
rect 58209 221155 58275 221158
rect 92709 221155 92775 221158
rect 143677 221218 143743 221221
rect 143677 221216 145044 221218
rect 143677 221160 143682 221216
rect 143738 221160 145044 221216
rect 143677 221158 145044 221160
rect 143677 221155 143743 221158
rect 18097 220946 18163 220949
rect 18097 220944 19924 220946
rect 18097 220888 18102 220944
rect 18158 220888 19924 220944
rect 18097 220886 19924 220888
rect 18097 220883 18163 220886
rect 50941 220810 51007 220813
rect 47892 220808 51007 220810
rect 47892 220752 50946 220808
rect 51002 220752 51007 220808
rect 47892 220750 51007 220752
rect 50941 220747 51007 220750
rect 101725 220674 101791 220677
rect 103982 220674 104042 221120
rect 174822 221082 174882 221188
rect 177717 221082 177783 221085
rect 174822 221080 177783 221082
rect 174822 221024 177722 221080
rect 177778 221024 177783 221080
rect 174822 221022 177783 221024
rect 177717 221019 177783 221022
rect 177625 220946 177691 220949
rect 174822 220944 177691 220946
rect 174822 220888 177630 220944
rect 177686 220888 177691 220944
rect 174822 220886 177691 220888
rect 135397 220810 135463 220813
rect 131796 220808 135463 220810
rect 131796 220752 135402 220808
rect 135458 220752 135463 220808
rect 131796 220750 135463 220752
rect 135397 220747 135463 220750
rect 101725 220672 104042 220674
rect 101725 220616 101730 220672
rect 101786 220616 104042 220672
rect 101725 220614 104042 220616
rect 101725 220611 101791 220614
rect 58209 220538 58275 220541
rect 93721 220538 93787 220541
rect 58209 220536 60956 220538
rect 58209 220480 58214 220536
rect 58270 220480 60956 220536
rect 58209 220478 60956 220480
rect 90764 220536 93787 220538
rect 90764 220480 93726 220536
rect 93782 220480 93787 220536
rect 90764 220478 93787 220480
rect 58209 220475 58275 220478
rect 93721 220475 93787 220478
rect 143585 220538 143651 220541
rect 143585 220536 145044 220538
rect 143585 220480 143590 220536
rect 143646 220480 145044 220536
rect 174822 220508 174882 220886
rect 177625 220883 177691 220886
rect 185169 220810 185235 220813
rect 220313 220810 220379 220813
rect 185169 220808 187916 220810
rect 185169 220752 185174 220808
rect 185230 220752 187916 220808
rect 185169 220750 187916 220752
rect 215884 220808 220379 220810
rect 215884 220752 220318 220808
rect 220374 220752 220379 220808
rect 215884 220750 220379 220752
rect 185169 220747 185235 220750
rect 220313 220747 220379 220750
rect 143585 220478 145044 220480
rect 143585 220475 143651 220478
rect 50205 220266 50271 220269
rect 47892 220264 50271 220266
rect 47892 220208 50210 220264
rect 50266 220208 50271 220264
rect 47892 220206 50271 220208
rect 50205 220203 50271 220206
rect 101817 220266 101883 220269
rect 103982 220266 104042 220440
rect 135305 220266 135371 220269
rect 177809 220266 177875 220269
rect 101817 220264 104042 220266
rect 101817 220208 101822 220264
rect 101878 220208 104042 220264
rect 101817 220206 104042 220208
rect 131796 220264 135371 220266
rect 131796 220208 135310 220264
rect 135366 220208 135371 220264
rect 131796 220206 135371 220208
rect 101817 220203 101883 220206
rect 135305 220203 135371 220206
rect 174822 220264 177875 220266
rect 174822 220208 177814 220264
rect 177870 220208 177875 220264
rect 174822 220206 177875 220208
rect 58301 219994 58367 219997
rect 93169 219994 93235 219997
rect 58301 219992 60956 219994
rect 58301 219936 58306 219992
rect 58362 219936 60956 219992
rect 58301 219934 60956 219936
rect 90764 219992 93235 219994
rect 90764 219936 93174 219992
rect 93230 219936 93235 219992
rect 90764 219934 93235 219936
rect 58301 219931 58367 219934
rect 93169 219931 93235 219934
rect 101909 219994 101975 219997
rect 143677 219994 143743 219997
rect 101909 219992 104012 219994
rect 101909 219936 101914 219992
rect 101970 219936 104012 219992
rect 101909 219934 104012 219936
rect 143677 219992 145044 219994
rect 143677 219936 143682 219992
rect 143738 219936 145044 219992
rect 174822 219964 174882 220206
rect 177809 220203 177875 220206
rect 185537 220266 185603 220269
rect 185537 220264 187916 220266
rect 185537 220208 185542 220264
rect 185598 220208 187916 220264
rect 185537 220206 187916 220208
rect 185537 220203 185603 220206
rect 143677 219934 145044 219936
rect 101909 219931 101975 219934
rect 143677 219931 143743 219934
rect 50849 219722 50915 219725
rect 135397 219722 135463 219725
rect 47892 219720 50915 219722
rect 47892 219664 50854 219720
rect 50910 219664 50915 219720
rect 47892 219662 50915 219664
rect 131796 219720 135463 219722
rect 131796 219664 135402 219720
rect 135458 219664 135463 219720
rect 131796 219662 135463 219664
rect 50849 219659 50915 219662
rect 135397 219659 135463 219662
rect 185721 219722 185787 219725
rect 185721 219720 187916 219722
rect 185721 219664 185726 219720
rect 185782 219664 187916 219720
rect 185721 219662 187916 219664
rect 185721 219659 185787 219662
rect 177717 219586 177783 219589
rect 174822 219584 177783 219586
rect 174822 219528 177722 219584
rect 177778 219528 177783 219584
rect 174822 219526 177783 219528
rect 58209 219314 58275 219317
rect 92801 219314 92867 219317
rect 58209 219312 60956 219314
rect 58209 219256 58214 219312
rect 58270 219256 60956 219312
rect 58209 219254 60956 219256
rect 90764 219312 92867 219314
rect 90764 219256 92806 219312
rect 92862 219256 92867 219312
rect 90764 219254 92867 219256
rect 58209 219251 58275 219254
rect 92801 219251 92867 219254
rect 50205 219178 50271 219181
rect 47892 219176 50271 219178
rect 47892 219120 50210 219176
rect 50266 219120 50271 219176
rect 47892 219118 50271 219120
rect 50205 219115 50271 219118
rect 101725 219042 101791 219045
rect 103982 219042 104042 219352
rect 143677 219314 143743 219317
rect 143677 219312 145044 219314
rect 143677 219256 143682 219312
rect 143738 219256 145044 219312
rect 174822 219284 174882 219526
rect 177717 219523 177783 219526
rect 143677 219254 145044 219256
rect 143677 219251 143743 219254
rect 135029 219178 135095 219181
rect 131796 219176 135095 219178
rect 131796 219120 135034 219176
rect 135090 219120 135095 219176
rect 131796 219118 135095 219120
rect 135029 219115 135095 219118
rect 185629 219178 185695 219181
rect 185629 219176 187916 219178
rect 185629 219120 185634 219176
rect 185690 219120 187916 219176
rect 185629 219118 187916 219120
rect 185629 219115 185695 219118
rect 177625 219042 177691 219045
rect 101725 219040 104042 219042
rect 101725 218984 101730 219040
rect 101786 218984 104042 219040
rect 101725 218982 104042 218984
rect 174822 219040 177691 219042
rect 174822 218984 177630 219040
rect 177686 218984 177691 219040
rect 174822 218982 177691 218984
rect 101725 218979 101791 218982
rect 58301 218770 58367 218773
rect 92709 218770 92775 218773
rect 58301 218768 60956 218770
rect 58301 218712 58306 218768
rect 58362 218712 60956 218768
rect 58301 218710 60956 218712
rect 90764 218768 92775 218770
rect 90764 218712 92714 218768
rect 92770 218712 92775 218768
rect 90764 218710 92775 218712
rect 58301 218707 58367 218710
rect 92709 218707 92775 218710
rect 51217 218634 51283 218637
rect 47892 218632 51283 218634
rect 47892 218576 51222 218632
rect 51278 218576 51283 218632
rect 47892 218574 51283 218576
rect 51217 218571 51283 218574
rect 102001 218634 102067 218637
rect 103982 218634 104042 218808
rect 143125 218770 143191 218773
rect 143125 218768 145044 218770
rect 143125 218712 143130 218768
rect 143186 218712 145044 218768
rect 174822 218740 174882 218982
rect 177625 218979 177691 218982
rect 143125 218710 145044 218712
rect 143125 218707 143191 218710
rect 135305 218634 135371 218637
rect 102001 218632 104042 218634
rect 102001 218576 102006 218632
rect 102062 218576 104042 218632
rect 102001 218574 104042 218576
rect 131796 218632 135371 218634
rect 131796 218576 135310 218632
rect 135366 218576 135371 218632
rect 131796 218574 135371 218576
rect 102001 218571 102067 218574
rect 135305 218571 135371 218574
rect 185905 218634 185971 218637
rect 185905 218632 187916 218634
rect 185905 218576 185910 218632
rect 185966 218576 187916 218632
rect 185905 218574 187916 218576
rect 185905 218571 185971 218574
rect 177717 218362 177783 218365
rect 174822 218360 177783 218362
rect 174822 218304 177722 218360
rect 177778 218304 177783 218360
rect 174822 218302 177783 218304
rect 58209 218226 58275 218229
rect 92801 218226 92867 218229
rect 58209 218224 60956 218226
rect 58209 218168 58214 218224
rect 58270 218168 60956 218224
rect 58209 218166 60956 218168
rect 90764 218224 92867 218226
rect 90764 218168 92806 218224
rect 92862 218168 92867 218224
rect 90764 218166 92867 218168
rect 58209 218163 58275 218166
rect 92801 218163 92867 218166
rect 51217 217954 51283 217957
rect 47892 217952 51283 217954
rect 47892 217896 51222 217952
rect 51278 217896 51283 217952
rect 47892 217894 51283 217896
rect 51217 217891 51283 217894
rect 101909 217954 101975 217957
rect 103982 217954 104042 218264
rect 143677 218226 143743 218229
rect 143677 218224 145044 218226
rect 143677 218168 143682 218224
rect 143738 218168 145044 218224
rect 174822 218196 174882 218302
rect 177717 218299 177783 218302
rect 143677 218166 145044 218168
rect 143677 218163 143743 218166
rect 135397 217954 135463 217957
rect 177625 217954 177691 217957
rect 101909 217952 104042 217954
rect 101909 217896 101914 217952
rect 101970 217896 104042 217952
rect 101909 217894 104042 217896
rect 131796 217952 135463 217954
rect 131796 217896 135402 217952
rect 135458 217896 135463 217952
rect 131796 217894 135463 217896
rect 101909 217891 101975 217894
rect 135397 217891 135463 217894
rect 174822 217952 177691 217954
rect 174822 217896 177630 217952
rect 177686 217896 177691 217952
rect 174822 217894 177691 217896
rect 58209 217546 58275 217549
rect 93721 217546 93787 217549
rect 58209 217544 60956 217546
rect 58209 217488 58214 217544
rect 58270 217488 60956 217544
rect 58209 217486 60956 217488
rect 90764 217544 93787 217546
rect 90764 217488 93726 217544
rect 93782 217488 93787 217544
rect 90764 217486 93787 217488
rect 58209 217483 58275 217486
rect 93721 217483 93787 217486
rect 101817 217546 101883 217549
rect 103982 217546 104042 217720
rect 101817 217544 104042 217546
rect 101817 217488 101822 217544
rect 101878 217488 104042 217544
rect 101817 217486 104042 217488
rect 143493 217546 143559 217549
rect 143493 217544 145044 217546
rect 143493 217488 143498 217544
rect 143554 217488 145044 217544
rect 174822 217516 174882 217894
rect 177625 217891 177691 217894
rect 185721 217954 185787 217957
rect 185721 217952 187916 217954
rect 185721 217896 185726 217952
rect 185782 217896 187916 217952
rect 185721 217894 187916 217896
rect 185721 217891 185787 217894
rect 143493 217486 145044 217488
rect 101817 217483 101883 217486
rect 143493 217483 143559 217486
rect 51217 217410 51283 217413
rect 135397 217410 135463 217413
rect 47892 217408 51283 217410
rect 47892 217352 51222 217408
rect 51278 217352 51283 217408
rect 47892 217350 51283 217352
rect 131796 217408 135463 217410
rect 131796 217352 135402 217408
rect 135458 217352 135463 217408
rect 131796 217350 135463 217352
rect 51217 217347 51283 217350
rect 135397 217347 135463 217350
rect 185537 217410 185603 217413
rect 185537 217408 187916 217410
rect 185537 217352 185542 217408
rect 185598 217352 187916 217408
rect 185537 217350 187916 217352
rect 185537 217347 185603 217350
rect 101725 217274 101791 217277
rect 101725 217272 104012 217274
rect 101725 217216 101730 217272
rect 101786 217216 104012 217272
rect 101725 217214 104012 217216
rect 101725 217211 101791 217214
rect 177717 217138 177783 217141
rect 174822 217136 177783 217138
rect 174822 217080 177722 217136
rect 177778 217080 177783 217136
rect 174822 217078 177783 217080
rect 58209 217002 58275 217005
rect 93905 217002 93971 217005
rect 58209 217000 60956 217002
rect 58209 216944 58214 217000
rect 58270 216944 60956 217000
rect 58209 216942 60956 216944
rect 90764 217000 93971 217002
rect 90764 216944 93910 217000
rect 93966 216944 93971 217000
rect 90764 216942 93971 216944
rect 58209 216939 58275 216942
rect 93905 216939 93971 216942
rect 143677 217002 143743 217005
rect 143677 217000 145044 217002
rect 143677 216944 143682 217000
rect 143738 216944 145044 217000
rect 174822 216972 174882 217078
rect 177717 217075 177783 217078
rect 143677 216942 145044 216944
rect 143677 216939 143743 216942
rect 51125 216866 51191 216869
rect 135397 216866 135463 216869
rect 47892 216864 51191 216866
rect 47892 216808 51130 216864
rect 51186 216808 51191 216864
rect 47892 216806 51191 216808
rect 131796 216864 135463 216866
rect 131796 216808 135402 216864
rect 135458 216808 135463 216864
rect 131796 216806 135463 216808
rect 51125 216803 51191 216806
rect 135397 216803 135463 216806
rect 185905 216866 185971 216869
rect 185905 216864 187916 216866
rect 185905 216808 185910 216864
rect 185966 216808 187916 216864
rect 185905 216806 187916 216808
rect 185905 216803 185971 216806
rect 177625 216730 177691 216733
rect 174822 216728 177691 216730
rect 174822 216672 177630 216728
rect 177686 216672 177691 216728
rect 174822 216670 177691 216672
rect 51217 216322 51283 216325
rect 47892 216320 51283 216322
rect 47892 216264 51222 216320
rect 51278 216264 51283 216320
rect 47892 216262 51283 216264
rect 51217 216259 51283 216262
rect 58301 216322 58367 216325
rect 92709 216322 92775 216325
rect 58301 216320 60956 216322
rect 58301 216264 58306 216320
rect 58362 216264 60956 216320
rect 58301 216262 60956 216264
rect 90764 216320 92775 216322
rect 90764 216264 92714 216320
rect 92770 216264 92775 216320
rect 90764 216262 92775 216264
rect 58301 216259 58367 216262
rect 92709 216259 92775 216262
rect 101817 216186 101883 216189
rect 103982 216186 104042 216632
rect 135489 216322 135555 216325
rect 131796 216320 135555 216322
rect 131796 216264 135494 216320
rect 135550 216264 135555 216320
rect 131796 216262 135555 216264
rect 135489 216259 135555 216262
rect 143125 216322 143191 216325
rect 143125 216320 145044 216322
rect 143125 216264 143130 216320
rect 143186 216264 145044 216320
rect 174822 216292 174882 216670
rect 177625 216667 177691 216670
rect 185721 216322 185787 216325
rect 185721 216320 187916 216322
rect 143125 216262 145044 216264
rect 185721 216264 185726 216320
rect 185782 216264 187916 216320
rect 185721 216262 187916 216264
rect 143125 216259 143191 216262
rect 185721 216259 185787 216262
rect 101817 216184 104042 216186
rect 101817 216128 101822 216184
rect 101878 216128 104042 216184
rect 101817 216126 104042 216128
rect 101817 216123 101883 216126
rect 101725 216050 101791 216053
rect 101725 216048 104012 216050
rect 101725 215992 101730 216048
rect 101786 215992 104012 216048
rect 101725 215990 104012 215992
rect 101725 215987 101791 215990
rect 51217 215778 51283 215781
rect 47892 215776 51283 215778
rect 47892 215720 51222 215776
rect 51278 215720 51283 215776
rect 47892 215718 51283 215720
rect 51217 215715 51283 215718
rect 58209 215778 58275 215781
rect 92709 215778 92775 215781
rect 135397 215778 135463 215781
rect 58209 215776 60956 215778
rect 58209 215720 58214 215776
rect 58270 215720 60956 215776
rect 58209 215718 60956 215720
rect 90764 215776 92775 215778
rect 90764 215720 92714 215776
rect 92770 215720 92775 215776
rect 90764 215718 92775 215720
rect 131796 215776 135463 215778
rect 131796 215720 135402 215776
rect 135458 215720 135463 215776
rect 131796 215718 135463 215720
rect 58209 215715 58275 215718
rect 92709 215715 92775 215718
rect 135397 215715 135463 215718
rect 143125 215778 143191 215781
rect 185629 215778 185695 215781
rect 143125 215776 145044 215778
rect 143125 215720 143130 215776
rect 143186 215720 145044 215776
rect 185629 215776 187916 215778
rect 143125 215718 145044 215720
rect 143125 215715 143191 215718
rect 174822 215642 174882 215748
rect 185629 215720 185634 215776
rect 185690 215720 187916 215776
rect 185629 215718 187916 215720
rect 185629 215715 185695 215718
rect 177717 215642 177783 215645
rect 174822 215640 177783 215642
rect 174822 215584 177722 215640
rect 177778 215584 177783 215640
rect 174822 215582 177783 215584
rect 177717 215579 177783 215582
rect 58301 215234 58367 215237
rect 92801 215234 92867 215237
rect 58301 215232 60956 215234
rect 58301 215176 58306 215232
rect 58362 215176 60956 215232
rect 58301 215174 60956 215176
rect 90764 215232 92867 215234
rect 90764 215176 92806 215232
rect 92862 215176 92867 215232
rect 90764 215174 92867 215176
rect 58301 215171 58367 215174
rect 92801 215171 92867 215174
rect 50389 215098 50455 215101
rect 47892 215096 50455 215098
rect 47892 215040 50394 215096
rect 50450 215040 50455 215096
rect 47892 215038 50455 215040
rect 50389 215035 50455 215038
rect 100989 215098 101055 215101
rect 103982 215098 104042 215408
rect 177717 215370 177783 215373
rect 174822 215368 177783 215370
rect 174822 215312 177722 215368
rect 177778 215312 177783 215368
rect 174822 215310 177783 215312
rect 142941 215234 143007 215237
rect 142941 215232 145044 215234
rect 142941 215176 142946 215232
rect 143002 215176 145044 215232
rect 174822 215204 174882 215310
rect 177717 215307 177783 215310
rect 142941 215174 145044 215176
rect 142941 215171 143007 215174
rect 134845 215098 134911 215101
rect 100989 215096 104042 215098
rect 100989 215040 100994 215096
rect 101050 215040 104042 215096
rect 100989 215038 104042 215040
rect 131796 215096 134911 215098
rect 131796 215040 134850 215096
rect 134906 215040 134911 215096
rect 131796 215038 134911 215040
rect 100989 215035 101055 215038
rect 134845 215035 134911 215038
rect 185721 215098 185787 215101
rect 185721 215096 187916 215098
rect 185721 215040 185726 215096
rect 185782 215040 187916 215096
rect 185721 215038 187916 215040
rect 185721 215035 185787 215038
rect 101817 214962 101883 214965
rect 177625 214962 177691 214965
rect 101817 214960 104012 214962
rect 101817 214904 101822 214960
rect 101878 214904 104012 214960
rect 101817 214902 104012 214904
rect 174822 214960 177691 214962
rect 174822 214904 177630 214960
rect 177686 214904 177691 214960
rect 174822 214902 177691 214904
rect 101817 214899 101883 214902
rect 51125 214554 51191 214557
rect 47892 214552 51191 214554
rect 47892 214496 51130 214552
rect 51186 214496 51191 214552
rect 47892 214494 51191 214496
rect 51125 214491 51191 214494
rect 58209 214554 58275 214557
rect 93537 214554 93603 214557
rect 135305 214554 135371 214557
rect 58209 214552 60956 214554
rect 58209 214496 58214 214552
rect 58270 214496 60956 214552
rect 58209 214494 60956 214496
rect 90764 214552 93603 214554
rect 90764 214496 93542 214552
rect 93598 214496 93603 214552
rect 90764 214494 93603 214496
rect 131796 214552 135371 214554
rect 131796 214496 135310 214552
rect 135366 214496 135371 214552
rect 131796 214494 135371 214496
rect 58209 214491 58275 214494
rect 93537 214491 93603 214494
rect 135305 214491 135371 214494
rect 143493 214554 143559 214557
rect 143493 214552 145044 214554
rect 143493 214496 143498 214552
rect 143554 214496 145044 214552
rect 174822 214524 174882 214902
rect 177625 214899 177691 214902
rect 185261 214554 185327 214557
rect 185261 214552 187916 214554
rect 143493 214494 145044 214496
rect 185261 214496 185266 214552
rect 185322 214496 187916 214552
rect 185261 214494 187916 214496
rect 143493 214491 143559 214494
rect 185261 214491 185327 214494
rect 50941 214010 51007 214013
rect 47892 214008 51007 214010
rect 47892 213952 50946 214008
rect 51002 213952 51007 214008
rect 47892 213950 51007 213952
rect 50941 213947 51007 213950
rect 58209 214010 58275 214013
rect 92801 214010 92867 214013
rect 58209 214008 60956 214010
rect 58209 213952 58214 214008
rect 58270 213952 60956 214008
rect 58209 213950 60956 213952
rect 90764 214008 92867 214010
rect 90764 213952 92806 214008
rect 92862 213952 92867 214008
rect 90764 213950 92867 213952
rect 58209 213947 58275 213950
rect 92801 213947 92867 213950
rect 100989 214010 101055 214013
rect 103982 214010 104042 214320
rect 177717 214146 177783 214149
rect 174822 214144 177783 214146
rect 174822 214088 177722 214144
rect 177778 214088 177783 214144
rect 174822 214086 177783 214088
rect 134661 214010 134727 214013
rect 100989 214008 104042 214010
rect 100989 213952 100994 214008
rect 101050 213952 104042 214008
rect 100989 213950 104042 213952
rect 131796 214008 134727 214010
rect 131796 213952 134666 214008
rect 134722 213952 134727 214008
rect 131796 213950 134727 213952
rect 100989 213947 101055 213950
rect 134661 213947 134727 213950
rect 142941 214010 143007 214013
rect 142941 214008 145044 214010
rect 142941 213952 142946 214008
rect 143002 213952 145044 214008
rect 174822 213980 174882 214086
rect 177717 214083 177783 214086
rect 185721 214010 185787 214013
rect 185721 214008 187916 214010
rect 142941 213950 145044 213952
rect 185721 213952 185726 214008
rect 185782 213952 187916 214008
rect 185721 213950 187916 213952
rect 142941 213947 143007 213950
rect 185721 213947 185787 213950
rect 50205 213466 50271 213469
rect 47892 213464 50271 213466
rect 47892 213408 50210 213464
rect 50266 213408 50271 213464
rect 47892 213406 50271 213408
rect 50205 213403 50271 213406
rect 101173 213466 101239 213469
rect 103982 213466 104042 213776
rect 177625 213738 177691 213741
rect 174822 213736 177691 213738
rect 174822 213680 177630 213736
rect 177686 213680 177691 213736
rect 174822 213678 177691 213680
rect 135397 213466 135463 213469
rect 101173 213464 104042 213466
rect 101173 213408 101178 213464
rect 101234 213408 104042 213464
rect 101173 213406 104042 213408
rect 131796 213464 135463 213466
rect 131796 213408 135402 213464
rect 135458 213408 135463 213464
rect 131796 213406 135463 213408
rect 101173 213403 101239 213406
rect 135397 213403 135463 213406
rect 58301 213330 58367 213333
rect 92709 213330 92775 213333
rect 58301 213328 60956 213330
rect 58301 213272 58306 213328
rect 58362 213272 60956 213328
rect 58301 213270 60956 213272
rect 90764 213328 92775 213330
rect 90764 213272 92714 213328
rect 92770 213272 92775 213328
rect 90764 213270 92775 213272
rect 58301 213267 58367 213270
rect 92709 213267 92775 213270
rect 143677 213330 143743 213333
rect 143677 213328 145044 213330
rect 143677 213272 143682 213328
rect 143738 213272 145044 213328
rect 174822 213300 174882 213678
rect 177625 213675 177691 213678
rect 185169 213466 185235 213469
rect 185169 213464 187916 213466
rect 185169 213408 185174 213464
rect 185230 213408 187916 213464
rect 185169 213406 187916 213408
rect 185169 213403 185235 213406
rect 143677 213270 145044 213272
rect 143677 213267 143743 213270
rect 103614 213202 104012 213262
rect 101081 213194 101147 213197
rect 103614 213194 103674 213202
rect 101081 213192 103674 213194
rect 101081 213136 101086 213192
rect 101142 213136 103674 213192
rect 101081 213134 103674 213136
rect 101081 213131 101147 213134
rect 50757 212922 50823 212925
rect 134845 212922 134911 212925
rect 177717 212922 177783 212925
rect 47892 212920 50823 212922
rect 47892 212864 50762 212920
rect 50818 212864 50823 212920
rect 47892 212862 50823 212864
rect 131796 212920 134911 212922
rect 131796 212864 134850 212920
rect 134906 212864 134911 212920
rect 131796 212862 134911 212864
rect 50757 212859 50823 212862
rect 134845 212859 134911 212862
rect 174822 212920 177783 212922
rect 174822 212864 177722 212920
rect 177778 212864 177783 212920
rect 174822 212862 177783 212864
rect 58209 212786 58275 212789
rect 92709 212786 92775 212789
rect 58209 212784 60956 212786
rect 58209 212728 58214 212784
rect 58270 212728 60956 212784
rect 58209 212726 60956 212728
rect 90764 212784 92775 212786
rect 90764 212728 92714 212784
rect 92770 212728 92775 212784
rect 90764 212726 92775 212728
rect 58209 212723 58275 212726
rect 92709 212723 92775 212726
rect 143677 212786 143743 212789
rect 143677 212784 145044 212786
rect 143677 212728 143682 212784
rect 143738 212728 145044 212784
rect 174822 212756 174882 212862
rect 177717 212859 177783 212862
rect 185721 212922 185787 212925
rect 185721 212920 187916 212922
rect 185721 212864 185726 212920
rect 185782 212864 187916 212920
rect 185721 212862 187916 212864
rect 185721 212859 185787 212862
rect 143677 212726 145044 212728
rect 143677 212723 143743 212726
rect 100989 212378 101055 212381
rect 103982 212378 104042 212688
rect 177717 212378 177783 212381
rect 100989 212376 104042 212378
rect 100989 212320 100994 212376
rect 101050 212320 104042 212376
rect 100989 212318 104042 212320
rect 174822 212376 177783 212378
rect 174822 212320 177722 212376
rect 177778 212320 177783 212376
rect 174822 212318 177783 212320
rect 100989 212315 101055 212318
rect 51217 212242 51283 212245
rect 47892 212240 51283 212242
rect 47892 212184 51222 212240
rect 51278 212184 51283 212240
rect 47892 212182 51283 212184
rect 51217 212179 51283 212182
rect 58301 212242 58367 212245
rect 93629 212242 93695 212245
rect 135397 212242 135463 212245
rect 58301 212240 60956 212242
rect 58301 212184 58306 212240
rect 58362 212184 60956 212240
rect 58301 212182 60956 212184
rect 90764 212240 93695 212242
rect 90764 212184 93634 212240
rect 93690 212184 93695 212240
rect 90764 212182 93695 212184
rect 131796 212240 135463 212242
rect 131796 212184 135402 212240
rect 135458 212184 135463 212240
rect 131796 212182 135463 212184
rect 58301 212179 58367 212182
rect 93629 212179 93695 212182
rect 135397 212179 135463 212182
rect 143493 212242 143559 212245
rect 143493 212240 145044 212242
rect 143493 212184 143498 212240
rect 143554 212184 145044 212240
rect 174822 212212 174882 212318
rect 177717 212315 177783 212318
rect 185905 212242 185971 212245
rect 185905 212240 187916 212242
rect 143493 212182 145044 212184
rect 185905 212184 185910 212240
rect 185966 212184 187916 212240
rect 185905 212182 187916 212184
rect 143493 212179 143559 212182
rect 185905 212179 185971 212182
rect 103614 212114 104012 212174
rect 101081 211970 101147 211973
rect 103614 211970 103674 212114
rect 101081 211968 103674 211970
rect 101081 211912 101086 211968
rect 101142 211912 103674 211968
rect 101081 211910 103674 211912
rect 101081 211907 101147 211910
rect 51125 211698 51191 211701
rect 135397 211698 135463 211701
rect 177717 211698 177783 211701
rect 47892 211696 51191 211698
rect 47892 211640 51130 211696
rect 51186 211640 51191 211696
rect 47892 211638 51191 211640
rect 131796 211696 135463 211698
rect 131796 211640 135402 211696
rect 135458 211640 135463 211696
rect 131796 211638 135463 211640
rect 51125 211635 51191 211638
rect 135397 211635 135463 211638
rect 174822 211696 177783 211698
rect 174822 211640 177722 211696
rect 177778 211640 177783 211696
rect 174822 211638 177783 211640
rect 58209 211562 58275 211565
rect 92709 211562 92775 211565
rect 58209 211560 60956 211562
rect 58209 211504 58214 211560
rect 58270 211504 60956 211560
rect 58209 211502 60956 211504
rect 90764 211560 92775 211562
rect 90764 211504 92714 211560
rect 92770 211504 92775 211560
rect 90764 211502 92775 211504
rect 58209 211499 58275 211502
rect 92709 211499 92775 211502
rect 143677 211562 143743 211565
rect 143677 211560 145044 211562
rect 143677 211504 143682 211560
rect 143738 211504 145044 211560
rect 174822 211532 174882 211638
rect 177717 211635 177783 211638
rect 185721 211698 185787 211701
rect 185721 211696 187916 211698
rect 185721 211640 185726 211696
rect 185782 211640 187916 211696
rect 185721 211638 187916 211640
rect 185721 211635 185787 211638
rect 216909 211562 216975 211565
rect 215884 211560 216975 211562
rect 143677 211502 145044 211504
rect 215884 211504 216914 211560
rect 216970 211504 216975 211560
rect 215884 211502 216975 211504
rect 143677 211499 143743 211502
rect 216909 211499 216975 211502
rect 50665 211154 50731 211157
rect 47892 211152 50731 211154
rect 47892 211096 50670 211152
rect 50726 211096 50731 211152
rect 47892 211094 50731 211096
rect 50665 211091 50731 211094
rect 101173 211154 101239 211157
rect 103982 211154 104042 211464
rect 135029 211154 135095 211157
rect 177717 211154 177783 211157
rect 101173 211152 104042 211154
rect 101173 211096 101178 211152
rect 101234 211096 104042 211152
rect 101173 211094 104042 211096
rect 131796 211152 135095 211154
rect 131796 211096 135034 211152
rect 135090 211096 135095 211152
rect 131796 211094 135095 211096
rect 101173 211091 101239 211094
rect 135029 211091 135095 211094
rect 174822 211152 177783 211154
rect 174822 211096 177722 211152
rect 177778 211096 177783 211152
rect 174822 211094 177783 211096
rect 58301 211018 58367 211021
rect 92801 211018 92867 211021
rect 58301 211016 60956 211018
rect 58301 210960 58306 211016
rect 58362 210960 60956 211016
rect 58301 210958 60956 210960
rect 90764 211016 92867 211018
rect 90764 210960 92806 211016
rect 92862 210960 92867 211016
rect 90764 210958 92867 210960
rect 58301 210955 58367 210958
rect 92801 210955 92867 210958
rect 143677 211018 143743 211021
rect 143677 211016 145044 211018
rect 143677 210960 143682 211016
rect 143738 210960 145044 211016
rect 174822 210988 174882 211094
rect 177717 211091 177783 211094
rect 185813 211154 185879 211157
rect 185813 211152 187916 211154
rect 185813 211096 185818 211152
rect 185874 211096 187916 211152
rect 185813 211094 187916 211096
rect 185813 211091 185879 211094
rect 143677 210958 145044 210960
rect 143677 210955 143743 210958
rect 101081 210746 101147 210749
rect 103982 210746 104042 210920
rect 177717 210746 177783 210749
rect 101081 210744 104042 210746
rect 101081 210688 101086 210744
rect 101142 210688 104042 210744
rect 101081 210686 104042 210688
rect 174822 210744 177783 210746
rect 174822 210688 177722 210744
rect 177778 210688 177783 210744
rect 174822 210686 177783 210688
rect 101081 210683 101147 210686
rect 50849 210610 50915 210613
rect 134845 210610 134911 210613
rect 47892 210608 50915 210610
rect 47892 210552 50854 210608
rect 50910 210552 50915 210608
rect 47892 210550 50915 210552
rect 131796 210608 134911 210610
rect 131796 210552 134850 210608
rect 134906 210552 134911 210608
rect 131796 210550 134911 210552
rect 50849 210547 50915 210550
rect 134845 210547 134911 210550
rect 100989 210474 101055 210477
rect 100989 210472 104012 210474
rect 100989 210416 100994 210472
rect 101050 210416 104012 210472
rect 100989 210414 104012 210416
rect 100989 210411 101055 210414
rect 58393 210338 58459 210341
rect 93537 210338 93603 210341
rect 58393 210336 60956 210338
rect 58393 210280 58398 210336
rect 58454 210280 60956 210336
rect 58393 210278 60956 210280
rect 90764 210336 93603 210338
rect 90764 210280 93542 210336
rect 93598 210280 93603 210336
rect 90764 210278 93603 210280
rect 58393 210275 58459 210278
rect 93537 210275 93603 210278
rect 143585 210338 143651 210341
rect 143585 210336 145044 210338
rect 143585 210280 143590 210336
rect 143646 210280 145044 210336
rect 174822 210308 174882 210686
rect 177717 210683 177783 210686
rect 185997 210610 186063 210613
rect 185997 210608 187916 210610
rect 185997 210552 186002 210608
rect 186058 210552 187916 210608
rect 185997 210550 187916 210552
rect 185997 210547 186063 210550
rect 143585 210278 145044 210280
rect 143585 210275 143651 210278
rect 50757 210066 50823 210069
rect 135121 210066 135187 210069
rect 47892 210064 50823 210066
rect 47892 210008 50762 210064
rect 50818 210008 50823 210064
rect 47892 210006 50823 210008
rect 131796 210064 135187 210066
rect 131796 210008 135126 210064
rect 135182 210008 135187 210064
rect 131796 210006 135187 210008
rect 50757 210003 50823 210006
rect 135121 210003 135187 210006
rect 185721 210066 185787 210069
rect 185721 210064 187916 210066
rect 185721 210008 185726 210064
rect 185782 210008 187916 210064
rect 185721 210006 187916 210008
rect 185721 210003 185787 210006
rect 177717 209930 177783 209933
rect 174822 209928 177783 209930
rect 174822 209872 177722 209928
rect 177778 209872 177783 209928
rect 174822 209870 177783 209872
rect 58209 209794 58275 209797
rect 92709 209794 92775 209797
rect 58209 209792 60956 209794
rect 58209 209736 58214 209792
rect 58270 209736 60956 209792
rect 58209 209734 60956 209736
rect 90764 209792 92775 209794
rect 90764 209736 92714 209792
rect 92770 209736 92775 209792
rect 90764 209734 92775 209736
rect 58209 209731 58275 209734
rect 92709 209731 92775 209734
rect 101081 209522 101147 209525
rect 103982 209522 104042 209832
rect 142941 209794 143007 209797
rect 142941 209792 145044 209794
rect 142941 209736 142946 209792
rect 143002 209736 145044 209792
rect 174822 209764 174882 209870
rect 177717 209867 177783 209870
rect 142941 209734 145044 209736
rect 142941 209731 143007 209734
rect 178177 209522 178243 209525
rect 101081 209520 104042 209522
rect 101081 209464 101086 209520
rect 101142 209464 104042 209520
rect 101081 209462 104042 209464
rect 174822 209520 178243 209522
rect 174822 209464 178182 209520
rect 178238 209464 178243 209520
rect 174822 209462 178243 209464
rect 101081 209459 101147 209462
rect 9896 209386 10376 209416
rect 13313 209386 13379 209389
rect 50941 209386 51007 209389
rect 134937 209386 135003 209389
rect 9896 209384 13379 209386
rect 9896 209328 13318 209384
rect 13374 209328 13379 209384
rect 9896 209326 13379 209328
rect 47892 209384 51007 209386
rect 47892 209328 50946 209384
rect 51002 209328 51007 209384
rect 47892 209326 51007 209328
rect 131796 209384 135003 209386
rect 131796 209328 134942 209384
rect 134998 209328 135003 209384
rect 131796 209326 135003 209328
rect 9896 209296 10376 209326
rect 13313 209323 13379 209326
rect 50941 209323 51007 209326
rect 134937 209323 135003 209326
rect 58301 209250 58367 209253
rect 94089 209250 94155 209253
rect 58301 209248 60956 209250
rect 58301 209192 58306 209248
rect 58362 209192 60956 209248
rect 58301 209190 60956 209192
rect 90764 209248 94155 209250
rect 90764 209192 94094 209248
rect 94150 209192 94155 209248
rect 90764 209190 94155 209192
rect 58301 209187 58367 209190
rect 94089 209187 94155 209190
rect 100989 209114 101055 209117
rect 103982 209114 104042 209288
rect 143677 209250 143743 209253
rect 143677 209248 145044 209250
rect 143677 209192 143682 209248
rect 143738 209192 145044 209248
rect 174822 209220 174882 209462
rect 178177 209459 178243 209462
rect 185813 209386 185879 209389
rect 185813 209384 187916 209386
rect 185813 209328 185818 209384
rect 185874 209328 187916 209384
rect 185813 209326 187916 209328
rect 185813 209323 185879 209326
rect 143677 209190 145044 209192
rect 143677 209187 143743 209190
rect 100989 209112 104042 209114
rect 100989 209056 100994 209112
rect 101050 209056 104042 209112
rect 100989 209054 104042 209056
rect 100989 209051 101055 209054
rect 169897 208978 169963 208981
rect 171134 208978 171140 208980
rect 169897 208976 171140 208978
rect 169897 208920 169902 208976
rect 169958 208920 171140 208976
rect 169897 208918 171140 208920
rect 169897 208915 169963 208918
rect 171134 208916 171140 208918
rect 171204 208916 171210 208980
rect 51125 208842 51191 208845
rect 135305 208842 135371 208845
rect 47892 208840 51191 208842
rect 47892 208784 51130 208840
rect 51186 208784 51191 208840
rect 47892 208782 51191 208784
rect 131796 208840 135371 208842
rect 131796 208784 135310 208840
rect 135366 208784 135371 208840
rect 131796 208782 135371 208784
rect 51125 208779 51191 208782
rect 135305 208779 135371 208782
rect 186089 208842 186155 208845
rect 186089 208840 187916 208842
rect 186089 208784 186094 208840
rect 186150 208784 187916 208840
rect 186089 208782 187916 208784
rect 186089 208779 186155 208782
rect 102093 208434 102159 208437
rect 103982 208434 104042 208744
rect 102093 208432 104042 208434
rect 102093 208376 102098 208432
rect 102154 208376 104042 208432
rect 102093 208374 104042 208376
rect 102093 208371 102159 208374
rect 51033 208298 51099 208301
rect 135213 208298 135279 208301
rect 47892 208296 51099 208298
rect 47892 208240 51038 208296
rect 51094 208240 51099 208296
rect 47892 208238 51099 208240
rect 131796 208296 135279 208298
rect 131796 208240 135218 208296
rect 135274 208240 135279 208296
rect 131796 208238 135279 208240
rect 51033 208235 51099 208238
rect 135213 208235 135279 208238
rect 186273 208298 186339 208301
rect 186273 208296 187916 208298
rect 186273 208240 186278 208296
rect 186334 208240 187916 208296
rect 186273 208238 187916 208240
rect 186273 208235 186339 208238
rect 101909 207890 101975 207893
rect 103982 207890 104042 208200
rect 101909 207888 104042 207890
rect 101909 207832 101914 207888
rect 101970 207832 104042 207888
rect 101909 207830 104042 207832
rect 101909 207827 101975 207830
rect 51217 207754 51283 207757
rect 135397 207754 135463 207757
rect 47892 207752 51283 207754
rect 47892 207696 51222 207752
rect 51278 207696 51283 207752
rect 47892 207694 51283 207696
rect 131796 207752 135463 207754
rect 131796 207696 135402 207752
rect 135458 207696 135463 207752
rect 131796 207694 135463 207696
rect 51217 207691 51283 207694
rect 135397 207691 135463 207694
rect 185997 207754 186063 207757
rect 185997 207752 187916 207754
rect 185997 207696 186002 207752
rect 186058 207696 187916 207752
rect 185997 207694 187916 207696
rect 185997 207691 186063 207694
rect 103614 207626 104012 207686
rect 101725 207618 101791 207621
rect 103614 207618 103674 207626
rect 101725 207616 103674 207618
rect 101725 207560 101730 207616
rect 101786 207560 103674 207616
rect 101725 207558 103674 207560
rect 101725 207555 101791 207558
rect 85717 207482 85783 207485
rect 88518 207482 88524 207484
rect 85717 207480 88524 207482
rect 85717 207424 85722 207480
rect 85778 207424 88524 207480
rect 85717 207422 88524 207424
rect 85717 207419 85783 207422
rect 88518 207420 88524 207422
rect 88588 207420 88594 207484
rect 51125 207210 51191 207213
rect 135305 207210 135371 207213
rect 47892 207208 51191 207210
rect 47892 207152 51130 207208
rect 51186 207152 51191 207208
rect 47892 207150 51191 207152
rect 131796 207208 135371 207210
rect 131796 207152 135310 207208
rect 135366 207152 135371 207208
rect 131796 207150 135371 207152
rect 51125 207147 51191 207150
rect 135305 207147 135371 207150
rect 185169 207210 185235 207213
rect 185169 207208 187916 207210
rect 185169 207152 185174 207208
rect 185230 207152 187916 207208
rect 185169 207150 187916 207152
rect 185169 207147 185235 207150
rect 100989 206530 101055 206533
rect 103982 206530 104042 207112
rect 187929 206938 187995 206941
rect 189166 206938 189172 206940
rect 187929 206936 189172 206938
rect 187929 206880 187934 206936
rect 187990 206880 189172 206936
rect 187929 206878 189172 206880
rect 187929 206875 187995 206878
rect 189166 206876 189172 206878
rect 189236 206876 189242 206940
rect 100989 206528 104042 206530
rect 100989 206472 100994 206528
rect 101050 206472 104042 206528
rect 100989 206470 104042 206472
rect 100989 206467 101055 206470
rect 220313 205442 220379 205445
rect 225416 205442 225896 205472
rect 220313 205440 225896 205442
rect 220313 205384 220318 205440
rect 220374 205384 225896 205440
rect 220313 205382 225896 205384
rect 220313 205379 220379 205382
rect 225416 205352 225896 205382
rect 140222 195180 140228 195244
rect 140292 195242 140298 195244
rect 167137 195242 167203 195245
rect 140292 195240 167203 195242
rect 140292 195184 167142 195240
rect 167198 195184 167203 195240
rect 140292 195182 167203 195184
rect 140292 195180 140298 195182
rect 167137 195179 167203 195182
rect 99517 193746 99583 193749
rect 95702 193744 99583 193746
rect 95702 193688 99522 193744
rect 99578 193688 99583 193744
rect 95702 193686 99583 193688
rect 95702 193240 95762 193686
rect 99517 193683 99583 193686
rect 182869 193202 182935 193205
rect 179820 193200 182935 193202
rect 179820 193144 182874 193200
rect 182930 193144 182935 193200
rect 179820 193142 182935 193144
rect 182869 193139 182935 193142
rect 191977 192794 192043 192797
rect 191977 192792 193988 192794
rect 191977 192736 191982 192792
rect 192038 192736 193988 192792
rect 191977 192734 193988 192736
rect 191977 192731 192043 192734
rect 105773 192522 105839 192525
rect 105773 192520 109900 192522
rect 105773 192464 105778 192520
rect 105834 192464 109900 192520
rect 105773 192462 109900 192464
rect 105773 192459 105839 192462
rect 99425 192386 99491 192389
rect 95702 192384 99491 192386
rect 95702 192328 99430 192384
rect 99486 192328 99491 192384
rect 95702 192326 99491 192328
rect 95702 192016 95762 192326
rect 99425 192323 99491 192326
rect 183605 191978 183671 191981
rect 179820 191976 183671 191978
rect 179820 191920 183610 191976
rect 183666 191920 183671 191976
rect 179820 191918 183671 191920
rect 183605 191915 183671 191918
rect 99241 190754 99307 190757
rect 183421 190754 183487 190757
rect 209917 190756 209983 190757
rect 209917 190754 209964 190756
rect 95732 190752 99307 190754
rect 95732 190696 99246 190752
rect 99302 190696 99307 190752
rect 95732 190694 99307 190696
rect 179820 190752 183487 190754
rect 179820 190696 183426 190752
rect 183482 190696 183487 190752
rect 209876 190752 209964 190754
rect 210028 190754 210034 190756
rect 179820 190694 183487 190696
rect 99241 190691 99307 190694
rect 183421 190691 183487 190694
rect 193958 190620 194018 190724
rect 209876 190696 209922 190752
rect 209876 190694 209964 190696
rect 209917 190692 209964 190694
rect 210028 190694 210110 190754
rect 210028 190692 210034 190694
rect 209917 190691 209983 190692
rect 193950 190556 193956 190620
rect 194020 190556 194026 190620
rect 22329 190482 22395 190485
rect 212125 190482 212191 190485
rect 22329 190480 25996 190482
rect 22329 190424 22334 190480
rect 22390 190424 25996 190480
rect 22329 190422 25996 190424
rect 209812 190480 212191 190482
rect 209812 190424 212130 190480
rect 212186 190424 212191 190480
rect 209812 190422 212191 190424
rect 22329 190419 22395 190422
rect 212125 190419 212191 190422
rect 107153 190210 107219 190213
rect 107153 190208 109900 190210
rect 107153 190152 107158 190208
rect 107214 190152 109900 190208
rect 107153 190150 109900 190152
rect 107153 190147 107219 190150
rect 99149 189530 99215 189533
rect 183329 189530 183395 189533
rect 95732 189528 99215 189530
rect 95732 189472 99154 189528
rect 99210 189472 99215 189528
rect 95732 189470 99215 189472
rect 179820 189528 183395 189530
rect 179820 189472 183334 189528
rect 183390 189472 183395 189528
rect 179820 189470 183395 189472
rect 99149 189467 99215 189470
rect 183329 189467 183395 189470
rect 41833 189258 41899 189261
rect 41790 189256 41899 189258
rect 41790 189200 41838 189256
rect 41894 189200 41899 189256
rect 41790 189195 41899 189200
rect 41790 188684 41850 189195
rect 99333 188986 99399 188989
rect 95702 188984 99399 188986
rect 95702 188928 99338 188984
rect 99394 188928 99399 188984
rect 95702 188926 99399 188928
rect 95702 188344 95762 188926
rect 99333 188923 99399 188926
rect 191977 188714 192043 188717
rect 191977 188712 193988 188714
rect 191977 188656 191982 188712
rect 192038 188656 193988 188712
rect 191977 188654 193988 188656
rect 191977 188651 192043 188654
rect 183513 188306 183579 188309
rect 179820 188304 183579 188306
rect 179820 188248 183518 188304
rect 183574 188248 183579 188304
rect 179820 188246 183579 188248
rect 183513 188243 183579 188246
rect 106785 187898 106851 187901
rect 106785 187896 109900 187898
rect 106785 187840 106790 187896
rect 106846 187840 109900 187896
rect 106785 187838 109900 187840
rect 106785 187835 106851 187838
rect 99057 187762 99123 187765
rect 95702 187760 99123 187762
rect 95702 187704 99062 187760
rect 99118 187704 99123 187760
rect 95702 187702 99123 187704
rect 95702 187120 95762 187702
rect 99057 187699 99123 187702
rect 183237 187082 183303 187085
rect 179820 187080 183303 187082
rect 179820 187024 183242 187080
rect 183298 187024 183303 187080
rect 179820 187022 183303 187024
rect 183237 187019 183303 187022
rect 191149 186810 191215 186813
rect 191149 186808 193988 186810
rect 191149 186752 191154 186808
rect 191210 186752 193988 186808
rect 191149 186750 193988 186752
rect 191149 186747 191215 186750
rect 98965 186538 99031 186541
rect 95702 186536 99031 186538
rect 95702 186480 98970 186536
rect 99026 186480 99031 186536
rect 95702 186478 99031 186480
rect 95702 185896 95762 186478
rect 98965 186475 99031 186478
rect 183145 185858 183211 185861
rect 179820 185856 183211 185858
rect 179820 185800 183150 185856
rect 183206 185800 183211 185856
rect 179820 185798 183211 185800
rect 183145 185795 183211 185798
rect 9896 185722 10376 185752
rect 13405 185722 13471 185725
rect 9896 185720 13471 185722
rect 9896 185664 13410 185720
rect 13466 185664 13471 185720
rect 9896 185662 13471 185664
rect 9896 185632 10376 185662
rect 13405 185659 13471 185662
rect 106785 185450 106851 185453
rect 106785 185448 109900 185450
rect 106785 185392 106790 185448
rect 106846 185392 109900 185448
rect 106785 185390 109900 185392
rect 106785 185387 106851 185390
rect 98873 185314 98939 185317
rect 95702 185312 98939 185314
rect 95702 185256 98878 185312
rect 98934 185256 98939 185312
rect 95702 185254 98939 185256
rect 95702 184672 95762 185254
rect 98873 185251 98939 185254
rect 191977 184770 192043 184773
rect 191977 184768 193988 184770
rect 191977 184712 191982 184768
rect 192038 184712 193988 184768
rect 191977 184710 193988 184712
rect 191977 184707 192043 184710
rect 183053 184634 183119 184637
rect 179820 184632 183119 184634
rect 179820 184576 183058 184632
rect 183114 184576 183119 184632
rect 179820 184574 183119 184576
rect 183053 184571 183119 184574
rect 22329 183818 22395 183821
rect 128497 183818 128563 183821
rect 212033 183818 212099 183821
rect 22329 183816 25996 183818
rect 22329 183760 22334 183816
rect 22390 183760 25996 183816
rect 22329 183758 25996 183760
rect 125724 183816 128563 183818
rect 125724 183760 128502 183816
rect 128558 183760 128563 183816
rect 125724 183758 128563 183760
rect 209812 183816 212099 183818
rect 209812 183760 212038 183816
rect 212094 183760 212099 183816
rect 209812 183758 212099 183760
rect 22329 183755 22395 183758
rect 128497 183755 128563 183758
rect 212033 183755 212099 183758
rect 99517 183682 99583 183685
rect 95702 183680 99583 183682
rect 95702 183624 99522 183680
rect 99578 183624 99583 183680
rect 95702 183622 99583 183624
rect 95702 183448 95762 183622
rect 99517 183619 99583 183622
rect 182869 183410 182935 183413
rect 179820 183408 182935 183410
rect 179820 183352 182874 183408
rect 182930 183352 182935 183408
rect 179820 183350 182935 183352
rect 182869 183347 182935 183350
rect 107153 183138 107219 183141
rect 107153 183136 109900 183138
rect 107153 183080 107158 183136
rect 107214 183080 109900 183136
rect 107153 183078 109900 183080
rect 107153 183075 107219 183078
rect 190597 182730 190663 182733
rect 190597 182728 193988 182730
rect 190597 182672 190602 182728
rect 190658 182672 193988 182728
rect 190597 182670 193988 182672
rect 190597 182667 190663 182670
rect 98597 182458 98663 182461
rect 95702 182456 98663 182458
rect 95702 182400 98602 182456
rect 98658 182400 98663 182456
rect 95702 182398 98663 182400
rect 95702 182224 95762 182398
rect 98597 182395 98663 182398
rect 183145 182186 183211 182189
rect 179820 182184 183211 182186
rect 179820 182128 183150 182184
rect 183206 182128 183211 182184
rect 179820 182126 183211 182128
rect 183145 182123 183211 182126
rect 99425 181098 99491 181101
rect 183697 181098 183763 181101
rect 95732 181096 99491 181098
rect 95732 181040 99430 181096
rect 99486 181040 99491 181096
rect 95732 181038 99491 181040
rect 179820 181096 183763 181098
rect 179820 181040 183702 181096
rect 183758 181040 183763 181096
rect 179820 181038 183763 181040
rect 99425 181035 99491 181038
rect 183697 181035 183763 181038
rect 106969 180826 107035 180829
rect 190689 180826 190755 180829
rect 106969 180824 109900 180826
rect 106969 180768 106974 180824
rect 107030 180768 109900 180824
rect 106969 180766 109900 180768
rect 190689 180824 193988 180826
rect 190689 180768 190694 180824
rect 190750 180768 193988 180824
rect 190689 180766 193988 180768
rect 106969 180763 107035 180766
rect 190689 180763 190755 180766
rect 99517 179874 99583 179877
rect 183697 179874 183763 179877
rect 95732 179872 99583 179874
rect 95732 179816 99522 179872
rect 99578 179816 99583 179872
rect 95732 179814 99583 179816
rect 179820 179872 183763 179874
rect 179820 179816 183702 179872
rect 183758 179816 183763 179872
rect 179820 179814 183763 179816
rect 99517 179811 99583 179814
rect 183697 179811 183763 179814
rect 98413 179330 98479 179333
rect 95702 179328 98479 179330
rect 95702 179272 98418 179328
rect 98474 179272 98479 179328
rect 95702 179270 98479 179272
rect 44409 178786 44475 178789
rect 41820 178784 44475 178786
rect 41820 178728 44414 178784
rect 44470 178728 44475 178784
rect 41820 178726 44475 178728
rect 44409 178723 44475 178726
rect 95702 178688 95762 179270
rect 98413 179267 98479 179270
rect 222337 179194 222403 179197
rect 225416 179194 225896 179224
rect 222337 179192 225896 179194
rect 222337 179136 222342 179192
rect 222398 179136 225896 179192
rect 222337 179134 225896 179136
rect 222337 179131 222403 179134
rect 225416 179104 225896 179134
rect 191977 178786 192043 178789
rect 191977 178784 193988 178786
rect 191977 178728 191982 178784
rect 192038 178728 193988 178784
rect 191977 178726 193988 178728
rect 191977 178723 192043 178726
rect 182501 178650 182567 178653
rect 179820 178648 182567 178650
rect 179820 178592 182506 178648
rect 182562 178592 182567 178648
rect 179820 178590 182567 178592
rect 182501 178587 182567 178590
rect 106785 178378 106851 178381
rect 106785 178376 109900 178378
rect 106785 178320 106790 178376
rect 106846 178320 109900 178376
rect 106785 178318 109900 178320
rect 106785 178315 106851 178318
rect 99517 177426 99583 177429
rect 182501 177426 182567 177429
rect 95732 177424 99583 177426
rect 95732 177368 99522 177424
rect 99578 177368 99583 177424
rect 95732 177366 99583 177368
rect 179820 177424 182567 177426
rect 179820 177368 182506 177424
rect 182562 177368 182567 177424
rect 179820 177366 182567 177368
rect 99517 177363 99583 177366
rect 182501 177363 182567 177366
rect 22329 177154 22395 177157
rect 211573 177154 211639 177157
rect 22329 177152 25996 177154
rect 22329 177096 22334 177152
rect 22390 177096 25996 177152
rect 22329 177094 25996 177096
rect 209812 177152 211639 177154
rect 209812 177096 211578 177152
rect 211634 177096 211639 177152
rect 209812 177094 211639 177096
rect 22329 177091 22395 177094
rect 211573 177091 211639 177094
rect 98597 176746 98663 176749
rect 95702 176744 98663 176746
rect 95702 176688 98602 176744
rect 98658 176688 98663 176744
rect 95702 176686 98663 176688
rect 95702 176240 95762 176686
rect 98597 176683 98663 176686
rect 191977 176746 192043 176749
rect 191977 176744 193988 176746
rect 191977 176688 191982 176744
rect 192038 176688 193988 176744
rect 191977 176686 193988 176688
rect 191977 176683 192043 176686
rect 183237 176202 183303 176205
rect 179820 176200 183303 176202
rect 179820 176144 183242 176200
rect 183298 176144 183303 176200
rect 179820 176142 183303 176144
rect 183237 176139 183303 176142
rect 106601 176066 106667 176069
rect 106601 176064 109900 176066
rect 106601 176008 106606 176064
rect 106662 176008 109900 176064
rect 106601 176006 109900 176008
rect 106601 176003 106667 176006
rect 98229 175386 98295 175389
rect 95702 175384 98295 175386
rect 95702 175328 98234 175384
rect 98290 175328 98295 175384
rect 95702 175326 98295 175328
rect 95702 175016 95762 175326
rect 98229 175323 98295 175326
rect 183697 174978 183763 174981
rect 179820 174976 183763 174978
rect 179820 174920 183702 174976
rect 183758 174920 183763 174976
rect 179820 174918 183763 174920
rect 183697 174915 183763 174918
rect 191517 174842 191583 174845
rect 191517 174840 193988 174842
rect 191517 174784 191522 174840
rect 191578 174784 193988 174840
rect 191517 174782 193988 174784
rect 191517 174779 191583 174782
rect 137513 174434 137579 174437
rect 137513 174432 140106 174434
rect 137513 174376 137518 174432
rect 137574 174376 140106 174432
rect 137513 174374 140106 174376
rect 137513 174371 137579 174374
rect 140046 173928 140106 174374
rect 52689 173890 52755 173893
rect 52689 173888 55988 173890
rect 52689 173832 52694 173888
rect 52750 173832 55988 173888
rect 52689 173830 55988 173832
rect 52689 173827 52755 173830
rect 99517 173754 99583 173757
rect 95732 173752 99583 173754
rect 95732 173696 99522 173752
rect 99578 173696 99583 173752
rect 95732 173694 99583 173696
rect 99517 173691 99583 173694
rect 106785 173754 106851 173757
rect 183329 173754 183395 173757
rect 106785 173752 109900 173754
rect 106785 173696 106790 173752
rect 106846 173696 109900 173752
rect 106785 173694 109900 173696
rect 179820 173752 183395 173754
rect 179820 173696 183334 173752
rect 183390 173696 183395 173752
rect 179820 173694 183395 173696
rect 106785 173691 106851 173694
rect 183329 173691 183395 173694
rect 191977 172802 192043 172805
rect 191977 172800 193988 172802
rect 191977 172744 191982 172800
rect 192038 172744 193988 172800
rect 191977 172742 193988 172744
rect 191977 172739 192043 172742
rect 99517 172530 99583 172533
rect 183513 172530 183579 172533
rect 95732 172528 99583 172530
rect 95732 172472 99522 172528
rect 99578 172472 99583 172528
rect 95732 172470 99583 172472
rect 179820 172528 183579 172530
rect 179820 172472 183518 172528
rect 183574 172472 183579 172528
rect 179820 172470 183579 172472
rect 99517 172467 99583 172470
rect 183513 172467 183579 172470
rect 106785 171442 106851 171445
rect 106785 171440 109900 171442
rect 106785 171384 106790 171440
rect 106846 171384 109900 171440
rect 106785 171382 109900 171384
rect 106785 171379 106851 171382
rect 99241 171306 99307 171309
rect 182685 171306 182751 171309
rect 95732 171304 99307 171306
rect 95732 171248 99246 171304
rect 99302 171248 99307 171304
rect 95732 171246 99307 171248
rect 179820 171304 182751 171306
rect 179820 171248 182690 171304
rect 182746 171248 182751 171304
rect 179820 171246 182751 171248
rect 99241 171243 99307 171246
rect 182685 171243 182751 171246
rect 209825 171034 209891 171037
rect 209782 171032 209891 171034
rect 209782 170976 209830 171032
rect 209886 170976 209891 171032
rect 209782 170971 209891 170976
rect 191149 170762 191215 170765
rect 191149 170760 193988 170762
rect 191149 170704 191154 170760
rect 191210 170704 193988 170760
rect 191149 170702 193988 170704
rect 191149 170699 191215 170702
rect 22973 170490 23039 170493
rect 22973 170488 25996 170490
rect 22973 170432 22978 170488
rect 23034 170432 25996 170488
rect 209782 170460 209842 170971
rect 22973 170430 25996 170432
rect 22973 170427 23039 170430
rect 99517 170082 99583 170085
rect 182501 170082 182567 170085
rect 95732 170080 99583 170082
rect 95732 170024 99522 170080
rect 99578 170024 99583 170080
rect 95732 170022 99583 170024
rect 179820 170080 182567 170082
rect 179820 170024 182506 170080
rect 182562 170024 182567 170080
rect 179820 170022 182567 170024
rect 99517 170019 99583 170022
rect 182501 170019 182567 170022
rect 106785 168994 106851 168997
rect 106785 168992 109900 168994
rect 106785 168936 106790 168992
rect 106846 168936 109900 168992
rect 106785 168934 109900 168936
rect 106785 168931 106851 168934
rect 99425 168858 99491 168861
rect 183697 168858 183763 168861
rect 95732 168856 99491 168858
rect 95732 168800 99430 168856
rect 99486 168800 99491 168856
rect 95732 168798 99491 168800
rect 179820 168856 183763 168858
rect 179820 168800 183702 168856
rect 183758 168800 183763 168856
rect 179820 168798 183763 168800
rect 99425 168795 99491 168798
rect 183697 168795 183763 168798
rect 44409 168722 44475 168725
rect 41820 168720 44475 168722
rect 41820 168664 44414 168720
rect 44470 168664 44475 168720
rect 41820 168662 44475 168664
rect 44409 168659 44475 168662
rect 191977 168722 192043 168725
rect 191977 168720 193988 168722
rect 191977 168664 191982 168720
rect 192038 168664 193988 168720
rect 191977 168662 193988 168664
rect 191977 168659 192043 168662
rect 99517 167770 99583 167773
rect 183789 167770 183855 167773
rect 95732 167768 99583 167770
rect 95732 167712 99522 167768
rect 99578 167712 99583 167768
rect 95732 167710 99583 167712
rect 179820 167768 183855 167770
rect 179820 167712 183794 167768
rect 183850 167712 183855 167768
rect 179820 167710 183855 167712
rect 99517 167707 99583 167710
rect 183789 167707 183855 167710
rect 191885 166818 191951 166821
rect 191885 166816 193988 166818
rect 191885 166760 191890 166816
rect 191946 166760 193988 166816
rect 191885 166758 193988 166760
rect 191885 166755 191951 166758
rect 106693 166682 106759 166685
rect 106693 166680 109900 166682
rect 106693 166624 106698 166680
rect 106754 166624 109900 166680
rect 106693 166622 109900 166624
rect 106693 166619 106759 166622
rect 99517 166546 99583 166549
rect 182869 166546 182935 166549
rect 95732 166544 99583 166546
rect 95732 166488 99522 166544
rect 99578 166488 99583 166544
rect 95732 166486 99583 166488
rect 179820 166544 182935 166546
rect 179820 166488 182874 166544
rect 182930 166488 182935 166544
rect 179820 166486 182935 166488
rect 99517 166483 99583 166486
rect 182869 166483 182935 166486
rect 99517 165322 99583 165325
rect 183697 165322 183763 165325
rect 95732 165320 99583 165322
rect 95732 165264 99522 165320
rect 99578 165264 99583 165320
rect 95732 165262 99583 165264
rect 179820 165320 183763 165322
rect 179820 165264 183702 165320
rect 183758 165264 183763 165320
rect 179820 165262 183763 165264
rect 99517 165259 99583 165262
rect 183697 165259 183763 165262
rect 191333 164778 191399 164781
rect 191333 164776 193988 164778
rect 191333 164720 191338 164776
rect 191394 164720 193988 164776
rect 191333 164718 193988 164720
rect 191333 164715 191399 164718
rect 106785 164370 106851 164373
rect 106785 164368 109900 164370
rect 106785 164312 106790 164368
rect 106846 164312 109900 164368
rect 106785 164310 109900 164312
rect 106785 164307 106851 164310
rect 99517 164098 99583 164101
rect 183053 164098 183119 164101
rect 95732 164096 99583 164098
rect 95732 164040 99522 164096
rect 99578 164040 99583 164096
rect 95732 164038 99583 164040
rect 179820 164096 183119 164098
rect 179820 164040 183058 164096
rect 183114 164040 183119 164096
rect 179820 164038 183119 164040
rect 99517 164035 99583 164038
rect 183053 164035 183119 164038
rect 23617 163826 23683 163829
rect 128497 163826 128563 163829
rect 211757 163826 211823 163829
rect 23617 163824 25996 163826
rect 23617 163768 23622 163824
rect 23678 163768 25996 163824
rect 23617 163766 25996 163768
rect 125724 163824 128563 163826
rect 125724 163768 128502 163824
rect 128558 163768 128563 163824
rect 125724 163766 128563 163768
rect 209812 163824 211823 163826
rect 209812 163768 211762 163824
rect 211818 163768 211823 163824
rect 209812 163766 211823 163768
rect 23617 163763 23683 163766
rect 128497 163763 128563 163766
rect 211757 163763 211823 163766
rect 98965 162874 99031 162877
rect 183053 162874 183119 162877
rect 95732 162872 99031 162874
rect 95732 162816 98970 162872
rect 99026 162816 99031 162872
rect 95732 162814 99031 162816
rect 179820 162872 183119 162874
rect 179820 162816 183058 162872
rect 183114 162816 183119 162872
rect 179820 162814 183119 162816
rect 98965 162811 99031 162814
rect 183053 162811 183119 162814
rect 191517 162738 191583 162741
rect 191517 162736 193988 162738
rect 191517 162680 191522 162736
rect 191578 162680 193988 162736
rect 191517 162678 193988 162680
rect 191517 162675 191583 162678
rect 9896 162194 10376 162224
rect 13129 162194 13195 162197
rect 9896 162192 13195 162194
rect 9896 162136 13134 162192
rect 13190 162136 13195 162192
rect 9896 162134 13195 162136
rect 9896 162104 10376 162134
rect 13129 162131 13195 162134
rect 106877 161922 106943 161925
rect 106877 161920 109900 161922
rect 106877 161864 106882 161920
rect 106938 161864 109900 161920
rect 106877 161862 109900 161864
rect 106877 161859 106943 161862
rect 99057 161650 99123 161653
rect 183145 161650 183211 161653
rect 95732 161648 99123 161650
rect 95732 161592 99062 161648
rect 99118 161592 99123 161648
rect 95732 161590 99123 161592
rect 179820 161648 183211 161650
rect 179820 161592 183150 161648
rect 183206 161592 183211 161648
rect 179820 161590 183211 161592
rect 99057 161587 99123 161590
rect 183145 161587 183211 161590
rect 191977 160834 192043 160837
rect 191977 160832 193988 160834
rect 191977 160776 191982 160832
rect 192038 160776 193988 160832
rect 191977 160774 193988 160776
rect 191977 160771 192043 160774
rect 53333 160562 53399 160565
rect 137513 160562 137579 160565
rect 53333 160560 55988 160562
rect 53333 160504 53338 160560
rect 53394 160504 55988 160560
rect 53333 160502 55988 160504
rect 137513 160560 140076 160562
rect 137513 160504 137518 160560
rect 137574 160504 140076 160560
rect 137513 160502 140076 160504
rect 53333 160499 53399 160502
rect 137513 160499 137579 160502
rect 99149 160426 99215 160429
rect 183237 160426 183303 160429
rect 95732 160424 99215 160426
rect 95732 160368 99154 160424
rect 99210 160368 99215 160424
rect 95732 160366 99215 160368
rect 179820 160424 183303 160426
rect 179820 160368 183242 160424
rect 183298 160368 183303 160424
rect 179820 160366 183303 160368
rect 99149 160363 99215 160366
rect 183237 160363 183303 160366
rect 107245 159610 107311 159613
rect 107245 159608 109900 159610
rect 107245 159552 107250 159608
rect 107306 159552 109900 159608
rect 107245 159550 109900 159552
rect 107245 159547 107311 159550
rect 99425 159202 99491 159205
rect 183513 159202 183579 159205
rect 95732 159200 99491 159202
rect 95732 159144 99430 159200
rect 99486 159144 99491 159200
rect 95732 159142 99491 159144
rect 179820 159200 183579 159202
rect 179820 159144 183518 159200
rect 183574 159144 183579 159200
rect 179820 159142 183579 159144
rect 99425 159139 99491 159142
rect 183513 159139 183579 159142
rect 44501 158794 44567 158797
rect 41820 158792 44567 158794
rect 41820 158736 44506 158792
rect 44562 158736 44567 158792
rect 41820 158734 44567 158736
rect 44501 158731 44567 158734
rect 190045 158794 190111 158797
rect 190045 158792 193988 158794
rect 190045 158736 190050 158792
rect 190106 158736 193988 158792
rect 190045 158734 193988 158736
rect 190045 158731 190111 158734
rect 99241 157978 99307 157981
rect 183329 157978 183395 157981
rect 95732 157976 99307 157978
rect 95732 157920 99246 157976
rect 99302 157920 99307 157976
rect 95732 157918 99307 157920
rect 179820 157976 183395 157978
rect 179820 157920 183334 157976
rect 183390 157920 183395 157976
rect 179820 157918 183395 157920
rect 99241 157915 99307 157918
rect 183329 157915 183395 157918
rect 107153 157298 107219 157301
rect 107153 157296 109900 157298
rect 107153 157240 107158 157296
rect 107214 157240 109900 157296
rect 107153 157238 109900 157240
rect 107153 157235 107219 157238
rect 23617 157162 23683 157165
rect 212677 157162 212743 157165
rect 23617 157160 25996 157162
rect 23617 157104 23622 157160
rect 23678 157104 25996 157160
rect 209812 157160 212743 157162
rect 209812 157132 212682 157160
rect 23617 157102 25996 157104
rect 209782 157104 212682 157132
rect 212738 157104 212743 157160
rect 209782 157102 212743 157104
rect 23617 157099 23683 157102
rect 99333 156754 99399 156757
rect 95732 156752 99399 156754
rect 95732 156696 99338 156752
rect 99394 156696 99399 156752
rect 95732 156694 99399 156696
rect 99333 156691 99399 156694
rect 137513 156754 137579 156757
rect 138014 156754 138020 156756
rect 137513 156752 138020 156754
rect 137513 156696 137518 156752
rect 137574 156696 138020 156752
rect 137513 156694 138020 156696
rect 137513 156691 137579 156694
rect 138014 156692 138020 156694
rect 138084 156692 138090 156756
rect 183421 156754 183487 156757
rect 179820 156752 183487 156754
rect 179820 156696 183426 156752
rect 183482 156696 183487 156752
rect 179820 156694 183487 156696
rect 183421 156691 183487 156694
rect 189953 156754 190019 156757
rect 209782 156756 209842 157102
rect 212677 157099 212743 157102
rect 189953 156752 193988 156754
rect 189953 156696 189958 156752
rect 190014 156696 193988 156752
rect 189953 156694 193988 156696
rect 189953 156691 190019 156694
rect 209774 156692 209780 156756
rect 209844 156692 209850 156756
rect 99517 155530 99583 155533
rect 182777 155530 182843 155533
rect 95732 155528 99583 155530
rect 95732 155472 99522 155528
rect 99578 155472 99583 155528
rect 95732 155470 99583 155472
rect 179820 155528 182843 155530
rect 179820 155472 182782 155528
rect 182838 155472 182843 155528
rect 179820 155470 182843 155472
rect 99517 155467 99583 155470
rect 182777 155467 182843 155470
rect 106509 154986 106575 154989
rect 106509 154984 109900 154986
rect 106509 154928 106514 154984
rect 106570 154928 109900 154984
rect 106509 154926 109900 154928
rect 106509 154923 106575 154926
rect 191977 154850 192043 154853
rect 191977 154848 193988 154850
rect 191977 154792 191982 154848
rect 192038 154792 193988 154848
rect 191977 154790 193988 154792
rect 191977 154787 192043 154790
rect 98781 154442 98847 154445
rect 183605 154442 183671 154445
rect 95732 154440 98847 154442
rect 95732 154384 98786 154440
rect 98842 154384 98847 154440
rect 95732 154382 98847 154384
rect 179820 154440 183671 154442
rect 179820 154384 183610 154440
rect 183666 154384 183671 154440
rect 179820 154382 183671 154384
rect 98781 154379 98847 154382
rect 183605 154379 183671 154382
rect 222245 152946 222311 152949
rect 225416 152946 225896 152976
rect 222245 152944 225896 152946
rect 222245 152888 222250 152944
rect 222306 152888 225896 152944
rect 222245 152886 225896 152888
rect 222245 152883 222311 152886
rect 225416 152856 225896 152886
rect 134845 140570 134911 140573
rect 131796 140568 134911 140570
rect 47862 140434 47922 140540
rect 131796 140512 134850 140568
rect 134906 140512 134911 140568
rect 131796 140510 134911 140512
rect 134845 140507 134911 140510
rect 49929 140434 49995 140437
rect 47862 140432 49995 140434
rect 47862 140376 49934 140432
rect 49990 140376 49995 140432
rect 47862 140374 49995 140376
rect 49929 140371 49995 140374
rect 49929 140162 49995 140165
rect 47678 140160 49995 140162
rect 47678 140104 49934 140160
rect 49990 140104 49995 140160
rect 47678 140102 49995 140104
rect 47678 139996 47738 140102
rect 49929 140099 49995 140102
rect 100805 140162 100871 140165
rect 103982 140162 104042 140472
rect 100805 140160 104042 140162
rect 100805 140104 100810 140160
rect 100866 140104 104042 140160
rect 100805 140102 104042 140104
rect 184985 140162 185051 140165
rect 187886 140162 187946 140540
rect 184985 140160 187946 140162
rect 184985 140104 184990 140160
rect 185046 140104 187946 140160
rect 184985 140102 187946 140104
rect 100805 140099 100871 140102
rect 184985 140099 185051 140102
rect 100897 140026 100963 140029
rect 135397 140026 135463 140029
rect 100897 140024 104012 140026
rect 100897 139968 100902 140024
rect 100958 139968 104012 140024
rect 100897 139966 104012 139968
rect 131796 140024 135463 140026
rect 131796 139968 135402 140024
rect 135458 139968 135463 140024
rect 131796 139966 135463 139968
rect 100897 139963 100963 139966
rect 135397 139963 135463 139966
rect 185077 140026 185143 140029
rect 185077 140024 187762 140026
rect 185077 139968 185082 140024
rect 185138 139968 187762 140024
rect 185077 139966 187762 139968
rect 185077 139963 185143 139966
rect 187702 139890 187762 139966
rect 187886 139890 187946 139996
rect 187702 139830 187946 139890
rect 134661 139482 134727 139485
rect 131796 139480 134727 139482
rect 47862 139074 47922 139452
rect 131796 139424 134666 139480
rect 134722 139424 134727 139480
rect 131796 139422 134727 139424
rect 134661 139419 134727 139422
rect 49653 139074 49719 139077
rect 47862 139072 49719 139074
rect 47862 139016 49658 139072
rect 49714 139016 49719 139072
rect 47862 139014 49719 139016
rect 49653 139011 49719 139014
rect 58485 138938 58551 138941
rect 101173 138938 101239 138941
rect 103982 138938 104042 139384
rect 58485 138936 60986 138938
rect 47862 138802 47922 138908
rect 58485 138880 58490 138936
rect 58546 138880 60986 138936
rect 58485 138878 60986 138880
rect 58485 138875 58551 138878
rect 49929 138802 49995 138805
rect 47862 138800 49995 138802
rect 47862 138744 49934 138800
rect 49990 138744 49995 138800
rect 47862 138742 49995 138744
rect 49929 138739 49995 138742
rect 9896 138530 10376 138560
rect 13313 138530 13379 138533
rect 9896 138528 13379 138530
rect 9896 138472 13318 138528
rect 13374 138472 13379 138528
rect 9896 138470 13379 138472
rect 9896 138440 10376 138470
rect 13313 138467 13379 138470
rect 60926 138364 60986 138878
rect 101173 138936 104042 138938
rect 101173 138880 101178 138936
rect 101234 138880 104042 138936
rect 101173 138878 104042 138880
rect 185353 138938 185419 138941
rect 187886 138938 187946 139452
rect 185353 138936 187946 138938
rect 185353 138880 185358 138936
rect 185414 138880 187946 138936
rect 185353 138878 187946 138880
rect 101173 138875 101239 138878
rect 185353 138875 185419 138878
rect 101081 138802 101147 138805
rect 135397 138802 135463 138805
rect 101081 138800 104012 138802
rect 101081 138744 101086 138800
rect 101142 138744 104012 138800
rect 101081 138742 104012 138744
rect 131796 138800 135463 138802
rect 131796 138744 135402 138800
rect 135458 138744 135463 138800
rect 131796 138742 135463 138744
rect 101081 138739 101147 138742
rect 135397 138739 135463 138742
rect 185261 138666 185327 138669
rect 187886 138666 187946 138772
rect 185261 138664 187946 138666
rect 185261 138608 185266 138664
rect 185322 138608 187946 138664
rect 185261 138606 187946 138608
rect 185261 138603 185327 138606
rect 92709 138530 92775 138533
rect 90734 138528 92775 138530
rect 90734 138472 92714 138528
rect 92770 138472 92775 138528
rect 90734 138470 92775 138472
rect 90734 138432 90794 138470
rect 92709 138467 92775 138470
rect 143585 138530 143651 138533
rect 177717 138530 177783 138533
rect 143585 138528 145074 138530
rect 143585 138472 143590 138528
rect 143646 138472 145074 138528
rect 143585 138470 145074 138472
rect 143585 138467 143651 138470
rect 145014 138432 145074 138470
rect 174822 138528 177783 138530
rect 174822 138472 177722 138528
rect 177778 138472 177783 138528
rect 174822 138470 177783 138472
rect 174822 138364 174882 138470
rect 177717 138467 177783 138470
rect 58945 138258 59011 138261
rect 134661 138258 134727 138261
rect 58945 138256 60986 138258
rect 47862 137850 47922 138228
rect 58945 138200 58950 138256
rect 59006 138200 60986 138256
rect 58945 138198 60986 138200
rect 131796 138256 134727 138258
rect 131796 138200 134666 138256
rect 134722 138200 134727 138256
rect 131796 138198 134727 138200
rect 58945 138195 59011 138198
rect 50021 137850 50087 137853
rect 47862 137848 50087 137850
rect 47862 137792 50026 137848
rect 50082 137792 50087 137848
rect 60926 137820 60986 138198
rect 134661 138195 134727 138198
rect 143309 138258 143375 138261
rect 177625 138258 177691 138261
rect 143309 138256 145074 138258
rect 143309 138200 143314 138256
rect 143370 138200 145074 138256
rect 143309 138198 145074 138200
rect 143309 138195 143375 138198
rect 92801 138122 92867 138125
rect 90734 138120 92867 138122
rect 90734 138064 92806 138120
rect 92862 138064 92867 138120
rect 90734 138062 92867 138064
rect 90734 137888 90794 138062
rect 92801 138059 92867 138062
rect 101817 137850 101883 137853
rect 103982 137850 104042 138160
rect 145014 137888 145074 138198
rect 174822 138256 177691 138258
rect 174822 138200 177630 138256
rect 177686 138200 177691 138256
rect 174822 138198 177691 138200
rect 101817 137848 104042 137850
rect 47862 137790 50087 137792
rect 50021 137787 50087 137790
rect 101817 137792 101822 137848
rect 101878 137792 104042 137848
rect 174822 137820 174882 138198
rect 177625 138195 177691 138198
rect 185169 137850 185235 137853
rect 187886 137850 187946 138228
rect 185169 137848 187946 137850
rect 101817 137790 104042 137792
rect 185169 137792 185174 137848
rect 185230 137792 187946 137848
rect 185169 137790 187946 137792
rect 101817 137787 101883 137790
rect 185169 137787 185235 137790
rect 101265 137714 101331 137717
rect 135397 137714 135463 137717
rect 101265 137712 104012 137714
rect 47862 137442 47922 137684
rect 101265 137656 101270 137712
rect 101326 137656 104012 137712
rect 101265 137654 104012 137656
rect 131796 137712 135463 137714
rect 131796 137656 135402 137712
rect 135458 137656 135463 137712
rect 131796 137654 135463 137656
rect 101265 137651 101331 137654
rect 135397 137651 135463 137654
rect 49929 137442 49995 137445
rect 47862 137440 49995 137442
rect 47862 137384 49934 137440
rect 49990 137384 49995 137440
rect 47862 137382 49995 137384
rect 49929 137379 49995 137382
rect 185445 137306 185511 137309
rect 187886 137306 187946 137684
rect 185445 137304 187946 137306
rect 185445 137248 185450 137304
rect 185506 137248 187946 137304
rect 185445 137246 187946 137248
rect 185445 137243 185511 137246
rect 58393 137170 58459 137173
rect 92709 137170 92775 137173
rect 58393 137168 60956 137170
rect 47862 136762 47922 137140
rect 58393 137112 58398 137168
rect 58454 137112 60956 137168
rect 58393 137110 60956 137112
rect 90764 137168 92775 137170
rect 90764 137112 92714 137168
rect 92770 137112 92775 137168
rect 90764 137110 92775 137112
rect 58393 137107 58459 137110
rect 92709 137107 92775 137110
rect 143585 137170 143651 137173
rect 143585 137168 145044 137170
rect 143585 137112 143590 137168
rect 143646 137112 145044 137168
rect 143585 137110 145044 137112
rect 143585 137107 143651 137110
rect 135029 137034 135095 137037
rect 131796 137032 135095 137034
rect 131796 136976 135034 137032
rect 135090 136976 135095 137032
rect 131796 136974 135095 136976
rect 174822 137034 174882 137140
rect 177717 137034 177783 137037
rect 174822 137032 177783 137034
rect 174822 136976 177722 137032
rect 177778 136976 177783 137032
rect 174822 136974 177783 136976
rect 135029 136971 135095 136974
rect 177717 136971 177783 136974
rect 92801 136898 92867 136901
rect 90734 136896 92867 136898
rect 90734 136840 92806 136896
rect 92862 136840 92867 136896
rect 90734 136838 92867 136840
rect 51033 136762 51099 136765
rect 47862 136760 51099 136762
rect 47862 136704 51038 136760
rect 51094 136704 51099 136760
rect 47862 136702 51099 136704
rect 51033 136699 51099 136702
rect 90734 136664 90794 136838
rect 92801 136835 92867 136838
rect 58209 136626 58275 136629
rect 101173 136626 101239 136629
rect 103982 136626 104042 136936
rect 143125 136898 143191 136901
rect 177625 136898 177691 136901
rect 143125 136896 145074 136898
rect 143125 136840 143130 136896
rect 143186 136840 145074 136896
rect 143125 136838 145074 136840
rect 143125 136835 143191 136838
rect 145014 136664 145074 136838
rect 174822 136896 177691 136898
rect 174822 136840 177630 136896
rect 177686 136840 177691 136896
rect 174822 136838 177691 136840
rect 58209 136624 60956 136626
rect 47862 136218 47922 136596
rect 58209 136568 58214 136624
rect 58270 136568 60956 136624
rect 58209 136566 60956 136568
rect 101173 136624 104042 136626
rect 101173 136568 101178 136624
rect 101234 136568 104042 136624
rect 174822 136596 174882 136838
rect 177625 136835 177691 136838
rect 185169 136626 185235 136629
rect 187886 136626 187946 137004
rect 185169 136624 187946 136626
rect 101173 136566 104042 136568
rect 185169 136568 185174 136624
rect 185230 136568 187946 136624
rect 185169 136566 187946 136568
rect 58209 136563 58275 136566
rect 101173 136563 101239 136566
rect 185169 136563 185235 136566
rect 92709 136490 92775 136493
rect 135305 136490 135371 136493
rect 90734 136488 92775 136490
rect 90734 136432 92714 136488
rect 92770 136432 92775 136488
rect 90734 136430 92775 136432
rect 131796 136488 135371 136490
rect 131796 136432 135310 136488
rect 135366 136432 135371 136488
rect 131796 136430 135371 136432
rect 51125 136218 51191 136221
rect 47862 136216 51191 136218
rect 47862 136160 51130 136216
rect 51186 136160 51191 136216
rect 47862 136158 51191 136160
rect 51125 136155 51191 136158
rect 90734 136120 90794 136430
rect 92709 136427 92775 136430
rect 135305 136427 135371 136430
rect 58301 136082 58367 136085
rect 101265 136082 101331 136085
rect 103982 136082 104042 136392
rect 143493 136354 143559 136357
rect 177717 136354 177783 136357
rect 143493 136352 145074 136354
rect 143493 136296 143498 136352
rect 143554 136296 145074 136352
rect 143493 136294 145074 136296
rect 143493 136291 143559 136294
rect 145014 136120 145074 136294
rect 174822 136352 177783 136354
rect 174822 136296 177722 136352
rect 177778 136296 177783 136352
rect 174822 136294 177783 136296
rect 58301 136080 60956 136082
rect 47862 135946 47922 136052
rect 58301 136024 58306 136080
rect 58362 136024 60956 136080
rect 58301 136022 60956 136024
rect 101265 136080 104042 136082
rect 101265 136024 101270 136080
rect 101326 136024 104042 136080
rect 174822 136052 174882 136294
rect 177717 136291 177783 136294
rect 185261 136082 185327 136085
rect 187886 136082 187946 136460
rect 185261 136080 187946 136082
rect 101265 136022 104042 136024
rect 185261 136024 185266 136080
rect 185322 136024 187946 136080
rect 185261 136022 187946 136024
rect 58301 136019 58367 136022
rect 101265 136019 101331 136022
rect 185261 136019 185327 136022
rect 51217 135946 51283 135949
rect 47862 135944 51283 135946
rect 47862 135888 51222 135944
rect 51278 135888 51283 135944
rect 47862 135886 51283 135888
rect 51217 135883 51283 135886
rect 101725 135946 101791 135949
rect 135397 135946 135463 135949
rect 101725 135944 104012 135946
rect 101725 135888 101730 135944
rect 101786 135888 104012 135944
rect 101725 135886 104012 135888
rect 131796 135944 135463 135946
rect 131796 135888 135402 135944
rect 135458 135888 135463 135944
rect 131796 135886 135463 135888
rect 101725 135883 101791 135886
rect 135397 135883 135463 135886
rect 185353 135946 185419 135949
rect 215854 135946 215914 136188
rect 218381 135946 218447 135949
rect 185353 135944 187762 135946
rect 185353 135888 185358 135944
rect 185414 135888 187762 135944
rect 215854 135944 218447 135946
rect 185353 135886 187762 135888
rect 185353 135883 185419 135886
rect 143401 135810 143467 135813
rect 187702 135810 187762 135886
rect 187886 135810 187946 135916
rect 215854 135888 218386 135944
rect 218442 135888 218447 135944
rect 215854 135886 218447 135888
rect 218381 135883 218447 135886
rect 143401 135808 145074 135810
rect 143401 135752 143406 135808
rect 143462 135752 145074 135808
rect 143401 135750 145074 135752
rect 187702 135750 187946 135810
rect 143401 135747 143467 135750
rect 92709 135538 92775 135541
rect 90734 135536 92775 135538
rect 90734 135480 92714 135536
rect 92770 135480 92775 135536
rect 90734 135478 92775 135480
rect 90734 135440 90794 135478
rect 92709 135475 92775 135478
rect 145014 135440 145074 135750
rect 177717 135538 177783 135541
rect 174822 135536 177783 135538
rect 174822 135480 177722 135536
rect 177778 135480 177783 135536
rect 174822 135478 177783 135480
rect 58209 135402 58275 135405
rect 134845 135402 134911 135405
rect 58209 135400 60956 135402
rect 47862 134994 47922 135372
rect 58209 135344 58214 135400
rect 58270 135344 60956 135400
rect 58209 135342 60956 135344
rect 131796 135400 134911 135402
rect 131796 135344 134850 135400
rect 134906 135344 134911 135400
rect 174822 135372 174882 135478
rect 177717 135475 177783 135478
rect 131796 135342 134911 135344
rect 58209 135339 58275 135342
rect 134845 135339 134911 135342
rect 92801 135266 92867 135269
rect 90734 135264 92867 135266
rect 90734 135208 92806 135264
rect 92862 135208 92867 135264
rect 90734 135206 92867 135208
rect 51125 134994 51191 134997
rect 47862 134992 51191 134994
rect 47862 134936 51130 134992
rect 51186 134936 51191 134992
rect 47862 134934 51191 134936
rect 51125 134931 51191 134934
rect 90734 134896 90794 135206
rect 92801 135203 92867 135206
rect 58301 134858 58367 134861
rect 101817 134858 101883 134861
rect 103982 134858 104042 135304
rect 143309 135266 143375 135269
rect 177625 135266 177691 135269
rect 143309 135264 145074 135266
rect 143309 135208 143314 135264
rect 143370 135208 145074 135264
rect 143309 135206 145074 135208
rect 143309 135203 143375 135206
rect 145014 134896 145074 135206
rect 174822 135264 177691 135266
rect 174822 135208 177630 135264
rect 177686 135208 177691 135264
rect 174822 135206 177691 135208
rect 58301 134856 60956 134858
rect 47862 134722 47922 134828
rect 58301 134800 58306 134856
rect 58362 134800 60956 134856
rect 58301 134798 60956 134800
rect 101817 134856 104042 134858
rect 101817 134800 101822 134856
rect 101878 134800 104042 134856
rect 174822 134828 174882 135206
rect 177625 135203 177691 135206
rect 185169 134858 185235 134861
rect 187886 134858 187946 135372
rect 185169 134856 187946 134858
rect 101817 134798 104042 134800
rect 185169 134800 185174 134856
rect 185230 134800 187946 134856
rect 185169 134798 187946 134800
rect 58301 134795 58367 134798
rect 101817 134795 101883 134798
rect 185169 134795 185235 134798
rect 51217 134722 51283 134725
rect 134477 134722 134543 134725
rect 47862 134720 51283 134722
rect 47862 134664 51222 134720
rect 51278 134664 51283 134720
rect 47862 134662 51283 134664
rect 131796 134720 134543 134722
rect 131796 134664 134482 134720
rect 134538 134664 134543 134720
rect 131796 134662 134543 134664
rect 51217 134659 51283 134662
rect 134477 134659 134543 134662
rect 100897 134450 100963 134453
rect 103982 134450 104042 134624
rect 100897 134448 104042 134450
rect 100897 134392 100902 134448
rect 100958 134392 104042 134448
rect 100897 134390 104042 134392
rect 185077 134450 185143 134453
rect 187886 134450 187946 134692
rect 185077 134448 187946 134450
rect 185077 134392 185082 134448
rect 185138 134392 187946 134448
rect 185077 134390 187946 134392
rect 100897 134387 100963 134390
rect 185077 134387 185143 134390
rect 143585 134314 143651 134317
rect 177717 134314 177783 134317
rect 143585 134312 145074 134314
rect 47862 133906 47922 134284
rect 143585 134256 143590 134312
rect 143646 134256 145074 134312
rect 143585 134254 145074 134256
rect 143585 134251 143651 134254
rect 145014 134216 145074 134254
rect 174822 134312 177783 134314
rect 174822 134256 177722 134312
rect 177778 134256 177783 134312
rect 174822 134254 177783 134256
rect 58393 134178 58459 134181
rect 92709 134178 92775 134181
rect 135397 134178 135463 134181
rect 58393 134176 60956 134178
rect 58393 134120 58398 134176
rect 58454 134120 60956 134176
rect 58393 134118 60956 134120
rect 90764 134176 92775 134178
rect 90764 134120 92714 134176
rect 92770 134120 92775 134176
rect 90764 134118 92775 134120
rect 131796 134176 135463 134178
rect 131796 134120 135402 134176
rect 135458 134120 135463 134176
rect 174822 134148 174882 134254
rect 177717 134251 177783 134254
rect 131796 134118 135463 134120
rect 58393 134115 58459 134118
rect 92709 134115 92775 134118
rect 135397 134115 135463 134118
rect 92801 134042 92867 134045
rect 90734 134040 92867 134042
rect 90734 133984 92806 134040
rect 92862 133984 92867 134040
rect 90734 133982 92867 133984
rect 50389 133906 50455 133909
rect 47862 133904 50455 133906
rect 18097 133362 18163 133365
rect 19894 133362 19954 133876
rect 47862 133848 50394 133904
rect 50450 133848 50455 133904
rect 47862 133846 50455 133848
rect 50389 133843 50455 133846
rect 18097 133360 19954 133362
rect 18097 133304 18102 133360
rect 18158 133304 19954 133360
rect 18097 133302 19954 133304
rect 47862 133362 47922 133740
rect 90734 133672 90794 133982
rect 92801 133979 92867 133982
rect 101357 133770 101423 133773
rect 103982 133770 104042 134080
rect 143217 134042 143283 134045
rect 143217 134040 145074 134042
rect 143217 133984 143222 134040
rect 143278 133984 145074 134040
rect 143217 133982 145074 133984
rect 143217 133979 143283 133982
rect 101357 133768 104042 133770
rect 101357 133712 101362 133768
rect 101418 133712 104042 133768
rect 101357 133710 104042 133712
rect 101357 133707 101423 133710
rect 145014 133672 145074 133982
rect 177717 133906 177783 133909
rect 174822 133904 177783 133906
rect 174822 133848 177722 133904
rect 177778 133848 177783 133904
rect 174822 133846 177783 133848
rect 58209 133634 58275 133637
rect 135029 133634 135095 133637
rect 58209 133632 60956 133634
rect 58209 133576 58214 133632
rect 58270 133576 60956 133632
rect 58209 133574 60956 133576
rect 131796 133632 135095 133634
rect 131796 133576 135034 133632
rect 135090 133576 135095 133632
rect 174822 133604 174882 133846
rect 177717 133843 177783 133846
rect 185169 133770 185235 133773
rect 187886 133770 187946 134148
rect 185169 133768 187946 133770
rect 185169 133712 185174 133768
rect 185230 133712 187946 133768
rect 185169 133710 187946 133712
rect 185169 133707 185235 133710
rect 131796 133574 135095 133576
rect 58209 133571 58275 133574
rect 135029 133571 135095 133574
rect 92893 133498 92959 133501
rect 90734 133496 92959 133498
rect 90734 133440 92898 133496
rect 92954 133440 92959 133496
rect 90734 133438 92959 133440
rect 51125 133362 51191 133365
rect 47862 133360 51191 133362
rect 47862 133304 51130 133360
rect 51186 133304 51191 133360
rect 47862 133302 51191 133304
rect 18097 133299 18163 133302
rect 51125 133299 51191 133302
rect 47862 133090 47922 133196
rect 90734 133128 90794 133438
rect 92893 133435 92959 133438
rect 51217 133090 51283 133093
rect 47862 133088 51283 133090
rect 47862 133032 51222 133088
rect 51278 133032 51283 133088
rect 47862 133030 51283 133032
rect 51217 133027 51283 133030
rect 58301 133090 58367 133093
rect 101725 133090 101791 133093
rect 103982 133090 104042 133536
rect 177625 133498 177691 133501
rect 174822 133496 177691 133498
rect 174822 133440 177630 133496
rect 177686 133440 177691 133496
rect 174822 133438 177691 133440
rect 142941 133362 143007 133365
rect 142941 133360 145074 133362
rect 142941 133304 142946 133360
rect 143002 133304 145074 133360
rect 142941 133302 145074 133304
rect 142941 133299 143007 133302
rect 145014 133128 145074 133302
rect 58301 133088 60956 133090
rect 58301 133032 58306 133088
rect 58362 133032 60956 133088
rect 58301 133030 60956 133032
rect 101725 133088 104042 133090
rect 101725 133032 101730 133088
rect 101786 133032 104042 133088
rect 174822 133060 174882 133438
rect 177625 133435 177691 133438
rect 185813 133090 185879 133093
rect 187886 133090 187946 133604
rect 185813 133088 187946 133090
rect 101725 133030 104042 133032
rect 185813 133032 185818 133088
rect 185874 133032 187946 133088
rect 185813 133030 187946 133032
rect 58301 133027 58367 133030
rect 101725 133027 101791 133030
rect 185813 133027 185879 133030
rect 135305 132954 135371 132957
rect 131796 132952 135371 132954
rect 131796 132896 135310 132952
rect 135366 132896 135371 132952
rect 131796 132894 135371 132896
rect 135305 132891 135371 132894
rect 92709 132682 92775 132685
rect 90734 132680 92775 132682
rect 90734 132624 92714 132680
rect 92770 132624 92775 132680
rect 90734 132622 92775 132624
rect 47862 132138 47922 132516
rect 90734 132448 90794 132622
rect 92709 132619 92775 132622
rect 101817 132546 101883 132549
rect 103982 132546 104042 132856
rect 143585 132818 143651 132821
rect 143585 132816 145074 132818
rect 143585 132760 143590 132816
rect 143646 132760 145074 132816
rect 143585 132758 145074 132760
rect 143585 132755 143651 132758
rect 101817 132544 104042 132546
rect 101817 132488 101822 132544
rect 101878 132488 104042 132544
rect 101817 132486 104042 132488
rect 101817 132483 101883 132486
rect 145014 132448 145074 132758
rect 177717 132682 177783 132685
rect 174822 132680 177783 132682
rect 174822 132624 177722 132680
rect 177778 132624 177783 132680
rect 174822 132622 177783 132624
rect 58301 132410 58367 132413
rect 135397 132410 135463 132413
rect 58301 132408 60956 132410
rect 58301 132352 58306 132408
rect 58362 132352 60956 132408
rect 58301 132350 60956 132352
rect 131796 132408 135463 132410
rect 131796 132352 135402 132408
rect 135458 132352 135463 132408
rect 174822 132380 174882 132622
rect 177717 132619 177783 132622
rect 185445 132546 185511 132549
rect 187886 132546 187946 132924
rect 185445 132544 187946 132546
rect 185445 132488 185450 132544
rect 185506 132488 187946 132544
rect 185445 132486 187946 132488
rect 185445 132483 185511 132486
rect 131796 132350 135463 132352
rect 58301 132347 58367 132350
rect 135397 132347 135463 132350
rect 92801 132274 92867 132277
rect 90734 132272 92867 132274
rect 90734 132216 92806 132272
rect 92862 132216 92867 132272
rect 90734 132214 92867 132216
rect 51125 132138 51191 132141
rect 47862 132136 51191 132138
rect 47862 132080 51130 132136
rect 51186 132080 51191 132136
rect 47862 132078 51191 132080
rect 51125 132075 51191 132078
rect 47862 131866 47922 131972
rect 90734 131904 90794 132214
rect 92801 132211 92867 132214
rect 101449 132002 101515 132005
rect 103982 132002 104042 132312
rect 143217 132274 143283 132277
rect 177625 132274 177691 132277
rect 143217 132272 145074 132274
rect 143217 132216 143222 132272
rect 143278 132216 145074 132272
rect 143217 132214 145074 132216
rect 143217 132211 143283 132214
rect 101449 132000 104042 132002
rect 101449 131944 101454 132000
rect 101510 131944 104042 132000
rect 101449 131942 104042 131944
rect 101449 131939 101515 131942
rect 145014 131904 145074 132214
rect 174822 132272 177691 132274
rect 174822 132216 177630 132272
rect 177686 132216 177691 132272
rect 174822 132214 177691 132216
rect 51217 131866 51283 131869
rect 47862 131864 51283 131866
rect 47862 131808 51222 131864
rect 51278 131808 51283 131864
rect 47862 131806 51283 131808
rect 51217 131803 51283 131806
rect 58209 131866 58275 131869
rect 101633 131866 101699 131869
rect 135029 131866 135095 131869
rect 58209 131864 60956 131866
rect 58209 131808 58214 131864
rect 58270 131808 60956 131864
rect 58209 131806 60956 131808
rect 101633 131864 104012 131866
rect 101633 131808 101638 131864
rect 101694 131808 104012 131864
rect 101633 131806 104012 131808
rect 131796 131864 135095 131866
rect 131796 131808 135034 131864
rect 135090 131808 135095 131864
rect 174822 131836 174882 132214
rect 177625 132211 177691 132214
rect 185721 132002 185787 132005
rect 187886 132002 187946 132380
rect 185721 132000 187946 132002
rect 185721 131944 185726 132000
rect 185782 131944 187946 132000
rect 185721 131942 187946 131944
rect 185721 131939 185787 131942
rect 131796 131806 135095 131808
rect 58209 131803 58275 131806
rect 101633 131803 101699 131806
rect 135029 131803 135095 131806
rect 185537 131730 185603 131733
rect 187886 131730 187946 131836
rect 185537 131728 187946 131730
rect 185537 131672 185542 131728
rect 185598 131672 187946 131728
rect 185537 131670 187946 131672
rect 185537 131667 185603 131670
rect 143585 131458 143651 131461
rect 143585 131456 145074 131458
rect 47862 131050 47922 131428
rect 143585 131400 143590 131456
rect 143646 131400 145074 131456
rect 143585 131398 145074 131400
rect 143585 131395 143651 131398
rect 92709 131322 92775 131325
rect 135029 131322 135095 131325
rect 90734 131320 92775 131322
rect 90734 131264 92714 131320
rect 92770 131264 92775 131320
rect 90734 131262 92775 131264
rect 131796 131320 135095 131322
rect 131796 131264 135034 131320
rect 135090 131264 135095 131320
rect 131796 131262 135095 131264
rect 90734 131224 90794 131262
rect 92709 131259 92775 131262
rect 135029 131259 135095 131262
rect 145014 131224 145074 131398
rect 177717 131322 177783 131325
rect 174822 131320 177783 131322
rect 174822 131264 177722 131320
rect 177778 131264 177783 131320
rect 174822 131262 177783 131264
rect 58209 131186 58275 131189
rect 58209 131184 60956 131186
rect 58209 131128 58214 131184
rect 58270 131128 60956 131184
rect 58209 131126 60956 131128
rect 58209 131123 58275 131126
rect 50205 131050 50271 131053
rect 92801 131050 92867 131053
rect 47862 131048 50271 131050
rect 47862 130992 50210 131048
rect 50266 130992 50271 131048
rect 47862 130990 50271 130992
rect 50205 130987 50271 130990
rect 90734 131048 92867 131050
rect 90734 130992 92806 131048
rect 92862 130992 92867 131048
rect 90734 130990 92867 130992
rect 47862 130642 47922 130884
rect 90734 130680 90794 130990
rect 92801 130987 92867 130990
rect 101725 130778 101791 130781
rect 103982 130778 104042 131224
rect 174822 131156 174882 131262
rect 177717 131259 177783 131262
rect 142481 131050 142547 131053
rect 177625 131050 177691 131053
rect 142481 131048 145074 131050
rect 142481 130992 142486 131048
rect 142542 130992 145074 131048
rect 142481 130990 145074 130992
rect 142481 130987 142547 130990
rect 101725 130776 104042 130778
rect 101725 130720 101730 130776
rect 101786 130720 104042 130776
rect 101725 130718 104042 130720
rect 101725 130715 101791 130718
rect 145014 130680 145074 130990
rect 174822 131048 177691 131050
rect 174822 130992 177630 131048
rect 177686 130992 177691 131048
rect 174822 130990 177691 130992
rect 51125 130642 51191 130645
rect 47862 130640 51191 130642
rect 47862 130584 51130 130640
rect 51186 130584 51191 130640
rect 47862 130582 51191 130584
rect 51125 130579 51191 130582
rect 58301 130642 58367 130645
rect 135397 130642 135463 130645
rect 58301 130640 60956 130642
rect 58301 130584 58306 130640
rect 58362 130584 60956 130640
rect 58301 130582 60956 130584
rect 131796 130640 135463 130642
rect 131796 130584 135402 130640
rect 135458 130584 135463 130640
rect 174822 130612 174882 130990
rect 177625 130987 177691 130990
rect 185261 130778 185327 130781
rect 187886 130778 187946 131292
rect 185261 130776 187946 130778
rect 185261 130720 185266 130776
rect 185322 130720 187946 130776
rect 185261 130718 187946 130720
rect 185261 130715 185327 130718
rect 131796 130582 135463 130584
rect 58301 130579 58367 130582
rect 135397 130579 135463 130582
rect 51217 130506 51283 130509
rect 47678 130504 51283 130506
rect 47678 130448 51222 130504
rect 51278 130448 51283 130504
rect 47678 130446 51283 130448
rect 47678 130340 47738 130446
rect 51217 130443 51283 130446
rect 101817 130370 101883 130373
rect 103982 130370 104042 130544
rect 101817 130368 104042 130370
rect 101817 130312 101822 130368
rect 101878 130312 104042 130368
rect 101817 130310 104042 130312
rect 185353 130370 185419 130373
rect 187886 130370 187946 130612
rect 185353 130368 187946 130370
rect 185353 130312 185358 130368
rect 185414 130312 187946 130368
rect 185353 130310 187946 130312
rect 101817 130307 101883 130310
rect 185353 130307 185419 130310
rect 143585 130234 143651 130237
rect 177717 130234 177783 130237
rect 143585 130232 145074 130234
rect 143585 130176 143590 130232
rect 143646 130176 145074 130232
rect 143585 130174 145074 130176
rect 143585 130171 143651 130174
rect 145014 130136 145074 130174
rect 174822 130232 177783 130234
rect 174822 130176 177722 130232
rect 177778 130176 177783 130232
rect 174822 130174 177783 130176
rect 58485 130098 58551 130101
rect 92709 130098 92775 130101
rect 135397 130098 135463 130101
rect 58485 130096 60956 130098
rect 58485 130040 58490 130096
rect 58546 130040 60956 130096
rect 58485 130038 60956 130040
rect 90764 130096 92775 130098
rect 90764 130040 92714 130096
rect 92770 130040 92775 130096
rect 90764 130038 92775 130040
rect 131796 130096 135463 130098
rect 131796 130040 135402 130096
rect 135458 130040 135463 130096
rect 174822 130068 174882 130174
rect 177717 130171 177783 130174
rect 131796 130038 135463 130040
rect 58485 130035 58551 130038
rect 92709 130035 92775 130038
rect 135397 130035 135463 130038
rect 92801 129826 92867 129829
rect 90734 129824 92867 129826
rect 90734 129768 92806 129824
rect 92862 129768 92867 129824
rect 90734 129766 92867 129768
rect 47862 129282 47922 129660
rect 90734 129456 90794 129766
rect 92801 129763 92867 129766
rect 101357 129690 101423 129693
rect 103982 129690 104042 130000
rect 143033 129962 143099 129965
rect 143033 129960 145074 129962
rect 143033 129904 143038 129960
rect 143094 129904 145074 129960
rect 143033 129902 145074 129904
rect 143033 129899 143099 129902
rect 101357 129688 104042 129690
rect 101357 129632 101362 129688
rect 101418 129632 104042 129688
rect 101357 129630 104042 129632
rect 101357 129627 101423 129630
rect 135305 129554 135371 129557
rect 131796 129552 135371 129554
rect 131796 129496 135310 129552
rect 135366 129496 135371 129552
rect 131796 129494 135371 129496
rect 135305 129491 135371 129494
rect 145014 129456 145074 129902
rect 177625 129826 177691 129829
rect 174822 129824 177691 129826
rect 174822 129768 177630 129824
rect 177686 129768 177691 129824
rect 174822 129766 177691 129768
rect 58209 129418 58275 129421
rect 58209 129416 60956 129418
rect 58209 129360 58214 129416
rect 58270 129360 60956 129416
rect 58209 129358 60956 129360
rect 58209 129355 58275 129358
rect 51125 129282 51191 129285
rect 47862 129280 51191 129282
rect 47862 129224 51130 129280
rect 51186 129224 51191 129280
rect 47862 129222 51191 129224
rect 51125 129219 51191 129222
rect 47862 129010 47922 129116
rect 51217 129010 51283 129013
rect 47862 129008 51283 129010
rect 47862 128952 51222 129008
rect 51278 128952 51283 129008
rect 47862 128950 51283 128952
rect 51217 128947 51283 128950
rect 101265 129010 101331 129013
rect 103982 129010 104042 129456
rect 174822 129388 174882 129766
rect 177625 129763 177691 129766
rect 185169 129690 185235 129693
rect 187886 129690 187946 130068
rect 185169 129688 187946 129690
rect 185169 129632 185174 129688
rect 185230 129632 187946 129688
rect 185169 129630 187946 129632
rect 185169 129627 185235 129630
rect 101265 129008 104042 129010
rect 101265 128952 101270 129008
rect 101326 128952 104042 129008
rect 101265 128950 104042 128952
rect 185445 129010 185511 129013
rect 187886 129010 187946 129524
rect 185445 129008 187946 129010
rect 185445 128952 185450 129008
rect 185506 128952 187946 129008
rect 185445 128950 187946 128952
rect 101265 128947 101331 128950
rect 185445 128947 185511 128950
rect 58209 128874 58275 128877
rect 92709 128874 92775 128877
rect 135397 128874 135463 128877
rect 58209 128872 60956 128874
rect 58209 128816 58214 128872
rect 58270 128816 60956 128872
rect 58209 128814 60956 128816
rect 90764 128872 92775 128874
rect 90764 128816 92714 128872
rect 92770 128816 92775 128872
rect 90764 128814 92775 128816
rect 131796 128872 135463 128874
rect 131796 128816 135402 128872
rect 135458 128816 135463 128872
rect 131796 128814 135463 128816
rect 58209 128811 58275 128814
rect 92709 128811 92775 128814
rect 135397 128811 135463 128814
rect 142757 128874 142823 128877
rect 142757 128872 145044 128874
rect 142757 128816 142762 128872
rect 142818 128816 145044 128872
rect 142757 128814 145044 128816
rect 142757 128811 142823 128814
rect 47862 128194 47922 128572
rect 92801 128466 92867 128469
rect 90734 128464 92867 128466
rect 90734 128408 92806 128464
rect 92862 128408 92867 128464
rect 90734 128406 92867 128408
rect 90734 128232 90794 128406
rect 92801 128403 92867 128406
rect 100989 128466 101055 128469
rect 103982 128466 104042 128776
rect 143585 128738 143651 128741
rect 174822 128738 174882 128844
rect 177717 128738 177783 128741
rect 143585 128736 145074 128738
rect 143585 128680 143590 128736
rect 143646 128680 145074 128736
rect 143585 128678 145074 128680
rect 174822 128736 177783 128738
rect 174822 128680 177722 128736
rect 177778 128680 177783 128736
rect 174822 128678 177783 128680
rect 143585 128675 143651 128678
rect 100989 128464 104042 128466
rect 100989 128408 100994 128464
rect 101050 128408 104042 128464
rect 100989 128406 104042 128408
rect 100989 128403 101055 128406
rect 134661 128330 134727 128333
rect 131796 128328 134727 128330
rect 131796 128272 134666 128328
rect 134722 128272 134727 128328
rect 131796 128270 134727 128272
rect 134661 128267 134727 128270
rect 145014 128232 145074 128678
rect 177717 128675 177783 128678
rect 177625 128466 177691 128469
rect 174822 128464 177691 128466
rect 174822 128408 177630 128464
rect 177686 128408 177691 128464
rect 174822 128406 177691 128408
rect 50757 128194 50823 128197
rect 47862 128192 50823 128194
rect 47862 128136 50762 128192
rect 50818 128136 50823 128192
rect 47862 128134 50823 128136
rect 50757 128131 50823 128134
rect 58393 128194 58459 128197
rect 58393 128192 60956 128194
rect 58393 128136 58398 128192
rect 58454 128136 60956 128192
rect 58393 128134 60956 128136
rect 58393 128131 58459 128134
rect 92893 128058 92959 128061
rect 90734 128056 92959 128058
rect 47862 127786 47922 128028
rect 90734 128000 92898 128056
rect 92954 128000 92959 128056
rect 90734 127998 92959 128000
rect 51217 127786 51283 127789
rect 47862 127784 51283 127786
rect 47862 127728 51222 127784
rect 51278 127728 51283 127784
rect 47862 127726 51283 127728
rect 51217 127723 51283 127726
rect 90734 127688 90794 127998
rect 92893 127995 92959 127998
rect 101173 127922 101239 127925
rect 103982 127922 104042 128232
rect 174822 128164 174882 128406
rect 177625 128403 177691 128406
rect 185169 128466 185235 128469
rect 187886 128466 187946 128844
rect 185169 128464 187946 128466
rect 185169 128408 185174 128464
rect 185230 128408 187946 128464
rect 185169 128406 187946 128408
rect 185169 128403 185235 128406
rect 143125 128058 143191 128061
rect 177809 128058 177875 128061
rect 143125 128056 145074 128058
rect 143125 128000 143130 128056
rect 143186 128000 145074 128056
rect 143125 127998 145074 128000
rect 143125 127995 143191 127998
rect 101173 127920 104042 127922
rect 101173 127864 101178 127920
rect 101234 127864 104042 127920
rect 101173 127862 104042 127864
rect 101173 127859 101239 127862
rect 101081 127786 101147 127789
rect 135305 127786 135371 127789
rect 101081 127784 104012 127786
rect 101081 127728 101086 127784
rect 101142 127728 104012 127784
rect 101081 127726 104012 127728
rect 131796 127784 135371 127786
rect 131796 127728 135310 127784
rect 135366 127728 135371 127784
rect 131796 127726 135371 127728
rect 101081 127723 101147 127726
rect 135305 127723 135371 127726
rect 145014 127688 145074 127998
rect 174822 128056 177875 128058
rect 174822 128000 177814 128056
rect 177870 128000 177875 128056
rect 174822 127998 177875 128000
rect 58301 127650 58367 127653
rect 58301 127648 60956 127650
rect 58301 127592 58306 127648
rect 58362 127592 60956 127648
rect 174822 127620 174882 127998
rect 177809 127995 177875 127998
rect 185353 127922 185419 127925
rect 187886 127922 187946 128300
rect 185353 127920 187946 127922
rect 185353 127864 185358 127920
rect 185414 127864 187946 127920
rect 185353 127862 187946 127864
rect 185353 127859 185419 127862
rect 185261 127650 185327 127653
rect 187886 127650 187946 127756
rect 185261 127648 187946 127650
rect 58301 127590 60956 127592
rect 185261 127592 185266 127648
rect 185322 127592 187946 127648
rect 185261 127590 187946 127592
rect 58301 127587 58367 127590
rect 185261 127587 185327 127590
rect 47862 126970 47922 127484
rect 142481 127378 142547 127381
rect 217001 127378 217067 127381
rect 142481 127376 145074 127378
rect 142481 127320 142486 127376
rect 142542 127320 145074 127376
rect 142481 127318 145074 127320
rect 142481 127315 142547 127318
rect 92709 127242 92775 127245
rect 135397 127242 135463 127245
rect 90734 127240 92775 127242
rect 90734 127184 92714 127240
rect 92770 127184 92775 127240
rect 90734 127182 92775 127184
rect 131796 127240 135463 127242
rect 131796 127184 135402 127240
rect 135458 127184 135463 127240
rect 131796 127182 135463 127184
rect 90734 127144 90794 127182
rect 92709 127179 92775 127182
rect 135397 127179 135463 127182
rect 145014 127144 145074 127318
rect 215670 127376 217067 127378
rect 215670 127320 217006 127376
rect 217062 127320 217067 127376
rect 215670 127318 217067 127320
rect 177165 127242 177231 127245
rect 174822 127240 177231 127242
rect 174822 127184 177170 127240
rect 177226 127184 177231 127240
rect 174822 127182 177231 127184
rect 58393 127106 58459 127109
rect 58393 127104 60956 127106
rect 58393 127048 58398 127104
rect 58454 127048 60956 127104
rect 58393 127046 60956 127048
rect 58393 127043 58459 127046
rect 50205 126970 50271 126973
rect 92801 126970 92867 126973
rect 47862 126968 50271 126970
rect 47862 126912 50210 126968
rect 50266 126912 50271 126968
rect 47862 126910 50271 126912
rect 50205 126907 50271 126910
rect 90734 126968 92867 126970
rect 90734 126912 92806 126968
rect 92862 126912 92867 126968
rect 90734 126910 92867 126912
rect 47862 126562 47922 126804
rect 50389 126562 50455 126565
rect 47862 126560 50455 126562
rect 47862 126504 50394 126560
rect 50450 126504 50455 126560
rect 47862 126502 50455 126504
rect 50389 126499 50455 126502
rect 90734 126464 90794 126910
rect 92801 126907 92867 126910
rect 101265 126698 101331 126701
rect 103982 126698 104042 127144
rect 174822 127076 174882 127182
rect 177165 127179 177231 127182
rect 143309 126970 143375 126973
rect 177717 126970 177783 126973
rect 143309 126968 145074 126970
rect 143309 126912 143314 126968
rect 143370 126912 145074 126968
rect 143309 126910 145074 126912
rect 143309 126907 143375 126910
rect 101265 126696 104042 126698
rect 101265 126640 101270 126696
rect 101326 126640 104042 126696
rect 101265 126638 104042 126640
rect 101265 126635 101331 126638
rect 135397 126562 135463 126565
rect 131796 126560 135463 126562
rect 131796 126504 135402 126560
rect 135458 126504 135463 126560
rect 131796 126502 135463 126504
rect 135397 126499 135463 126502
rect 145014 126464 145074 126910
rect 174822 126968 177783 126970
rect 174822 126912 177722 126968
rect 177778 126912 177783 126968
rect 174822 126910 177783 126912
rect 58209 126426 58275 126429
rect 58209 126424 60956 126426
rect 58209 126368 58214 126424
rect 58270 126368 60956 126424
rect 58209 126366 60956 126368
rect 58209 126363 58275 126366
rect 100989 126290 101055 126293
rect 103982 126290 104042 126464
rect 174822 126396 174882 126910
rect 177717 126907 177783 126910
rect 185445 126698 185511 126701
rect 187886 126698 187946 127212
rect 215670 126804 215730 127318
rect 217001 127315 217067 127318
rect 222337 126834 222403 126837
rect 225416 126834 225896 126864
rect 222337 126832 225896 126834
rect 222337 126776 222342 126832
rect 222398 126776 225896 126832
rect 222337 126774 225896 126776
rect 222337 126771 222403 126774
rect 225416 126744 225896 126774
rect 185445 126696 187946 126698
rect 185445 126640 185450 126696
rect 185506 126640 187946 126696
rect 185445 126638 187946 126640
rect 185445 126635 185511 126638
rect 100989 126288 104042 126290
rect 47862 126154 47922 126260
rect 100989 126232 100994 126288
rect 101050 126232 104042 126288
rect 100989 126230 104042 126232
rect 185169 126290 185235 126293
rect 187886 126290 187946 126532
rect 185169 126288 187946 126290
rect 185169 126232 185174 126288
rect 185230 126232 187946 126288
rect 185169 126230 187946 126232
rect 100989 126227 101055 126230
rect 185169 126227 185235 126230
rect 51217 126154 51283 126157
rect 47862 126152 51283 126154
rect 47862 126096 51222 126152
rect 51278 126096 51283 126152
rect 47862 126094 51283 126096
rect 51217 126091 51283 126094
rect 92709 126018 92775 126021
rect 135213 126018 135279 126021
rect 90734 126016 92775 126018
rect 90734 125960 92714 126016
rect 92770 125960 92775 126016
rect 90734 125958 92775 125960
rect 131796 126016 135279 126018
rect 131796 125960 135218 126016
rect 135274 125960 135279 126016
rect 131796 125958 135279 125960
rect 90734 125920 90794 125958
rect 92709 125955 92775 125958
rect 135213 125955 135279 125958
rect 143585 126018 143651 126021
rect 177717 126018 177783 126021
rect 143585 126016 145074 126018
rect 143585 125960 143590 126016
rect 143646 125960 145074 126016
rect 143585 125958 145074 125960
rect 143585 125955 143651 125958
rect 145014 125920 145074 125958
rect 174822 126016 177783 126018
rect 174822 125960 177722 126016
rect 177778 125960 177783 126016
rect 174822 125958 177783 125960
rect 58301 125882 58367 125885
rect 58301 125880 60956 125882
rect 58301 125824 58306 125880
rect 58362 125824 60956 125880
rect 58301 125822 60956 125824
rect 58301 125819 58367 125822
rect 47862 125338 47922 125716
rect 92801 125610 92867 125613
rect 90734 125608 92867 125610
rect 90734 125552 92806 125608
rect 92862 125552 92867 125608
rect 90734 125550 92867 125552
rect 51125 125338 51191 125341
rect 47862 125336 51191 125338
rect 47862 125280 51130 125336
rect 51186 125280 51191 125336
rect 47862 125278 51191 125280
rect 51125 125275 51191 125278
rect 90734 125240 90794 125550
rect 92801 125547 92867 125550
rect 100989 125610 101055 125613
rect 103982 125610 104042 125920
rect 174822 125852 174882 125958
rect 177717 125955 177783 125958
rect 100989 125608 104042 125610
rect 100989 125552 100994 125608
rect 101050 125552 104042 125608
rect 100989 125550 104042 125552
rect 143493 125610 143559 125613
rect 177625 125610 177691 125613
rect 143493 125608 145074 125610
rect 143493 125552 143498 125608
rect 143554 125552 145074 125608
rect 143493 125550 145074 125552
rect 100989 125547 101055 125550
rect 143493 125547 143559 125550
rect 135397 125474 135463 125477
rect 131796 125472 135463 125474
rect 131796 125416 135402 125472
rect 135458 125416 135463 125472
rect 131796 125414 135463 125416
rect 135397 125411 135463 125414
rect 58209 125202 58275 125205
rect 58209 125200 60956 125202
rect 47862 125066 47922 125172
rect 58209 125144 58214 125200
rect 58270 125144 60956 125200
rect 58209 125142 60956 125144
rect 58209 125139 58275 125142
rect 51217 125066 51283 125069
rect 47862 125064 51283 125066
rect 47862 125008 51222 125064
rect 51278 125008 51283 125064
rect 47862 125006 51283 125008
rect 51217 125003 51283 125006
rect 101265 125066 101331 125069
rect 103982 125066 104042 125376
rect 145014 125240 145074 125550
rect 174822 125608 177691 125610
rect 174822 125552 177630 125608
rect 177686 125552 177691 125608
rect 174822 125550 177691 125552
rect 174822 125172 174882 125550
rect 177625 125547 177691 125550
rect 185169 125610 185235 125613
rect 187886 125610 187946 125988
rect 185169 125608 187946 125610
rect 185169 125552 185174 125608
rect 185230 125552 187946 125608
rect 185169 125550 187946 125552
rect 185169 125547 185235 125550
rect 101265 125064 104042 125066
rect 101265 125008 101270 125064
rect 101326 125008 104042 125064
rect 101265 125006 104042 125008
rect 101265 125003 101331 125006
rect 185445 124930 185511 124933
rect 187886 124930 187946 125444
rect 185445 124928 187946 124930
rect 185445 124872 185450 124928
rect 185506 124872 187946 124928
rect 185445 124870 187946 124872
rect 185445 124867 185511 124870
rect 101081 124794 101147 124797
rect 135397 124794 135463 124797
rect 101081 124792 104012 124794
rect 101081 124736 101086 124792
rect 101142 124736 104012 124792
rect 101081 124734 104012 124736
rect 131796 124792 135463 124794
rect 131796 124736 135402 124792
rect 135458 124736 135463 124792
rect 131796 124734 135463 124736
rect 101081 124731 101147 124734
rect 135397 124731 135463 124734
rect 185353 124794 185419 124797
rect 185353 124792 187762 124794
rect 185353 124736 185358 124792
rect 185414 124736 187762 124792
rect 185353 124734 187762 124736
rect 185353 124731 185419 124734
rect 58301 124658 58367 124661
rect 92709 124658 92775 124661
rect 58301 124656 60956 124658
rect 47862 124114 47922 124628
rect 58301 124600 58306 124656
rect 58362 124600 60956 124656
rect 58301 124598 60956 124600
rect 90764 124656 92775 124658
rect 90764 124600 92714 124656
rect 92770 124600 92775 124656
rect 90764 124598 92775 124600
rect 58301 124595 58367 124598
rect 92709 124595 92775 124598
rect 143585 124658 143651 124661
rect 187702 124658 187762 124734
rect 187886 124658 187946 124764
rect 143585 124656 145044 124658
rect 143585 124600 143590 124656
rect 143646 124600 145044 124656
rect 143585 124598 145044 124600
rect 143585 124595 143651 124598
rect 174822 124522 174882 124628
rect 187702 124598 187946 124658
rect 177717 124522 177783 124525
rect 174822 124520 177783 124522
rect 174822 124464 177722 124520
rect 177778 124464 177783 124520
rect 174822 124462 177783 124464
rect 177717 124459 177783 124462
rect 92801 124386 92867 124389
rect 90734 124384 92867 124386
rect 90734 124328 92806 124384
rect 92862 124328 92867 124384
rect 90734 124326 92867 124328
rect 90734 124152 90794 124326
rect 92801 124323 92867 124326
rect 142481 124386 142547 124389
rect 142481 124384 145074 124386
rect 142481 124328 142486 124384
rect 142542 124328 145074 124384
rect 142481 124326 145074 124328
rect 142481 124323 142547 124326
rect 134109 124250 134175 124253
rect 131796 124248 134175 124250
rect 131796 124192 134114 124248
rect 134170 124192 134175 124248
rect 131796 124190 134175 124192
rect 134109 124187 134175 124190
rect 145014 124152 145074 124326
rect 177165 124250 177231 124253
rect 174822 124248 177231 124250
rect 174822 124192 177170 124248
rect 177226 124192 177231 124248
rect 174822 124190 177231 124192
rect 50205 124114 50271 124117
rect 47862 124112 50271 124114
rect 47862 124056 50210 124112
rect 50266 124056 50271 124112
rect 47862 124054 50271 124056
rect 50205 124051 50271 124054
rect 58485 124114 58551 124117
rect 58485 124112 60956 124114
rect 58485 124056 58490 124112
rect 58546 124056 60956 124112
rect 58485 124054 60956 124056
rect 58485 124051 58551 124054
rect 92893 123978 92959 123981
rect 90734 123976 92959 123978
rect 47862 123842 47922 123948
rect 90734 123920 92898 123976
rect 92954 123920 92959 123976
rect 90734 123918 92959 123920
rect 51217 123842 51283 123845
rect 47862 123840 51283 123842
rect 47862 123784 51222 123840
rect 51278 123784 51283 123840
rect 47862 123782 51283 123784
rect 51217 123779 51283 123782
rect 51217 123570 51283 123573
rect 47678 123568 51283 123570
rect 47678 123512 51222 123568
rect 51278 123512 51283 123568
rect 47678 123510 51283 123512
rect 47678 123404 47738 123510
rect 51217 123507 51283 123510
rect 90734 123472 90794 123918
rect 92893 123915 92959 123918
rect 101173 123842 101239 123845
rect 103982 123842 104042 124152
rect 174822 124084 174882 124190
rect 177165 124187 177231 124190
rect 142757 123978 142823 123981
rect 177625 123978 177691 123981
rect 142757 123976 145074 123978
rect 142757 123920 142762 123976
rect 142818 123920 145074 123976
rect 142757 123918 145074 123920
rect 142757 123915 142823 123918
rect 101173 123840 104042 123842
rect 101173 123784 101178 123840
rect 101234 123784 104042 123840
rect 101173 123782 104042 123784
rect 101173 123779 101239 123782
rect 135029 123706 135095 123709
rect 131796 123704 135095 123706
rect 131796 123648 135034 123704
rect 135090 123648 135095 123704
rect 131796 123646 135095 123648
rect 135029 123643 135095 123646
rect 58209 123434 58275 123437
rect 100989 123434 101055 123437
rect 103982 123434 104042 123608
rect 145014 123472 145074 123918
rect 174822 123976 177691 123978
rect 174822 123920 177630 123976
rect 177686 123920 177691 123976
rect 174822 123918 177691 123920
rect 58209 123432 60956 123434
rect 58209 123376 58214 123432
rect 58270 123376 60956 123432
rect 58209 123374 60956 123376
rect 100989 123432 104042 123434
rect 100989 123376 100994 123432
rect 101050 123376 104042 123432
rect 174822 123404 174882 123918
rect 177625 123915 177691 123918
rect 185813 123842 185879 123845
rect 187886 123842 187946 124220
rect 185813 123840 187946 123842
rect 185813 123784 185818 123840
rect 185874 123784 187946 123840
rect 185813 123782 187946 123784
rect 185813 123779 185879 123782
rect 185261 123434 185327 123437
rect 187886 123434 187946 123676
rect 185261 123432 187946 123434
rect 100989 123374 104042 123376
rect 185261 123376 185266 123432
rect 185322 123376 187946 123432
rect 185261 123374 187946 123376
rect 58209 123371 58275 123374
rect 100989 123371 101055 123374
rect 185261 123371 185327 123374
rect 143585 123298 143651 123301
rect 143585 123296 145074 123298
rect 143585 123240 143590 123296
rect 143646 123240 145074 123296
rect 143585 123238 145074 123240
rect 143585 123235 143651 123238
rect 92709 123026 92775 123029
rect 135213 123026 135279 123029
rect 90734 123024 92775 123026
rect 90734 122968 92714 123024
rect 92770 122968 92775 123024
rect 90734 122966 92775 122968
rect 131796 123024 135279 123026
rect 131796 122968 135218 123024
rect 135274 122968 135279 123024
rect 131796 122966 135279 122968
rect 90734 122928 90794 122966
rect 92709 122963 92775 122966
rect 135213 122963 135279 122966
rect 145014 122928 145074 123238
rect 177717 123026 177783 123029
rect 174822 123024 177783 123026
rect 174822 122968 177722 123024
rect 177778 122968 177783 123024
rect 174822 122966 177783 122968
rect 58393 122890 58459 122893
rect 58393 122888 60956 122890
rect 47862 122482 47922 122860
rect 58393 122832 58398 122888
rect 58454 122832 60956 122888
rect 58393 122830 60956 122832
rect 58393 122827 58459 122830
rect 92801 122754 92867 122757
rect 90734 122752 92867 122754
rect 90734 122696 92806 122752
rect 92862 122696 92867 122752
rect 90734 122694 92867 122696
rect 51125 122482 51191 122485
rect 47862 122480 51191 122482
rect 47862 122424 51130 122480
rect 51186 122424 51191 122480
rect 47862 122422 51191 122424
rect 51125 122419 51191 122422
rect 47862 122210 47922 122316
rect 90734 122248 90794 122694
rect 92801 122691 92867 122694
rect 101265 122618 101331 122621
rect 103982 122618 104042 122928
rect 174822 122860 174882 122966
rect 177717 122963 177783 122966
rect 177625 122754 177691 122757
rect 101265 122616 104042 122618
rect 101265 122560 101270 122616
rect 101326 122560 104042 122616
rect 101265 122558 104042 122560
rect 174822 122752 177691 122754
rect 174822 122696 177630 122752
rect 177686 122696 177691 122752
rect 174822 122694 177691 122696
rect 101265 122555 101331 122558
rect 135213 122482 135279 122485
rect 131796 122480 135279 122482
rect 131796 122424 135218 122480
rect 135274 122424 135279 122480
rect 131796 122422 135279 122424
rect 135213 122419 135279 122422
rect 143585 122482 143651 122485
rect 143585 122480 145074 122482
rect 143585 122424 143590 122480
rect 143646 122424 145074 122480
rect 143585 122422 145074 122424
rect 143585 122419 143651 122422
rect 51217 122210 51283 122213
rect 47862 122208 51283 122210
rect 47862 122152 51222 122208
rect 51278 122152 51283 122208
rect 47862 122150 51283 122152
rect 51217 122147 51283 122150
rect 58209 122210 58275 122213
rect 58209 122208 60956 122210
rect 58209 122152 58214 122208
rect 58270 122152 60956 122208
rect 58209 122150 60956 122152
rect 58209 122147 58275 122150
rect 101081 122074 101147 122077
rect 103982 122074 104042 122384
rect 145014 122248 145074 122422
rect 174822 122180 174882 122694
rect 177625 122691 177691 122694
rect 185629 122618 185695 122621
rect 187886 122618 187946 122996
rect 185629 122616 187946 122618
rect 185629 122560 185634 122616
rect 185690 122560 187946 122616
rect 185629 122558 187946 122560
rect 185629 122555 185695 122558
rect 185905 122210 185971 122213
rect 187886 122210 187946 122452
rect 185905 122208 187946 122210
rect 185905 122152 185910 122208
rect 185966 122152 187946 122208
rect 185905 122150 187946 122152
rect 185905 122147 185971 122150
rect 101081 122072 104042 122074
rect 101081 122016 101086 122072
rect 101142 122016 104042 122072
rect 101081 122014 104042 122016
rect 101081 122011 101147 122014
rect 134845 121938 134911 121941
rect 131796 121936 134911 121938
rect 131796 121880 134850 121936
rect 134906 121880 134911 121936
rect 131796 121878 134911 121880
rect 134845 121875 134911 121878
rect 92709 121802 92775 121805
rect 90734 121800 92775 121802
rect 47862 121258 47922 121772
rect 90734 121744 92714 121800
rect 92770 121744 92775 121800
rect 90734 121742 92775 121744
rect 90734 121704 90794 121742
rect 92709 121739 92775 121742
rect 58209 121666 58275 121669
rect 58209 121664 60956 121666
rect 58209 121608 58214 121664
rect 58270 121608 60956 121664
rect 58209 121606 60956 121608
rect 58209 121603 58275 121606
rect 92801 121530 92867 121533
rect 90734 121528 92867 121530
rect 90734 121472 92806 121528
rect 92862 121472 92867 121528
rect 90734 121470 92867 121472
rect 51125 121258 51191 121261
rect 47862 121256 51191 121258
rect 47862 121200 51130 121256
rect 51186 121200 51191 121256
rect 47862 121198 51191 121200
rect 51125 121195 51191 121198
rect 90734 121160 90794 121470
rect 92801 121467 92867 121470
rect 100989 121530 101055 121533
rect 103982 121530 104042 121840
rect 143033 121802 143099 121805
rect 177717 121802 177783 121805
rect 143033 121800 145074 121802
rect 143033 121744 143038 121800
rect 143094 121744 145074 121800
rect 143033 121742 145074 121744
rect 143033 121739 143099 121742
rect 145014 121704 145074 121742
rect 174822 121800 177783 121802
rect 174822 121744 177722 121800
rect 177778 121744 177783 121800
rect 174822 121742 177783 121744
rect 174822 121636 174882 121742
rect 177717 121739 177783 121742
rect 100989 121528 104042 121530
rect 100989 121472 100994 121528
rect 101050 121472 104042 121528
rect 100989 121470 104042 121472
rect 142757 121530 142823 121533
rect 177349 121530 177415 121533
rect 142757 121528 145074 121530
rect 142757 121472 142762 121528
rect 142818 121472 145074 121528
rect 142757 121470 145074 121472
rect 100989 121467 101055 121470
rect 142757 121467 142823 121470
rect 134661 121394 134727 121397
rect 131796 121392 134727 121394
rect 131796 121336 134666 121392
rect 134722 121336 134727 121392
rect 131796 121334 134727 121336
rect 134661 121331 134727 121334
rect 58209 121122 58275 121125
rect 58209 121120 60956 121122
rect 47862 120986 47922 121092
rect 58209 121064 58214 121120
rect 58270 121064 60956 121120
rect 58209 121062 60956 121064
rect 58209 121059 58275 121062
rect 51217 120986 51283 120989
rect 47862 120984 51283 120986
rect 47862 120928 51222 120984
rect 51278 120928 51283 120984
rect 47862 120926 51283 120928
rect 51217 120923 51283 120926
rect 101173 120850 101239 120853
rect 103982 120850 104042 121296
rect 145014 121160 145074 121470
rect 174822 121528 177415 121530
rect 174822 121472 177354 121528
rect 177410 121472 177415 121528
rect 174822 121470 177415 121472
rect 174822 121092 174882 121470
rect 177349 121467 177415 121470
rect 185353 121530 185419 121533
rect 187886 121530 187946 121908
rect 185353 121528 187946 121530
rect 185353 121472 185358 121528
rect 185414 121472 187946 121528
rect 185353 121470 187946 121472
rect 185353 121467 185419 121470
rect 101173 120848 104042 120850
rect 101173 120792 101178 120848
rect 101234 120792 104042 120848
rect 101173 120790 104042 120792
rect 185169 120850 185235 120853
rect 187886 120850 187946 121364
rect 185169 120848 187946 120850
rect 185169 120792 185174 120848
rect 185230 120792 187946 120848
rect 185169 120790 187946 120792
rect 101173 120787 101239 120790
rect 185169 120787 185235 120790
rect 100989 120714 101055 120717
rect 135397 120714 135463 120717
rect 100989 120712 104012 120714
rect 100989 120656 100994 120712
rect 101050 120656 104012 120712
rect 100989 120654 104012 120656
rect 131796 120712 135463 120714
rect 131796 120656 135402 120712
rect 135458 120656 135463 120712
rect 131796 120654 135463 120656
rect 100989 120651 101055 120654
rect 135397 120651 135463 120654
rect 185261 120714 185327 120717
rect 185261 120712 187762 120714
rect 185261 120656 185266 120712
rect 185322 120656 187762 120712
rect 185261 120654 187762 120656
rect 185261 120651 185327 120654
rect 142941 120578 143007 120581
rect 177717 120578 177783 120581
rect 142941 120576 145074 120578
rect 47862 120170 47922 120548
rect 142941 120520 142946 120576
rect 143002 120520 145074 120576
rect 142941 120518 145074 120520
rect 142941 120515 143007 120518
rect 145014 120480 145074 120518
rect 174822 120576 177783 120578
rect 174822 120520 177722 120576
rect 177778 120520 177783 120576
rect 174822 120518 177783 120520
rect 187702 120578 187762 120654
rect 187886 120578 187946 120684
rect 187702 120518 187946 120578
rect 58209 120442 58275 120445
rect 92709 120442 92775 120445
rect 58209 120440 60956 120442
rect 58209 120384 58214 120440
rect 58270 120384 60956 120440
rect 58209 120382 60956 120384
rect 90764 120440 92775 120442
rect 90764 120384 92714 120440
rect 92770 120384 92775 120440
rect 174822 120412 174882 120518
rect 177717 120515 177783 120518
rect 90764 120382 92775 120384
rect 58209 120379 58275 120382
rect 92709 120379 92775 120382
rect 143585 120306 143651 120309
rect 177625 120306 177691 120309
rect 143585 120304 145074 120306
rect 143585 120248 143590 120304
rect 143646 120248 145074 120304
rect 143585 120246 145074 120248
rect 143585 120243 143651 120246
rect 50205 120170 50271 120173
rect 134293 120170 134359 120173
rect 47862 120168 50271 120170
rect 47862 120112 50210 120168
rect 50266 120112 50271 120168
rect 47862 120110 50271 120112
rect 131796 120168 134359 120170
rect 131796 120112 134298 120168
rect 134354 120112 134359 120168
rect 131796 120110 134359 120112
rect 50205 120107 50271 120110
rect 134293 120107 134359 120110
rect 92801 120034 92867 120037
rect 90734 120032 92867 120034
rect 18005 119354 18071 119357
rect 19894 119354 19954 119868
rect 47862 119762 47922 120004
rect 90734 119976 92806 120032
rect 92862 119976 92867 120032
rect 90734 119974 92867 119976
rect 90734 119936 90794 119974
rect 92801 119971 92867 119974
rect 58393 119898 58459 119901
rect 58393 119896 60956 119898
rect 58393 119840 58398 119896
rect 58454 119840 60956 119896
rect 58393 119838 60956 119840
rect 58393 119835 58459 119838
rect 51217 119762 51283 119765
rect 47862 119760 51283 119762
rect 47862 119704 51222 119760
rect 51278 119704 51283 119760
rect 47862 119702 51283 119704
rect 51217 119699 51283 119702
rect 101081 119762 101147 119765
rect 103982 119762 104042 120072
rect 145014 119936 145074 120246
rect 174822 120304 177691 120306
rect 174822 120248 177630 120304
rect 177686 120248 177691 120304
rect 174822 120246 177691 120248
rect 174822 119868 174882 120246
rect 177625 120243 177691 120246
rect 101081 119760 104042 119762
rect 101081 119704 101086 119760
rect 101142 119704 104042 119760
rect 101081 119702 104042 119704
rect 185261 119762 185327 119765
rect 187886 119762 187946 120140
rect 185261 119760 187946 119762
rect 185261 119704 185266 119760
rect 185322 119704 187946 119760
rect 185261 119702 187946 119704
rect 101081 119699 101147 119702
rect 185261 119699 185327 119702
rect 135397 119626 135463 119629
rect 131796 119624 135463 119626
rect 131796 119568 135402 119624
rect 135458 119568 135463 119624
rect 131796 119566 135463 119568
rect 135397 119563 135463 119566
rect 18005 119352 19954 119354
rect 18005 119296 18010 119352
rect 18066 119296 19954 119352
rect 18005 119294 19954 119296
rect 47862 119354 47922 119460
rect 51217 119354 51283 119357
rect 47862 119352 51283 119354
rect 47862 119296 51222 119352
rect 51278 119296 51283 119352
rect 47862 119294 51283 119296
rect 18005 119291 18071 119294
rect 51217 119291 51283 119294
rect 100989 119354 101055 119357
rect 103982 119354 104042 119528
rect 100989 119352 104042 119354
rect 100989 119296 100994 119352
rect 101050 119296 104042 119352
rect 100989 119294 104042 119296
rect 185169 119354 185235 119357
rect 187886 119354 187946 119596
rect 185169 119352 187946 119354
rect 185169 119296 185174 119352
rect 185230 119296 187946 119352
rect 185169 119294 187946 119296
rect 100989 119291 101055 119294
rect 185169 119291 185235 119294
rect 58301 119218 58367 119221
rect 92709 119218 92775 119221
rect 58301 119216 60956 119218
rect 58301 119160 58306 119216
rect 58362 119160 60956 119216
rect 58301 119158 60956 119160
rect 90764 119216 92775 119218
rect 90764 119160 92714 119216
rect 92770 119160 92775 119216
rect 90764 119158 92775 119160
rect 58301 119155 58367 119158
rect 92709 119155 92775 119158
rect 143585 119218 143651 119221
rect 143585 119216 145044 119218
rect 143585 119160 143590 119216
rect 143646 119160 145044 119216
rect 143585 119158 145044 119160
rect 143585 119155 143651 119158
rect 174822 119082 174882 119188
rect 177717 119082 177783 119085
rect 174822 119080 177783 119082
rect 174822 119024 177722 119080
rect 177778 119024 177783 119080
rect 174822 119022 177783 119024
rect 177717 119019 177783 119022
rect 92801 118946 92867 118949
rect 134845 118946 134911 118949
rect 90734 118944 92867 118946
rect 47862 118402 47922 118916
rect 90734 118888 92806 118944
rect 92862 118888 92867 118944
rect 90734 118886 92867 118888
rect 131796 118944 134911 118946
rect 131796 118888 134850 118944
rect 134906 118888 134911 118944
rect 131796 118886 134911 118888
rect 90734 118712 90794 118886
rect 92801 118883 92867 118886
rect 134845 118883 134911 118886
rect 143033 118946 143099 118949
rect 143033 118944 145074 118946
rect 143033 118888 143038 118944
rect 143094 118888 145074 118944
rect 143033 118886 145074 118888
rect 143033 118883 143099 118886
rect 58485 118674 58551 118677
rect 58485 118672 60956 118674
rect 58485 118616 58490 118672
rect 58546 118616 60956 118672
rect 58485 118614 60956 118616
rect 58485 118611 58551 118614
rect 92893 118538 92959 118541
rect 90734 118536 92959 118538
rect 90734 118480 92898 118536
rect 92954 118480 92959 118536
rect 90734 118478 92959 118480
rect 50573 118402 50639 118405
rect 47862 118400 50639 118402
rect 47862 118344 50578 118400
rect 50634 118344 50639 118400
rect 47862 118342 50639 118344
rect 50573 118339 50639 118342
rect 47862 118130 47922 118236
rect 90734 118168 90794 118478
rect 92893 118475 92959 118478
rect 101081 118538 101147 118541
rect 103982 118538 104042 118848
rect 145014 118712 145074 118886
rect 177717 118810 177783 118813
rect 174822 118808 177783 118810
rect 174822 118752 177722 118808
rect 177778 118752 177783 118808
rect 174822 118750 177783 118752
rect 174822 118644 174882 118750
rect 177717 118747 177783 118750
rect 101081 118536 104042 118538
rect 101081 118480 101086 118536
rect 101142 118480 104042 118536
rect 101081 118478 104042 118480
rect 143309 118538 143375 118541
rect 177625 118538 177691 118541
rect 143309 118536 145074 118538
rect 143309 118480 143314 118536
rect 143370 118480 145074 118536
rect 143309 118478 145074 118480
rect 101081 118475 101147 118478
rect 143309 118475 143375 118478
rect 134477 118402 134543 118405
rect 131796 118400 134543 118402
rect 131796 118344 134482 118400
rect 134538 118344 134543 118400
rect 131796 118342 134543 118344
rect 134477 118339 134543 118342
rect 51217 118130 51283 118133
rect 47862 118128 51283 118130
rect 47862 118072 51222 118128
rect 51278 118072 51283 118128
rect 47862 118070 51283 118072
rect 51217 118067 51283 118070
rect 58209 118130 58275 118133
rect 58209 118128 60956 118130
rect 58209 118072 58214 118128
rect 58270 118072 60956 118128
rect 58209 118070 60956 118072
rect 58209 118067 58275 118070
rect 100989 117994 101055 117997
rect 103982 117994 104042 118304
rect 145014 118168 145074 118478
rect 174822 118536 177691 118538
rect 174822 118480 177630 118536
rect 177686 118480 177691 118536
rect 174822 118478 177691 118480
rect 174822 118100 174882 118478
rect 177625 118475 177691 118478
rect 185261 118538 185327 118541
rect 187886 118538 187946 118916
rect 185261 118536 187946 118538
rect 185261 118480 185266 118536
rect 185322 118480 187946 118536
rect 185261 118478 187946 118480
rect 185261 118475 185327 118478
rect 100989 117992 104042 117994
rect 100989 117936 100994 117992
rect 101050 117936 104042 117992
rect 100989 117934 104042 117936
rect 185169 117994 185235 117997
rect 187886 117994 187946 118372
rect 185169 117992 187946 117994
rect 185169 117936 185174 117992
rect 185230 117936 187946 117992
rect 185169 117934 187946 117936
rect 100989 117931 101055 117934
rect 185169 117931 185235 117934
rect 134845 117858 134911 117861
rect 218289 117858 218355 117861
rect 131796 117856 134911 117858
rect 131796 117800 134850 117856
rect 134906 117800 134911 117856
rect 215670 117856 218355 117858
rect 131796 117798 134911 117800
rect 134845 117795 134911 117798
rect 47862 117314 47922 117692
rect 92709 117586 92775 117589
rect 90734 117584 92775 117586
rect 90734 117528 92714 117584
rect 92770 117528 92775 117584
rect 90734 117526 92775 117528
rect 90734 117488 90794 117526
rect 92709 117523 92775 117526
rect 58209 117450 58275 117453
rect 101173 117450 101239 117453
rect 103982 117450 104042 117760
rect 142573 117722 142639 117725
rect 142573 117720 145074 117722
rect 142573 117664 142578 117720
rect 142634 117664 145074 117720
rect 142573 117662 145074 117664
rect 142573 117659 142639 117662
rect 145014 117488 145074 117662
rect 177717 117586 177783 117589
rect 174822 117584 177783 117586
rect 174822 117528 177722 117584
rect 177778 117528 177783 117584
rect 174822 117526 177783 117528
rect 58209 117448 60956 117450
rect 58209 117392 58214 117448
rect 58270 117392 60956 117448
rect 58209 117390 60956 117392
rect 101173 117448 104042 117450
rect 101173 117392 101178 117448
rect 101234 117392 104042 117448
rect 174822 117420 174882 117526
rect 177717 117523 177783 117526
rect 185353 117450 185419 117453
rect 187886 117450 187946 117828
rect 215670 117800 218294 117856
rect 218350 117800 218355 117856
rect 215670 117798 218355 117800
rect 215670 117556 215730 117798
rect 218289 117795 218355 117798
rect 185353 117448 187946 117450
rect 101173 117390 104042 117392
rect 185353 117392 185358 117448
rect 185414 117392 187946 117448
rect 185353 117390 187946 117392
rect 58209 117387 58275 117390
rect 101173 117387 101239 117390
rect 185353 117387 185419 117390
rect 50021 117314 50087 117317
rect 134937 117314 135003 117317
rect 47862 117312 50087 117314
rect 47862 117256 50026 117312
rect 50082 117256 50087 117312
rect 47862 117254 50087 117256
rect 131796 117312 135003 117314
rect 131796 117256 134942 117312
rect 134998 117256 135003 117312
rect 131796 117254 135003 117256
rect 50021 117251 50087 117254
rect 134937 117251 135003 117254
rect 143217 117314 143283 117317
rect 143217 117312 145074 117314
rect 143217 117256 143222 117312
rect 143278 117256 145074 117312
rect 143217 117254 145074 117256
rect 143217 117251 143283 117254
rect 92801 117178 92867 117181
rect 90734 117176 92867 117178
rect 47862 116770 47922 117148
rect 90734 117120 92806 117176
rect 92862 117120 92867 117176
rect 90734 117118 92867 117120
rect 90734 116944 90794 117118
rect 92801 117115 92867 117118
rect 58301 116906 58367 116909
rect 58301 116904 60956 116906
rect 58301 116848 58306 116904
rect 58362 116848 60956 116904
rect 58301 116846 60956 116848
rect 58301 116843 58367 116846
rect 50573 116770 50639 116773
rect 47862 116768 50639 116770
rect 47862 116712 50578 116768
rect 50634 116712 50639 116768
rect 47862 116710 50639 116712
rect 50573 116707 50639 116710
rect 101081 116770 101147 116773
rect 103982 116770 104042 117216
rect 145014 116944 145074 117254
rect 177165 117178 177231 117181
rect 174822 117176 177231 117178
rect 174822 117120 177170 117176
rect 177226 117120 177231 117176
rect 174822 117118 177231 117120
rect 174822 116876 174882 117118
rect 177165 117115 177231 117118
rect 101081 116768 104042 116770
rect 101081 116712 101086 116768
rect 101142 116712 104042 116768
rect 101081 116710 104042 116712
rect 185261 116770 185327 116773
rect 187886 116770 187946 117284
rect 185261 116768 187946 116770
rect 185261 116712 185266 116768
rect 185322 116712 187946 116768
rect 185261 116710 187946 116712
rect 101081 116707 101147 116710
rect 185261 116707 185327 116710
rect 100989 116634 101055 116637
rect 134753 116634 134819 116637
rect 100989 116632 104012 116634
rect 47862 116498 47922 116604
rect 100989 116576 100994 116632
rect 101050 116576 104012 116632
rect 100989 116574 104012 116576
rect 131796 116632 134819 116634
rect 131796 116576 134758 116632
rect 134814 116576 134819 116632
rect 131796 116574 134819 116576
rect 100989 116571 101055 116574
rect 134753 116571 134819 116574
rect 50757 116498 50823 116501
rect 47862 116496 50823 116498
rect 47862 116440 50762 116496
rect 50818 116440 50823 116496
rect 47862 116438 50823 116440
rect 50757 116435 50823 116438
rect 185169 116498 185235 116501
rect 187886 116498 187946 116604
rect 185169 116496 187946 116498
rect 185169 116440 185174 116496
rect 185230 116440 187946 116496
rect 185169 116438 187946 116440
rect 185169 116435 185235 116438
rect 142941 116362 143007 116365
rect 177717 116362 177783 116365
rect 142941 116360 145074 116362
rect 142941 116304 142946 116360
rect 143002 116304 145074 116360
rect 142941 116302 145074 116304
rect 142941 116299 143007 116302
rect 145014 116264 145074 116302
rect 174822 116360 177783 116362
rect 174822 116304 177722 116360
rect 177778 116304 177783 116360
rect 174822 116302 177783 116304
rect 58301 116226 58367 116229
rect 92709 116226 92775 116229
rect 58301 116224 60956 116226
rect 58301 116168 58306 116224
rect 58362 116168 60956 116224
rect 58301 116166 60956 116168
rect 90764 116224 92775 116226
rect 90764 116168 92714 116224
rect 92770 116168 92775 116224
rect 174822 116196 174882 116302
rect 177717 116299 177783 116302
rect 90764 116166 92775 116168
rect 58301 116163 58367 116166
rect 92709 116163 92775 116166
rect 134845 116090 134911 116093
rect 131796 116088 134911 116090
rect 47862 115546 47922 116060
rect 131796 116032 134850 116088
rect 134906 116032 134911 116088
rect 131796 116030 134911 116032
rect 134845 116027 134911 116030
rect 143585 116090 143651 116093
rect 143585 116088 145074 116090
rect 143585 116032 143590 116088
rect 143646 116032 145074 116088
rect 143585 116030 145074 116032
rect 143585 116027 143651 116030
rect 92801 115818 92867 115821
rect 90734 115816 92867 115818
rect 90734 115760 92806 115816
rect 92862 115760 92867 115816
rect 90734 115758 92867 115760
rect 90734 115720 90794 115758
rect 92801 115755 92867 115758
rect 58393 115682 58459 115685
rect 101081 115682 101147 115685
rect 103982 115682 104042 115992
rect 145014 115720 145074 116030
rect 177717 115954 177783 115957
rect 174822 115952 177783 115954
rect 174822 115896 177722 115952
rect 177778 115896 177783 115952
rect 174822 115894 177783 115896
rect 58393 115680 60956 115682
rect 58393 115624 58398 115680
rect 58454 115624 60956 115680
rect 58393 115622 60956 115624
rect 101081 115680 104042 115682
rect 101081 115624 101086 115680
rect 101142 115624 104042 115680
rect 174822 115652 174882 115894
rect 177717 115891 177783 115894
rect 185261 115682 185327 115685
rect 187886 115682 187946 116060
rect 185261 115680 187946 115682
rect 101081 115622 104042 115624
rect 185261 115624 185266 115680
rect 185322 115624 187946 115680
rect 185261 115622 187946 115624
rect 58393 115619 58459 115622
rect 101081 115619 101147 115622
rect 185261 115619 185327 115622
rect 50665 115546 50731 115549
rect 92893 115546 92959 115549
rect 135029 115546 135095 115549
rect 47862 115544 50731 115546
rect 47862 115488 50670 115544
rect 50726 115488 50731 115544
rect 47862 115486 50731 115488
rect 50665 115483 50731 115486
rect 90734 115544 92959 115546
rect 90734 115488 92898 115544
rect 92954 115488 92959 115544
rect 90734 115486 92959 115488
rect 131796 115544 135095 115546
rect 131796 115488 135034 115544
rect 135090 115488 135095 115544
rect 131796 115486 135095 115488
rect 47862 115138 47922 115380
rect 90734 115176 90794 115486
rect 92893 115483 92959 115486
rect 135029 115483 135095 115486
rect 142757 115546 142823 115549
rect 177073 115546 177139 115549
rect 142757 115544 145074 115546
rect 142757 115488 142762 115544
rect 142818 115488 145074 115544
rect 142757 115486 145074 115488
rect 142757 115483 142823 115486
rect 100989 115274 101055 115277
rect 103982 115274 104042 115448
rect 100989 115272 104042 115274
rect 100989 115216 100994 115272
rect 101050 115216 104042 115272
rect 100989 115214 104042 115216
rect 100989 115211 101055 115214
rect 145014 115176 145074 115486
rect 174822 115544 177139 115546
rect 174822 115488 177078 115544
rect 177134 115488 177139 115544
rect 174822 115486 177139 115488
rect 50849 115138 50915 115141
rect 47862 115136 50915 115138
rect 47862 115080 50854 115136
rect 50910 115080 50915 115136
rect 47862 115078 50915 115080
rect 50849 115075 50915 115078
rect 58209 115138 58275 115141
rect 58209 115136 60956 115138
rect 58209 115080 58214 115136
rect 58270 115080 60956 115136
rect 174822 115108 174882 115486
rect 177073 115483 177139 115486
rect 185169 115274 185235 115277
rect 187886 115274 187946 115516
rect 185169 115272 187946 115274
rect 185169 115216 185174 115272
rect 185230 115216 187946 115272
rect 185169 115214 187946 115216
rect 185169 115211 185235 115214
rect 58209 115078 60956 115080
rect 58209 115075 58275 115078
rect 9896 115002 10376 115032
rect 13405 115002 13471 115005
rect 9896 115000 13471 115002
rect 9896 114944 13410 115000
rect 13466 114944 13471 115000
rect 9896 114942 13471 114944
rect 9896 114912 10376 114942
rect 13405 114939 13471 114942
rect 135121 114866 135187 114869
rect 131796 114864 135187 114866
rect 47862 114458 47922 114836
rect 131796 114808 135126 114864
rect 135182 114808 135187 114864
rect 131796 114806 135187 114808
rect 135121 114803 135187 114806
rect 51125 114458 51191 114461
rect 47862 114456 51191 114458
rect 47862 114400 51130 114456
rect 51186 114400 51191 114456
rect 47862 114398 51191 114400
rect 51125 114395 51191 114398
rect 102001 114458 102067 114461
rect 103982 114458 104042 114768
rect 102001 114456 104042 114458
rect 102001 114400 102006 114456
rect 102062 114400 104042 114456
rect 102001 114398 104042 114400
rect 185997 114458 186063 114461
rect 187886 114458 187946 114836
rect 185997 114456 187946 114458
rect 185997 114400 186002 114456
rect 186058 114400 187946 114456
rect 185997 114398 187946 114400
rect 102001 114395 102067 114398
rect 185997 114395 186063 114398
rect 135305 114322 135371 114325
rect 131796 114320 135371 114322
rect 47862 113914 47922 114292
rect 131796 114264 135310 114320
rect 135366 114264 135371 114320
rect 131796 114262 135371 114264
rect 135305 114259 135371 114262
rect 50481 113914 50547 113917
rect 47862 113912 50547 113914
rect 47862 113856 50486 113912
rect 50542 113856 50547 113912
rect 47862 113854 50547 113856
rect 50481 113851 50547 113854
rect 101633 113914 101699 113917
rect 103982 113914 104042 114224
rect 101633 113912 104042 113914
rect 101633 113856 101638 113912
rect 101694 113856 104042 113912
rect 101633 113854 104042 113856
rect 185813 113914 185879 113917
rect 187886 113914 187946 114292
rect 185813 113912 187946 113914
rect 185813 113856 185818 113912
rect 185874 113856 187946 113912
rect 185813 113854 187946 113856
rect 101633 113851 101699 113854
rect 185813 113851 185879 113854
rect 50941 113778 51007 113781
rect 48046 113776 51007 113778
rect 47862 113642 47922 113748
rect 48046 113720 50946 113776
rect 51002 113720 51007 113776
rect 48046 113718 51007 113720
rect 48046 113642 48106 113718
rect 50941 113715 51007 113718
rect 101817 113778 101883 113781
rect 135397 113778 135463 113781
rect 101817 113776 104012 113778
rect 101817 113720 101822 113776
rect 101878 113720 104012 113776
rect 101817 113718 104012 113720
rect 131796 113776 135463 113778
rect 131796 113720 135402 113776
rect 135458 113720 135463 113776
rect 131796 113718 135463 113720
rect 101817 113715 101883 113718
rect 135397 113715 135463 113718
rect 186181 113778 186247 113781
rect 186181 113776 187762 113778
rect 186181 113720 186186 113776
rect 186242 113720 187762 113776
rect 186181 113718 187762 113720
rect 186181 113715 186247 113718
rect 47862 113582 48106 113642
rect 187702 113642 187762 113718
rect 187886 113642 187946 113748
rect 187702 113582 187946 113642
rect 135213 113234 135279 113237
rect 131796 113232 135279 113234
rect 47862 112826 47922 113204
rect 131796 113176 135218 113232
rect 135274 113176 135279 113232
rect 131796 113174 135279 113176
rect 135213 113171 135279 113174
rect 51217 112826 51283 112829
rect 47862 112824 51283 112826
rect 47862 112768 51222 112824
rect 51278 112768 51283 112824
rect 47862 112766 51283 112768
rect 51217 112763 51283 112766
rect 100989 112554 101055 112557
rect 103982 112554 104042 113136
rect 185169 112690 185235 112693
rect 187886 112690 187946 113204
rect 185169 112688 187946 112690
rect 185169 112632 185174 112688
rect 185230 112632 187946 112688
rect 185169 112630 187946 112632
rect 185169 112627 185235 112630
rect 100989 112552 104042 112554
rect 100989 112496 100994 112552
rect 101050 112496 104042 112552
rect 100989 112494 104042 112496
rect 100989 112491 101055 112494
rect 220957 100586 221023 100589
rect 225416 100586 225896 100616
rect 220957 100584 225896 100586
rect 220957 100528 220962 100584
rect 221018 100528 225896 100584
rect 220957 100526 225896 100528
rect 220957 100523 221023 100526
rect 225416 100496 225896 100526
rect 98781 99770 98847 99773
rect 95702 99768 98847 99770
rect 95702 99712 98786 99768
rect 98842 99712 98847 99768
rect 95702 99710 98847 99712
rect 95702 99224 95762 99710
rect 98781 99707 98847 99710
rect 183697 99226 183763 99229
rect 179820 99224 183763 99226
rect 179820 99168 183702 99224
rect 183758 99168 183763 99224
rect 179820 99166 183763 99168
rect 183697 99163 183763 99166
rect 191977 98818 192043 98821
rect 191977 98816 193988 98818
rect 191977 98760 191982 98816
rect 192038 98760 193988 98816
rect 191977 98758 193988 98760
rect 191977 98755 192043 98758
rect 99517 98546 99583 98549
rect 95702 98544 99583 98546
rect 95702 98488 99522 98544
rect 99578 98488 99583 98544
rect 95702 98486 99583 98488
rect 95702 98000 95762 98486
rect 99517 98483 99583 98486
rect 106785 98546 106851 98549
rect 106785 98544 109900 98546
rect 106785 98488 106790 98544
rect 106846 98488 109900 98544
rect 106785 98486 109900 98488
rect 106785 98483 106851 98486
rect 183605 98002 183671 98005
rect 179820 98000 183671 98002
rect 179820 97944 183610 98000
rect 183666 97944 183671 98000
rect 179820 97942 183671 97944
rect 183605 97939 183671 97942
rect 99425 97050 99491 97053
rect 95702 97048 99491 97050
rect 95702 96992 99430 97048
rect 99486 96992 99491 97048
rect 95702 96990 99491 96992
rect 95702 96776 95762 96990
rect 99425 96987 99491 96990
rect 193766 96852 193772 96916
rect 193836 96852 193842 96916
rect 209825 96914 209891 96917
rect 209782 96912 209891 96914
rect 209782 96856 209830 96912
rect 209886 96856 209891 96912
rect 183513 96778 183579 96781
rect 179820 96776 183579 96778
rect 179820 96720 183518 96776
rect 183574 96720 183579 96776
rect 179820 96718 183579 96720
rect 193774 96778 193834 96852
rect 209782 96851 209891 96856
rect 209782 96780 209842 96851
rect 193774 96718 193988 96778
rect 183513 96715 183579 96718
rect 209774 96716 209780 96780
rect 209844 96716 209850 96780
rect 22329 96506 22395 96509
rect 212309 96506 212375 96509
rect 22329 96504 25996 96506
rect 22329 96448 22334 96504
rect 22390 96448 25996 96504
rect 22329 96446 25996 96448
rect 209812 96504 212375 96506
rect 209812 96448 212314 96504
rect 212370 96448 212375 96504
rect 209812 96446 212375 96448
rect 22329 96443 22395 96446
rect 212309 96443 212375 96446
rect 106785 96234 106851 96237
rect 106785 96232 109900 96234
rect 106785 96176 106790 96232
rect 106846 96176 109900 96232
rect 106785 96174 109900 96176
rect 106785 96171 106851 96174
rect 99241 95554 99307 95557
rect 183329 95554 183395 95557
rect 95732 95552 99307 95554
rect 95732 95496 99246 95552
rect 99302 95496 99307 95552
rect 95732 95494 99307 95496
rect 179820 95552 183395 95554
rect 179820 95496 183334 95552
rect 183390 95496 183395 95552
rect 179820 95494 183395 95496
rect 99241 95491 99307 95494
rect 183329 95491 183395 95494
rect 41833 95282 41899 95285
rect 41790 95280 41899 95282
rect 41790 95224 41838 95280
rect 41894 95224 41899 95280
rect 41790 95219 41899 95224
rect 41790 94708 41850 95219
rect 191977 94738 192043 94741
rect 191977 94736 193988 94738
rect 191977 94680 191982 94736
rect 192038 94680 193988 94736
rect 191977 94678 193988 94680
rect 191977 94675 192043 94678
rect 99149 94330 99215 94333
rect 183237 94330 183303 94333
rect 95732 94328 99215 94330
rect 95732 94272 99154 94328
rect 99210 94272 99215 94328
rect 95732 94270 99215 94272
rect 179820 94328 183303 94330
rect 179820 94272 183242 94328
rect 183298 94272 183303 94328
rect 179820 94270 183303 94272
rect 99149 94267 99215 94270
rect 183237 94267 183303 94270
rect 106509 93922 106575 93925
rect 106509 93920 109900 93922
rect 106509 93864 106514 93920
rect 106570 93864 109900 93920
rect 106509 93862 109900 93864
rect 106509 93859 106575 93862
rect 99333 93650 99399 93653
rect 95702 93648 99399 93650
rect 95702 93592 99338 93648
rect 99394 93592 99399 93648
rect 95702 93590 99399 93592
rect 95702 93104 95762 93590
rect 99333 93587 99399 93590
rect 183421 93106 183487 93109
rect 179820 93104 183487 93106
rect 179820 93048 183426 93104
rect 183482 93048 183487 93104
rect 179820 93046 183487 93048
rect 183421 93043 183487 93046
rect 191149 92834 191215 92837
rect 191149 92832 193988 92834
rect 191149 92776 191154 92832
rect 191210 92776 193988 92832
rect 191149 92774 193988 92776
rect 191149 92771 191215 92774
rect 99057 92426 99123 92429
rect 95702 92424 99123 92426
rect 95702 92368 99062 92424
rect 99118 92368 99123 92424
rect 95702 92366 99123 92368
rect 95702 91880 95762 92366
rect 99057 92363 99123 92366
rect 183145 91882 183211 91885
rect 179820 91880 183211 91882
rect 179820 91824 183150 91880
rect 183206 91824 183211 91880
rect 179820 91822 183211 91824
rect 183145 91819 183211 91822
rect 106785 91474 106851 91477
rect 106785 91472 109900 91474
rect 106785 91416 106790 91472
rect 106846 91416 109900 91472
rect 106785 91414 109900 91416
rect 106785 91411 106851 91414
rect 9896 91338 10376 91368
rect 13497 91338 13563 91341
rect 9896 91336 13563 91338
rect 9896 91280 13502 91336
rect 13558 91280 13563 91336
rect 9896 91278 13563 91280
rect 9896 91248 10376 91278
rect 13497 91275 13563 91278
rect 98965 91202 99031 91205
rect 95702 91200 99031 91202
rect 95702 91144 98970 91200
rect 99026 91144 99031 91200
rect 95702 91142 99031 91144
rect 95702 90656 95762 91142
rect 98965 91139 99031 91142
rect 190781 90794 190847 90797
rect 190781 90792 193988 90794
rect 190781 90736 190786 90792
rect 190842 90736 193988 90792
rect 190781 90734 193988 90736
rect 190781 90731 190847 90734
rect 183053 90658 183119 90661
rect 179820 90656 183119 90658
rect 179820 90600 183058 90656
rect 183114 90600 183119 90656
rect 179820 90598 183119 90600
rect 183053 90595 183119 90598
rect 98781 89978 98847 89981
rect 95702 89976 98847 89978
rect 95702 89920 98786 89976
rect 98842 89920 98847 89976
rect 95702 89918 98847 89920
rect 22329 89842 22395 89845
rect 22329 89840 25996 89842
rect 22329 89784 22334 89840
rect 22390 89784 25996 89840
rect 22329 89782 25996 89784
rect 22329 89779 22395 89782
rect 95702 89432 95762 89918
rect 98781 89915 98847 89918
rect 128497 89842 128563 89845
rect 212125 89842 212191 89845
rect 125724 89840 128563 89842
rect 125724 89784 128502 89840
rect 128558 89784 128563 89840
rect 125724 89782 128563 89784
rect 209812 89840 212191 89842
rect 209812 89784 212130 89840
rect 212186 89784 212191 89840
rect 209812 89782 212191 89784
rect 128497 89779 128563 89782
rect 212125 89779 212191 89782
rect 182869 89434 182935 89437
rect 179820 89432 182935 89434
rect 179820 89376 182874 89432
rect 182930 89376 182935 89432
rect 179820 89374 182935 89376
rect 182869 89371 182935 89374
rect 106785 89162 106851 89165
rect 106785 89160 109900 89162
rect 106785 89104 106790 89160
rect 106846 89104 109900 89160
rect 106785 89102 109900 89104
rect 106785 89099 106851 89102
rect 99517 88754 99583 88757
rect 95702 88752 99583 88754
rect 95702 88696 99522 88752
rect 99578 88696 99583 88752
rect 95702 88694 99583 88696
rect 95702 88208 95762 88694
rect 99517 88691 99583 88694
rect 191701 88754 191767 88757
rect 191701 88752 193988 88754
rect 191701 88696 191706 88752
rect 191762 88696 193988 88752
rect 191701 88694 193988 88696
rect 191701 88691 191767 88694
rect 183513 88210 183579 88213
rect 179820 88208 183579 88210
rect 179820 88152 183518 88208
rect 183574 88152 183579 88208
rect 179820 88150 183579 88152
rect 183513 88147 183579 88150
rect 98689 87394 98755 87397
rect 95702 87392 98755 87394
rect 95702 87336 98694 87392
rect 98750 87336 98755 87392
rect 95702 87334 98755 87336
rect 95702 87120 95762 87334
rect 98689 87331 98755 87334
rect 183697 87122 183763 87125
rect 179820 87120 183763 87122
rect 179820 87064 183702 87120
rect 183758 87064 183763 87120
rect 179820 87062 183763 87064
rect 183697 87059 183763 87062
rect 106785 86850 106851 86853
rect 191609 86850 191675 86853
rect 106785 86848 109900 86850
rect 106785 86792 106790 86848
rect 106846 86792 109900 86848
rect 106785 86790 109900 86792
rect 191609 86848 193988 86850
rect 191609 86792 191614 86848
rect 191670 86792 193988 86848
rect 191609 86790 193988 86792
rect 106785 86787 106851 86790
rect 191609 86787 191675 86790
rect 183697 85898 183763 85901
rect 179820 85896 183763 85898
rect 179820 85840 183702 85896
rect 183758 85840 183763 85896
rect 95702 85354 95762 85840
rect 179820 85838 183763 85840
rect 183697 85835 183763 85838
rect 99517 85354 99583 85357
rect 95702 85352 99583 85354
rect 95702 85296 99522 85352
rect 99578 85296 99583 85352
rect 95702 85294 99583 85296
rect 99517 85291 99583 85294
rect 44409 84810 44475 84813
rect 41820 84808 44475 84810
rect 41820 84752 44414 84808
rect 44470 84752 44475 84808
rect 41820 84750 44475 84752
rect 44409 84747 44475 84750
rect 191977 84810 192043 84813
rect 191977 84808 193988 84810
rect 191977 84752 191982 84808
rect 192038 84752 193988 84808
rect 191977 84750 193988 84752
rect 191977 84747 192043 84750
rect 99517 84674 99583 84677
rect 183697 84674 183763 84677
rect 95732 84672 99583 84674
rect 95732 84616 99522 84672
rect 99578 84616 99583 84672
rect 95732 84614 99583 84616
rect 179820 84672 183763 84674
rect 179820 84616 183702 84672
rect 183758 84616 183763 84672
rect 179820 84614 183763 84616
rect 99517 84611 99583 84614
rect 183697 84611 183763 84614
rect 107797 84402 107863 84405
rect 107797 84400 109900 84402
rect 107797 84344 107802 84400
rect 107858 84344 109900 84400
rect 107797 84342 109900 84344
rect 107797 84339 107863 84342
rect 99425 83994 99491 83997
rect 95702 83992 99491 83994
rect 95702 83936 99430 83992
rect 99486 83936 99491 83992
rect 95702 83934 99491 83936
rect 95702 83448 95762 83934
rect 99425 83931 99491 83934
rect 182501 83450 182567 83453
rect 179820 83448 182567 83450
rect 179820 83392 182506 83448
rect 182562 83392 182567 83448
rect 179820 83390 182567 83392
rect 182501 83387 182567 83390
rect 22329 83178 22395 83181
rect 212033 83178 212099 83181
rect 22329 83176 25996 83178
rect 22329 83120 22334 83176
rect 22390 83120 25996 83176
rect 22329 83118 25996 83120
rect 209812 83176 212099 83178
rect 209812 83120 212038 83176
rect 212094 83120 212099 83176
rect 209812 83118 212099 83120
rect 22329 83115 22395 83118
rect 212033 83115 212099 83118
rect 99517 82770 99583 82773
rect 95702 82768 99583 82770
rect 95702 82712 99522 82768
rect 99578 82712 99583 82768
rect 95702 82710 99583 82712
rect 95702 82224 95762 82710
rect 99517 82707 99583 82710
rect 191977 82770 192043 82773
rect 191977 82768 193988 82770
rect 191977 82712 191982 82768
rect 192038 82712 193988 82768
rect 191977 82710 193988 82712
rect 191977 82707 192043 82710
rect 183697 82226 183763 82229
rect 179820 82224 183763 82226
rect 179820 82168 183702 82224
rect 183758 82168 183763 82224
rect 179820 82166 183763 82168
rect 183697 82163 183763 82166
rect 106785 82090 106851 82093
rect 106785 82088 109900 82090
rect 106785 82032 106790 82088
rect 106846 82032 109900 82088
rect 106785 82030 109900 82032
rect 106785 82027 106851 82030
rect 99517 81546 99583 81549
rect 95702 81544 99583 81546
rect 95702 81488 99522 81544
rect 99578 81488 99583 81544
rect 95702 81486 99583 81488
rect 95702 81000 95762 81486
rect 99517 81483 99583 81486
rect 183237 81002 183303 81005
rect 179820 81000 183303 81002
rect 179820 80944 183242 81000
rect 183298 80944 183303 81000
rect 179820 80942 183303 80944
rect 183237 80939 183303 80942
rect 191885 80866 191951 80869
rect 191885 80864 193988 80866
rect 191885 80808 191890 80864
rect 191946 80808 193988 80864
rect 191885 80806 193988 80808
rect 191885 80803 191951 80806
rect 136869 80458 136935 80461
rect 136869 80456 140106 80458
rect 136869 80400 136874 80456
rect 136930 80400 140106 80456
rect 136869 80398 140106 80400
rect 136869 80395 136935 80398
rect 52689 79914 52755 79917
rect 52689 79912 55988 79914
rect 140046 79912 140106 80398
rect 52689 79856 52694 79912
rect 52750 79856 55988 79912
rect 52689 79854 55988 79856
rect 52689 79851 52755 79854
rect 99517 79778 99583 79781
rect 95732 79776 99583 79778
rect 95732 79720 99522 79776
rect 99578 79720 99583 79776
rect 95732 79718 99583 79720
rect 99517 79715 99583 79718
rect 106785 79778 106851 79781
rect 183697 79778 183763 79781
rect 106785 79776 109900 79778
rect 106785 79720 106790 79776
rect 106846 79720 109900 79776
rect 106785 79718 109900 79720
rect 179820 79776 183763 79778
rect 179820 79720 183702 79776
rect 183758 79720 183763 79776
rect 179820 79718 183763 79720
rect 106785 79715 106851 79718
rect 183697 79715 183763 79718
rect 191977 78826 192043 78829
rect 191977 78824 193988 78826
rect 191977 78768 191982 78824
rect 192038 78768 193988 78824
rect 191977 78766 193988 78768
rect 191977 78763 192043 78766
rect 183513 78554 183579 78557
rect 179820 78552 183579 78554
rect 179820 78496 183518 78552
rect 183574 78496 183579 78552
rect 95702 78010 95762 78496
rect 179820 78494 183579 78496
rect 183513 78491 183579 78494
rect 99517 78010 99583 78013
rect 95702 78008 99583 78010
rect 95702 77952 99522 78008
rect 99578 77952 99583 78008
rect 95702 77950 99583 77952
rect 99517 77947 99583 77950
rect 106509 77466 106575 77469
rect 106509 77464 109900 77466
rect 106509 77408 106514 77464
rect 106570 77408 109900 77464
rect 106509 77406 109900 77408
rect 106509 77403 106575 77406
rect 183053 77330 183119 77333
rect 179820 77328 183119 77330
rect 179820 77272 183058 77328
rect 183114 77272 183119 77328
rect 95702 76786 95762 77272
rect 179820 77270 183119 77272
rect 183053 77267 183119 77270
rect 209825 76922 209891 76925
rect 209782 76920 209891 76922
rect 209782 76864 209830 76920
rect 209886 76864 209891 76920
rect 209782 76859 209891 76864
rect 99517 76786 99583 76789
rect 95702 76784 99583 76786
rect 95702 76728 99522 76784
rect 99578 76728 99583 76784
rect 95702 76726 99583 76728
rect 99517 76723 99583 76726
rect 191977 76786 192043 76789
rect 191977 76784 193988 76786
rect 191977 76728 191982 76784
rect 192038 76728 193988 76784
rect 191977 76726 193988 76728
rect 191977 76723 192043 76726
rect 22329 76514 22395 76517
rect 22329 76512 25996 76514
rect 22329 76456 22334 76512
rect 22390 76456 25996 76512
rect 209782 76484 209842 76859
rect 22329 76454 25996 76456
rect 22329 76451 22395 76454
rect 183237 76106 183303 76109
rect 179820 76104 183303 76106
rect 179820 76048 183242 76104
rect 183298 76048 183303 76104
rect 95702 75562 95762 76048
rect 179820 76046 183303 76048
rect 183237 76043 183303 76046
rect 98229 75562 98295 75565
rect 95702 75560 98295 75562
rect 95702 75504 98234 75560
rect 98290 75504 98295 75560
rect 95702 75502 98295 75504
rect 98229 75499 98295 75502
rect 106785 75018 106851 75021
rect 106785 75016 109900 75018
rect 106785 74960 106790 75016
rect 106846 74960 109900 75016
rect 106785 74958 109900 74960
rect 106785 74955 106851 74958
rect 183697 74882 183763 74885
rect 179820 74880 183763 74882
rect 179820 74824 183702 74880
rect 183758 74824 183763 74880
rect 44409 74746 44475 74749
rect 41820 74744 44475 74746
rect 41820 74688 44414 74744
rect 44470 74688 44475 74744
rect 41820 74686 44475 74688
rect 44409 74683 44475 74686
rect 95702 74338 95762 74824
rect 179820 74822 183763 74824
rect 183697 74819 183763 74822
rect 191517 74746 191583 74749
rect 191517 74744 193988 74746
rect 191517 74688 191522 74744
rect 191578 74688 193988 74744
rect 191517 74686 193988 74688
rect 191517 74683 191583 74686
rect 99425 74338 99491 74341
rect 95702 74336 99491 74338
rect 95702 74280 99430 74336
rect 99486 74280 99491 74336
rect 95702 74278 99491 74280
rect 99425 74275 99491 74278
rect 222337 74338 222403 74341
rect 225416 74338 225896 74368
rect 222337 74336 225896 74338
rect 222337 74280 222342 74336
rect 222398 74280 225896 74336
rect 222337 74278 225896 74280
rect 222337 74275 222403 74278
rect 225416 74248 225896 74278
rect 99517 73794 99583 73797
rect 183697 73794 183763 73797
rect 95732 73792 99583 73794
rect 95732 73736 99522 73792
rect 99578 73736 99583 73792
rect 95732 73734 99583 73736
rect 179820 73792 183763 73794
rect 179820 73736 183702 73792
rect 183758 73736 183763 73792
rect 179820 73734 183763 73736
rect 99517 73731 99583 73734
rect 183697 73731 183763 73734
rect 191977 72842 192043 72845
rect 191977 72840 193988 72842
rect 191977 72784 191982 72840
rect 192038 72784 193988 72840
rect 191977 72782 193988 72784
rect 191977 72779 192043 72782
rect 106785 72706 106851 72709
rect 106785 72704 109900 72706
rect 106785 72648 106790 72704
rect 106846 72648 109900 72704
rect 106785 72646 109900 72648
rect 106785 72643 106851 72646
rect 99517 72570 99583 72573
rect 183697 72570 183763 72573
rect 95732 72568 99583 72570
rect 95732 72512 99522 72568
rect 99578 72512 99583 72568
rect 95732 72510 99583 72512
rect 179820 72568 183763 72570
rect 179820 72512 183702 72568
rect 183758 72512 183763 72568
rect 179820 72510 183763 72512
rect 99517 72507 99583 72510
rect 183697 72507 183763 72510
rect 183697 71346 183763 71349
rect 179820 71344 183763 71346
rect 179820 71288 183702 71344
rect 183758 71288 183763 71344
rect 95702 71074 95762 71288
rect 179820 71286 183763 71288
rect 183697 71283 183763 71286
rect 99517 71074 99583 71077
rect 95702 71072 99583 71074
rect 95702 71016 99522 71072
rect 99578 71016 99583 71072
rect 95702 71014 99583 71016
rect 99517 71011 99583 71014
rect 190781 70802 190847 70805
rect 190781 70800 193988 70802
rect 190781 70744 190786 70800
rect 190842 70744 193988 70800
rect 190781 70742 193988 70744
rect 190781 70739 190847 70742
rect 106693 70394 106759 70397
rect 106693 70392 109900 70394
rect 106693 70336 106698 70392
rect 106754 70336 109900 70392
rect 106693 70334 109900 70336
rect 106693 70331 106759 70334
rect 182869 70122 182935 70125
rect 179820 70120 182935 70122
rect 179820 70064 182874 70120
rect 182930 70064 182935 70120
rect 23617 69850 23683 69853
rect 95702 69850 95762 70064
rect 179820 70062 182935 70064
rect 182869 70059 182935 70062
rect 99517 69850 99583 69853
rect 128497 69850 128563 69853
rect 212677 69850 212743 69853
rect 23617 69848 25996 69850
rect 23617 69792 23622 69848
rect 23678 69792 25996 69848
rect 23617 69790 25996 69792
rect 95702 69848 99583 69850
rect 95702 69792 99522 69848
rect 99578 69792 99583 69848
rect 95702 69790 99583 69792
rect 125724 69848 128563 69850
rect 125724 69792 128502 69848
rect 128558 69792 128563 69848
rect 125724 69790 128563 69792
rect 209812 69848 212743 69850
rect 209812 69792 212682 69848
rect 212738 69792 212743 69848
rect 209812 69790 212743 69792
rect 23617 69787 23683 69790
rect 99517 69787 99583 69790
rect 128497 69787 128563 69790
rect 212677 69787 212743 69790
rect 183053 68898 183119 68901
rect 179820 68896 183119 68898
rect 179820 68840 183058 68896
rect 183114 68840 183119 68896
rect 95702 68354 95762 68840
rect 179820 68838 183119 68840
rect 183053 68835 183119 68838
rect 190965 68762 191031 68765
rect 190965 68760 193988 68762
rect 190965 68704 190970 68760
rect 191026 68704 193988 68760
rect 190965 68702 193988 68704
rect 190965 68699 191031 68702
rect 98965 68354 99031 68357
rect 95702 68352 99031 68354
rect 95702 68296 98970 68352
rect 99026 68296 99031 68352
rect 95702 68294 99031 68296
rect 98965 68291 99031 68294
rect 106601 67946 106667 67949
rect 106601 67944 109900 67946
rect 106601 67888 106606 67944
rect 106662 67888 109900 67944
rect 106601 67886 109900 67888
rect 106601 67883 106667 67886
rect 9896 67810 10376 67840
rect 13262 67810 13268 67812
rect 9896 67750 13268 67810
rect 9896 67720 10376 67750
rect 13262 67748 13268 67750
rect 13332 67748 13338 67812
rect 183145 67674 183211 67677
rect 179820 67672 183211 67674
rect 179820 67616 183150 67672
rect 183206 67616 183211 67672
rect 95702 67130 95762 67616
rect 179820 67614 183211 67616
rect 183145 67611 183211 67614
rect 99057 67130 99123 67133
rect 95702 67128 99123 67130
rect 95702 67072 99062 67128
rect 99118 67072 99123 67128
rect 95702 67070 99123 67072
rect 99057 67067 99123 67070
rect 191333 66858 191399 66861
rect 191333 66856 193988 66858
rect 191333 66800 191338 66856
rect 191394 66800 193988 66856
rect 191333 66798 193988 66800
rect 191333 66795 191399 66798
rect 53333 66586 53399 66589
rect 136869 66586 136935 66589
rect 137973 66586 138039 66589
rect 53333 66584 55988 66586
rect 53333 66528 53338 66584
rect 53394 66528 55988 66584
rect 53333 66526 55988 66528
rect 136869 66584 140076 66586
rect 136869 66528 136874 66584
rect 136930 66528 137978 66584
rect 138034 66528 140076 66584
rect 136869 66526 140076 66528
rect 53333 66523 53399 66526
rect 136869 66523 136935 66526
rect 137973 66523 138039 66526
rect 183237 66450 183303 66453
rect 179820 66448 183303 66450
rect 179820 66392 183242 66448
rect 183298 66392 183303 66448
rect 95702 65906 95762 66392
rect 179820 66390 183303 66392
rect 183237 66387 183303 66390
rect 99149 65906 99215 65909
rect 95702 65904 99215 65906
rect 95702 65848 99154 65904
rect 99210 65848 99215 65904
rect 95702 65846 99215 65848
rect 99149 65843 99215 65846
rect 106509 65634 106575 65637
rect 106509 65632 109900 65634
rect 106509 65576 106514 65632
rect 106570 65576 109900 65632
rect 106509 65574 109900 65576
rect 106509 65571 106575 65574
rect 183329 65226 183395 65229
rect 179820 65224 183395 65226
rect 179820 65168 183334 65224
rect 183390 65168 183395 65224
rect 44409 64818 44475 64821
rect 41820 64816 44475 64818
rect 41820 64760 44414 64816
rect 44470 64760 44475 64816
rect 41820 64758 44475 64760
rect 44409 64755 44475 64758
rect 95702 64682 95762 65168
rect 179820 65166 183395 65168
rect 183329 65163 183395 65166
rect 191517 64818 191583 64821
rect 191517 64816 193988 64818
rect 191517 64760 191522 64816
rect 191578 64760 193988 64816
rect 191517 64758 193988 64760
rect 191517 64755 191583 64758
rect 99241 64682 99307 64685
rect 95702 64680 99307 64682
rect 95702 64624 99246 64680
rect 99302 64624 99307 64680
rect 95702 64622 99307 64624
rect 99241 64619 99307 64622
rect 183605 64002 183671 64005
rect 179820 64000 183671 64002
rect 179820 63944 183610 64000
rect 183666 63944 183671 64000
rect 95702 63458 95762 63944
rect 179820 63942 183671 63944
rect 183605 63939 183671 63942
rect 99517 63458 99583 63461
rect 95702 63456 99583 63458
rect 95702 63400 99522 63456
rect 99578 63400 99583 63456
rect 95702 63398 99583 63400
rect 99517 63395 99583 63398
rect 106601 63322 106667 63325
rect 106601 63320 109900 63322
rect 106601 63264 106606 63320
rect 106662 63264 109900 63320
rect 106601 63262 109900 63264
rect 106601 63259 106667 63262
rect 23617 63186 23683 63189
rect 212350 63186 212356 63188
rect 23617 63184 25996 63186
rect 23617 63128 23622 63184
rect 23678 63128 25996 63184
rect 23617 63126 25996 63128
rect 209812 63126 212356 63186
rect 23617 63123 23683 63126
rect 212350 63124 212356 63126
rect 212420 63124 212426 63188
rect 99333 62778 99399 62781
rect 183421 62778 183487 62781
rect 95732 62776 99399 62778
rect 95732 62720 99338 62776
rect 99394 62720 99399 62776
rect 95732 62718 99399 62720
rect 179820 62776 183487 62778
rect 179820 62720 183426 62776
rect 183482 62720 183487 62776
rect 179820 62718 183487 62720
rect 99333 62715 99399 62718
rect 183421 62715 183487 62718
rect 189953 62778 190019 62781
rect 189953 62776 193988 62778
rect 189953 62720 189958 62776
rect 190014 62720 193988 62776
rect 189953 62718 193988 62720
rect 189953 62715 190019 62718
rect 99517 61554 99583 61557
rect 183697 61554 183763 61557
rect 95732 61552 99583 61554
rect 95732 61496 99522 61552
rect 99578 61496 99583 61552
rect 95732 61494 99583 61496
rect 179820 61552 183763 61554
rect 179820 61496 183702 61552
rect 183758 61496 183763 61552
rect 179820 61494 183763 61496
rect 99517 61491 99583 61494
rect 183697 61491 183763 61494
rect 107153 61010 107219 61013
rect 107153 61008 109900 61010
rect 107153 60952 107158 61008
rect 107214 60952 109900 61008
rect 107153 60950 109900 60952
rect 107153 60947 107219 60950
rect 191977 60874 192043 60877
rect 191977 60872 193988 60874
rect 191977 60816 191982 60872
rect 192038 60816 193988 60872
rect 191977 60814 193988 60816
rect 191977 60811 192043 60814
rect 182685 60466 182751 60469
rect 179820 60464 182751 60466
rect 179820 60408 182690 60464
rect 182746 60408 182751 60464
rect 95702 59922 95762 60408
rect 179820 60406 182751 60408
rect 182685 60403 182751 60406
rect 100253 59922 100319 59925
rect 95702 59920 100319 59922
rect 95702 59864 100258 59920
rect 100314 59864 100319 59920
rect 95702 59862 100319 59864
rect 100253 59859 100319 59862
rect 59221 58426 59287 58429
rect 140222 58426 140228 58428
rect 59221 58424 140228 58426
rect 59221 58368 59226 58424
rect 59282 58368 140228 58424
rect 59221 58366 140228 58368
rect 59221 58363 59287 58366
rect 140222 58364 140228 58366
rect 140292 58364 140298 58428
rect 55950 58228 55956 58292
rect 56020 58290 56026 58292
rect 79185 58290 79251 58293
rect 56020 58288 79251 58290
rect 56020 58232 79190 58288
rect 79246 58232 79251 58288
rect 56020 58230 79251 58232
rect 56020 58228 56026 58230
rect 79185 58227 79251 58230
rect 222245 48090 222311 48093
rect 225416 48090 225896 48120
rect 222245 48088 225896 48090
rect 222245 48032 222250 48088
rect 222306 48032 225896 48088
rect 222245 48030 225896 48032
rect 222245 48027 222311 48030
rect 225416 48000 225896 48030
rect 50389 46866 50455 46869
rect 47862 46864 50455 46866
rect 47862 46808 50394 46864
rect 50450 46808 50455 46864
rect 47862 46806 50455 46808
rect 47862 46224 47922 46806
rect 50389 46803 50455 46806
rect 64966 46804 64972 46868
rect 65036 46866 65042 46868
rect 79277 46866 79343 46869
rect 65036 46864 79343 46866
rect 65036 46808 79282 46864
rect 79338 46808 79343 46864
rect 65036 46806 79343 46808
rect 65036 46804 65042 46806
rect 79277 46803 79343 46806
rect 159542 46804 159548 46868
rect 159612 46866 159618 46868
rect 164745 46866 164811 46869
rect 159612 46864 164811 46866
rect 159612 46808 164750 46864
rect 164806 46808 164811 46864
rect 159612 46806 164811 46808
rect 159612 46804 159618 46806
rect 164745 46803 164811 46806
rect 63494 46668 63500 46732
rect 63564 46730 63570 46732
rect 80749 46730 80815 46733
rect 63564 46728 80815 46730
rect 63564 46672 80754 46728
rect 80810 46672 80815 46728
rect 63564 46670 80815 46672
rect 63564 46668 63570 46670
rect 80749 46667 80815 46670
rect 149054 46668 149060 46732
rect 149124 46730 149130 46732
rect 161893 46730 161959 46733
rect 149124 46728 161959 46730
rect 149124 46672 161898 46728
rect 161954 46672 161959 46728
rect 149124 46670 161959 46672
rect 149124 46668 149130 46670
rect 161893 46667 161959 46670
rect 62206 46532 62212 46596
rect 62276 46594 62282 46596
rect 73389 46594 73455 46597
rect 62276 46592 73455 46594
rect 62276 46536 73394 46592
rect 73450 46536 73455 46592
rect 62276 46534 73455 46536
rect 62276 46532 62282 46534
rect 73389 46531 73455 46534
rect 146294 46532 146300 46596
rect 146364 46594 146370 46596
rect 158949 46594 159015 46597
rect 146364 46592 159015 46594
rect 146364 46536 158954 46592
rect 159010 46536 159015 46592
rect 146364 46534 159015 46536
rect 146364 46532 146370 46534
rect 158949 46531 159015 46534
rect 63126 46396 63132 46460
rect 63196 46458 63202 46460
rect 76333 46458 76399 46461
rect 63196 46456 76399 46458
rect 63196 46400 76338 46456
rect 76394 46400 76399 46456
rect 63196 46398 76399 46400
rect 63196 46396 63202 46398
rect 76333 46395 76399 46398
rect 63310 46260 63316 46324
rect 63380 46322 63386 46324
rect 74861 46322 74927 46325
rect 63380 46320 74927 46322
rect 63380 46264 74866 46320
rect 74922 46264 74927 46320
rect 63380 46262 74927 46264
rect 63380 46260 63386 46262
rect 74861 46259 74927 46262
rect 85717 46322 85783 46325
rect 89806 46322 89812 46324
rect 85717 46320 89812 46322
rect 85717 46264 85722 46320
rect 85778 46264 89812 46320
rect 85717 46262 89812 46264
rect 85717 46259 85783 46262
rect 89806 46260 89812 46262
rect 89876 46260 89882 46324
rect 64782 46124 64788 46188
rect 64852 46186 64858 46188
rect 77805 46186 77871 46189
rect 64852 46184 77871 46186
rect 64852 46128 77810 46184
rect 77866 46128 77871 46184
rect 64852 46126 77871 46128
rect 64852 46124 64858 46126
rect 77805 46123 77871 46126
rect 87097 46186 87163 46189
rect 89070 46186 89076 46188
rect 87097 46184 89076 46186
rect 87097 46128 87102 46184
rect 87158 46128 89076 46184
rect 87097 46126 89076 46128
rect 87097 46123 87163 46126
rect 89070 46124 89076 46126
rect 89140 46124 89146 46188
rect 101173 46186 101239 46189
rect 103982 46186 104042 46496
rect 131766 46458 131826 46496
rect 134753 46458 134819 46461
rect 131766 46456 134819 46458
rect 131766 46400 134758 46456
rect 134814 46400 134819 46456
rect 131766 46398 134819 46400
rect 134753 46395 134819 46398
rect 147766 46396 147772 46460
rect 147836 46458 147842 46460
rect 160329 46458 160395 46461
rect 147836 46456 160395 46458
rect 147836 46400 160334 46456
rect 160390 46400 160395 46456
rect 147836 46398 160395 46400
rect 147836 46396 147842 46398
rect 160329 46395 160395 46398
rect 146110 46260 146116 46324
rect 146180 46322 146186 46324
rect 157569 46322 157635 46325
rect 163273 46322 163339 46325
rect 146180 46320 157635 46322
rect 146180 46264 157574 46320
rect 157630 46264 157635 46320
rect 146180 46262 157635 46264
rect 146180 46260 146186 46262
rect 157569 46259 157635 46262
rect 157710 46320 163339 46322
rect 157710 46264 163278 46320
rect 163334 46264 163339 46320
rect 157710 46262 163339 46264
rect 138341 46186 138407 46189
rect 101173 46184 104042 46186
rect 101173 46128 101178 46184
rect 101234 46128 104042 46184
rect 138206 46184 138407 46186
rect 101173 46126 104042 46128
rect 138065 46152 138131 46155
rect 138206 46152 138346 46184
rect 138065 46150 138346 46152
rect 101173 46123 101239 46126
rect 138065 46094 138070 46150
rect 138126 46128 138346 46150
rect 138402 46128 138407 46184
rect 138126 46126 138407 46128
rect 138126 46094 138266 46126
rect 138341 46123 138407 46126
rect 147030 46124 147036 46188
rect 147100 46186 147106 46188
rect 154257 46186 154323 46189
rect 147100 46184 154323 46186
rect 147100 46128 154262 46184
rect 154318 46128 154323 46184
rect 147100 46126 154323 46128
rect 147100 46124 147106 46126
rect 154257 46123 154323 46126
rect 138065 46092 138266 46094
rect 138065 46089 138131 46092
rect 154942 45988 154948 46052
rect 155012 46050 155018 46052
rect 157710 46050 157770 46262
rect 163273 46259 163339 46262
rect 169897 46322 169963 46325
rect 173158 46322 173164 46324
rect 169897 46320 173164 46322
rect 169897 46264 169902 46320
rect 169958 46264 173164 46320
rect 169897 46262 173164 46264
rect 169897 46259 169963 46262
rect 173158 46260 173164 46262
rect 173228 46260 173234 46324
rect 171093 46186 171159 46189
rect 173526 46186 173532 46188
rect 171093 46184 173532 46186
rect 171093 46128 171098 46184
rect 171154 46128 173532 46184
rect 171093 46126 173532 46128
rect 171093 46123 171159 46126
rect 173526 46124 173532 46126
rect 173596 46124 173602 46188
rect 185813 46186 185879 46189
rect 187886 46186 187946 46496
rect 185813 46184 187946 46186
rect 185813 46128 185818 46184
rect 185874 46128 187946 46184
rect 185813 46126 187946 46128
rect 185813 46123 185879 46126
rect 155012 45990 157770 46050
rect 155012 45988 155018 45990
rect 47862 45234 47922 45680
rect 100989 45506 101055 45509
rect 103982 45506 104042 45952
rect 100989 45504 104042 45506
rect 100989 45448 100994 45504
rect 101050 45448 104042 45504
rect 100989 45446 104042 45448
rect 131766 45506 131826 45952
rect 134845 45506 134911 45509
rect 131766 45504 134911 45506
rect 131766 45448 134850 45504
rect 134906 45448 134911 45504
rect 131766 45446 134911 45448
rect 100989 45443 101055 45446
rect 134845 45443 134911 45446
rect 185169 45506 185235 45509
rect 187886 45506 187946 45952
rect 185169 45504 187946 45506
rect 185169 45448 185174 45504
rect 185230 45448 187946 45504
rect 185169 45446 187946 45448
rect 185169 45443 185235 45446
rect 51309 45234 51375 45237
rect 47862 45232 51375 45234
rect 47862 45176 51314 45232
rect 51370 45176 51375 45232
rect 47862 45174 51375 45176
rect 51309 45171 51375 45174
rect 47862 44826 47922 45000
rect 101265 44962 101331 44965
rect 103982 44962 104042 45272
rect 131766 45098 131826 45272
rect 134293 45098 134359 45101
rect 131766 45096 134359 45098
rect 131766 45040 134298 45096
rect 134354 45040 134359 45096
rect 131766 45038 134359 45040
rect 134293 45035 134359 45038
rect 101265 44960 104042 44962
rect 101265 44904 101270 44960
rect 101326 44904 104042 44960
rect 101265 44902 104042 44904
rect 185445 44962 185511 44965
rect 187886 44962 187946 45272
rect 185445 44960 187946 44962
rect 185445 44904 185450 44960
rect 185506 44904 187946 44960
rect 185445 44902 187946 44904
rect 101265 44899 101331 44902
rect 185445 44899 185511 44902
rect 51217 44826 51283 44829
rect 47862 44824 51283 44826
rect 47862 44768 51222 44824
rect 51278 44768 51283 44824
rect 47862 44766 51283 44768
rect 51217 44763 51283 44766
rect 101081 44826 101147 44829
rect 134753 44826 134819 44829
rect 101081 44824 104042 44826
rect 101081 44768 101086 44824
rect 101142 44768 104042 44824
rect 101081 44766 104042 44768
rect 101081 44763 101147 44766
rect 103982 44732 104042 44766
rect 131766 44824 134819 44826
rect 131766 44768 134758 44824
rect 134814 44768 134819 44824
rect 131766 44766 134819 44768
rect 131766 44728 131826 44766
rect 134753 44763 134819 44766
rect 185537 44826 185603 44829
rect 185537 44824 187946 44826
rect 185537 44768 185542 44824
rect 185598 44768 187946 44824
rect 185537 44766 187946 44768
rect 185537 44763 185603 44766
rect 187886 44728 187946 44766
rect 172933 44690 172999 44693
rect 173894 44690 173900 44692
rect 172933 44688 173900 44690
rect 172933 44632 172938 44688
rect 172994 44632 173900 44688
rect 172933 44630 173900 44632
rect 172933 44627 172999 44630
rect 173894 44628 173900 44630
rect 173964 44628 173970 44692
rect 9896 44146 10376 44176
rect 13313 44146 13379 44149
rect 9896 44144 13379 44146
rect 9896 44088 13318 44144
rect 13374 44088 13379 44144
rect 9896 44086 13379 44088
rect 47862 44146 47922 44456
rect 58209 44418 58275 44421
rect 93997 44418 94063 44421
rect 58209 44416 60956 44418
rect 58209 44360 58214 44416
rect 58270 44360 60956 44416
rect 58209 44358 60956 44360
rect 90764 44416 94063 44418
rect 90764 44360 94002 44416
rect 94058 44360 94063 44416
rect 90764 44358 94063 44360
rect 58209 44355 58275 44358
rect 93997 44355 94063 44358
rect 142573 44418 142639 44421
rect 177717 44418 177783 44421
rect 142573 44416 145044 44418
rect 142573 44360 142578 44416
rect 142634 44360 145044 44416
rect 142573 44358 145044 44360
rect 174852 44416 177783 44418
rect 174852 44360 177722 44416
rect 177778 44360 177783 44416
rect 174852 44358 177783 44360
rect 142573 44355 142639 44358
rect 177717 44355 177783 44358
rect 93905 44282 93971 44285
rect 90734 44280 93971 44282
rect 90734 44224 93910 44280
rect 93966 44224 93971 44280
rect 90734 44222 93971 44224
rect 51217 44146 51283 44149
rect 47862 44144 51283 44146
rect 47862 44088 51222 44144
rect 51278 44088 51283 44144
rect 47862 44086 51283 44088
rect 9896 44056 10376 44086
rect 13313 44083 13379 44086
rect 51217 44083 51283 44086
rect 90734 43912 90794 44222
rect 93905 44219 93971 44222
rect 142389 44282 142455 44285
rect 142389 44280 145074 44282
rect 142389 44224 142394 44280
rect 142450 44224 145074 44280
rect 142389 44222 145074 44224
rect 142389 44219 142455 44222
rect 47862 43738 47922 43912
rect 58301 43874 58367 43877
rect 58301 43872 60956 43874
rect 58301 43816 58306 43872
rect 58362 43816 60956 43872
rect 58301 43814 60956 43816
rect 58301 43811 58367 43814
rect 50021 43738 50087 43741
rect 47862 43736 50087 43738
rect 47862 43680 50026 43736
rect 50082 43680 50087 43736
rect 47862 43678 50087 43680
rect 50021 43675 50087 43678
rect 100989 43738 101055 43741
rect 103982 43738 104042 44048
rect 131766 43874 131826 44048
rect 145014 43912 145074 44222
rect 134753 43874 134819 43877
rect 177717 43874 177783 43877
rect 131766 43872 134819 43874
rect 131766 43816 134758 43872
rect 134814 43816 134819 43872
rect 131766 43814 134819 43816
rect 174852 43872 177783 43874
rect 174852 43816 177722 43872
rect 177778 43816 177783 43872
rect 174852 43814 177783 43816
rect 134753 43811 134819 43814
rect 177717 43811 177783 43814
rect 100989 43736 104042 43738
rect 100989 43680 100994 43736
rect 101050 43680 104042 43736
rect 100989 43678 104042 43680
rect 185169 43738 185235 43741
rect 187886 43738 187946 44048
rect 185169 43736 187946 43738
rect 185169 43680 185174 43736
rect 185230 43680 187946 43736
rect 185169 43678 187946 43680
rect 100989 43675 101055 43678
rect 185169 43675 185235 43678
rect 100805 43466 100871 43469
rect 103982 43466 104042 43504
rect 100805 43464 104042 43466
rect 100805 43408 100810 43464
rect 100866 43408 104042 43464
rect 100805 43406 104042 43408
rect 131766 43466 131826 43504
rect 134753 43466 134819 43469
rect 131766 43464 134819 43466
rect 131766 43408 134758 43464
rect 134814 43408 134819 43464
rect 131766 43406 134819 43408
rect 100805 43403 100871 43406
rect 134753 43403 134819 43406
rect 184985 43466 185051 43469
rect 187886 43466 187946 43504
rect 184985 43464 187946 43466
rect 184985 43408 184990 43464
rect 185046 43408 187946 43464
rect 184985 43406 187946 43408
rect 184985 43403 185051 43406
rect 47862 42922 47922 43232
rect 58209 43194 58275 43197
rect 93997 43194 94063 43197
rect 58209 43192 60956 43194
rect 58209 43136 58214 43192
rect 58270 43136 60956 43192
rect 58209 43134 60956 43136
rect 90764 43192 94063 43194
rect 90764 43136 94002 43192
rect 94058 43136 94063 43192
rect 90764 43134 94063 43136
rect 58209 43131 58275 43134
rect 93997 43131 94063 43134
rect 142481 43194 142547 43197
rect 177717 43194 177783 43197
rect 142481 43192 145044 43194
rect 142481 43136 142486 43192
rect 142542 43136 145044 43192
rect 142481 43134 145044 43136
rect 174852 43192 177783 43194
rect 174852 43136 177722 43192
rect 177778 43136 177783 43192
rect 174852 43134 177783 43136
rect 142481 43131 142547 43134
rect 177717 43131 177783 43134
rect 142665 43058 142731 43061
rect 142665 43056 145074 43058
rect 142665 43000 142670 43056
rect 142726 43000 145074 43056
rect 142665 42998 145074 43000
rect 142665 42995 142731 42998
rect 50205 42922 50271 42925
rect 93905 42922 93971 42925
rect 47862 42920 50271 42922
rect 47862 42864 50210 42920
rect 50266 42864 50271 42920
rect 47862 42862 50271 42864
rect 50205 42859 50271 42862
rect 90734 42920 93971 42922
rect 90734 42864 93910 42920
rect 93966 42864 93971 42920
rect 90734 42862 93971 42864
rect 90734 42688 90794 42862
rect 93905 42859 93971 42862
rect 47862 42378 47922 42688
rect 58301 42650 58367 42653
rect 58301 42648 60956 42650
rect 58301 42592 58306 42648
rect 58362 42592 60956 42648
rect 58301 42590 60956 42592
rect 58301 42587 58367 42590
rect 93997 42514 94063 42517
rect 90734 42512 94063 42514
rect 90734 42456 94002 42512
rect 94058 42456 94063 42512
rect 90734 42454 94063 42456
rect 51125 42378 51191 42381
rect 47862 42376 51191 42378
rect 47862 42320 51130 42376
rect 51186 42320 51191 42376
rect 47862 42318 51191 42320
rect 51125 42315 51191 42318
rect 90734 42144 90794 42454
rect 93997 42451 94063 42454
rect 100989 42514 101055 42517
rect 103982 42514 104042 42824
rect 131766 42650 131826 42824
rect 145014 42688 145074 42998
rect 134753 42650 134819 42653
rect 177625 42650 177691 42653
rect 131766 42648 134819 42650
rect 131766 42592 134758 42648
rect 134814 42592 134819 42648
rect 131766 42590 134819 42592
rect 174852 42648 177691 42650
rect 174852 42592 177630 42648
rect 177686 42592 177691 42648
rect 174852 42590 177691 42592
rect 134753 42587 134819 42590
rect 177625 42587 177691 42590
rect 100989 42512 104042 42514
rect 100989 42456 100994 42512
rect 101050 42456 104042 42512
rect 100989 42454 104042 42456
rect 143125 42514 143191 42517
rect 185169 42514 185235 42517
rect 187886 42514 187946 42824
rect 143125 42512 145074 42514
rect 143125 42456 143130 42512
rect 143186 42456 145074 42512
rect 143125 42454 145074 42456
rect 100989 42451 101055 42454
rect 143125 42451 143191 42454
rect 51217 42106 51283 42109
rect 47862 42104 51283 42106
rect 47862 42048 51222 42104
rect 51278 42048 51283 42104
rect 47862 42046 51283 42048
rect 47862 42008 47922 42046
rect 51217 42043 51283 42046
rect 58209 42106 58275 42109
rect 100897 42106 100963 42109
rect 103982 42106 104042 42280
rect 58209 42104 60956 42106
rect 58209 42048 58214 42104
rect 58270 42048 60956 42104
rect 58209 42046 60956 42048
rect 100897 42104 104042 42106
rect 100897 42048 100902 42104
rect 100958 42048 104042 42104
rect 100897 42046 104042 42048
rect 131766 42106 131826 42280
rect 145014 42144 145074 42454
rect 185169 42512 187946 42514
rect 185169 42456 185174 42512
rect 185230 42456 187946 42512
rect 185169 42454 187946 42456
rect 185169 42451 185235 42454
rect 134753 42106 134819 42109
rect 177717 42106 177783 42109
rect 131766 42104 134819 42106
rect 131766 42048 134758 42104
rect 134814 42048 134819 42104
rect 131766 42046 134819 42048
rect 174852 42104 177783 42106
rect 174852 42048 177722 42104
rect 177778 42048 177783 42104
rect 174852 42046 177783 42048
rect 58209 42043 58275 42046
rect 100897 42043 100963 42046
rect 134753 42043 134819 42046
rect 177717 42043 177783 42046
rect 185077 42106 185143 42109
rect 187886 42106 187946 42280
rect 185077 42104 187946 42106
rect 185077 42048 185082 42104
rect 185138 42048 187946 42104
rect 185077 42046 187946 42048
rect 185077 42043 185143 42046
rect 143493 41970 143559 41973
rect 143493 41968 145074 41970
rect 143493 41912 143498 41968
rect 143554 41912 145074 41968
rect 143493 41910 145074 41912
rect 143493 41907 143559 41910
rect 93997 41698 94063 41701
rect 90734 41696 94063 41698
rect 90734 41640 94002 41696
rect 94058 41640 94063 41696
rect 90734 41638 94063 41640
rect 90734 41464 90794 41638
rect 93997 41635 94063 41638
rect 47862 41154 47922 41464
rect 58209 41426 58275 41429
rect 58209 41424 60956 41426
rect 58209 41368 58214 41424
rect 58270 41368 60956 41424
rect 58209 41366 60956 41368
rect 58209 41363 58275 41366
rect 92709 41290 92775 41293
rect 90734 41288 92775 41290
rect 90734 41232 92714 41288
rect 92770 41232 92775 41288
rect 90734 41230 92775 41232
rect 51125 41154 51191 41157
rect 47862 41152 51191 41154
rect 47862 41096 51130 41152
rect 51186 41096 51191 41152
rect 47862 41094 51191 41096
rect 51125 41091 51191 41094
rect 90734 40920 90794 41230
rect 92709 41227 92775 41230
rect 100989 41290 101055 41293
rect 103982 41290 104042 41600
rect 100989 41288 104042 41290
rect 100989 41232 100994 41288
rect 101050 41232 104042 41288
rect 100989 41230 104042 41232
rect 131766 41290 131826 41600
rect 145014 41464 145074 41910
rect 177717 41426 177783 41429
rect 174852 41424 177783 41426
rect 174852 41368 177722 41424
rect 177778 41368 177783 41424
rect 174852 41366 177783 41368
rect 177717 41363 177783 41366
rect 134661 41290 134727 41293
rect 131766 41288 134727 41290
rect 131766 41232 134666 41288
rect 134722 41232 134727 41288
rect 131766 41230 134727 41232
rect 100989 41227 101055 41230
rect 134661 41227 134727 41230
rect 142757 41290 142823 41293
rect 185169 41290 185235 41293
rect 187886 41290 187946 41600
rect 142757 41288 145074 41290
rect 142757 41232 142762 41288
rect 142818 41232 145074 41288
rect 142757 41230 145074 41232
rect 142757 41227 142823 41230
rect 47862 40882 47922 40920
rect 51217 40882 51283 40885
rect 47862 40880 51283 40882
rect 47862 40824 51222 40880
rect 51278 40824 51283 40880
rect 47862 40822 51283 40824
rect 51217 40819 51283 40822
rect 58301 40882 58367 40885
rect 58301 40880 60956 40882
rect 58301 40824 58306 40880
rect 58362 40824 60956 40880
rect 58301 40822 60956 40824
rect 58301 40819 58367 40822
rect 100805 40610 100871 40613
rect 103982 40610 104042 41056
rect 131766 41018 131826 41056
rect 134753 41018 134819 41021
rect 131766 41016 134819 41018
rect 131766 40960 134758 41016
rect 134814 40960 134819 41016
rect 131766 40958 134819 40960
rect 134753 40955 134819 40958
rect 145014 40920 145074 41230
rect 185169 41288 187946 41290
rect 185169 41232 185174 41288
rect 185230 41232 187946 41288
rect 185169 41230 187946 41232
rect 185169 41227 185235 41230
rect 177625 40882 177691 40885
rect 174852 40880 177691 40882
rect 174852 40824 177630 40880
rect 177686 40824 177691 40880
rect 174852 40822 177691 40824
rect 177625 40819 177691 40822
rect 100805 40608 104042 40610
rect 100805 40552 100810 40608
rect 100866 40552 104042 40608
rect 100805 40550 104042 40552
rect 184985 40610 185051 40613
rect 187886 40610 187946 41056
rect 184985 40608 187946 40610
rect 184985 40552 184990 40608
rect 185046 40552 187946 40608
rect 184985 40550 187946 40552
rect 100805 40547 100871 40550
rect 184985 40547 185051 40550
rect 47862 39930 47922 40240
rect 58209 40202 58275 40205
rect 93997 40202 94063 40205
rect 58209 40200 60956 40202
rect 58209 40144 58214 40200
rect 58270 40144 60956 40200
rect 58209 40142 60956 40144
rect 90764 40200 94063 40202
rect 90764 40144 94002 40200
rect 94058 40144 94063 40200
rect 90764 40142 94063 40144
rect 58209 40139 58275 40142
rect 93997 40139 94063 40142
rect 92709 40066 92775 40069
rect 90734 40064 92775 40066
rect 90734 40008 92714 40064
rect 92770 40008 92775 40064
rect 90734 40006 92775 40008
rect 51125 39930 51191 39933
rect 47862 39928 51191 39930
rect 47862 39872 51130 39928
rect 51186 39872 51191 39928
rect 47862 39870 51191 39872
rect 51125 39867 51191 39870
rect 90734 39696 90794 40006
rect 92709 40003 92775 40006
rect 101081 40066 101147 40069
rect 103982 40066 104042 40376
rect 101081 40064 104042 40066
rect 101081 40008 101086 40064
rect 101142 40008 104042 40064
rect 101081 40006 104042 40008
rect 131766 40066 131826 40376
rect 143677 40202 143743 40205
rect 177717 40202 177783 40205
rect 143677 40200 145044 40202
rect 143677 40144 143682 40200
rect 143738 40144 145044 40200
rect 143677 40142 145044 40144
rect 174852 40200 177783 40202
rect 174852 40144 177722 40200
rect 177778 40144 177783 40200
rect 174852 40142 177783 40144
rect 143677 40139 143743 40142
rect 177717 40139 177783 40142
rect 134569 40066 134635 40069
rect 131766 40064 134635 40066
rect 131766 40008 134574 40064
rect 134630 40008 134635 40064
rect 131766 40006 134635 40008
rect 101081 40003 101147 40006
rect 134569 40003 134635 40006
rect 142389 40066 142455 40069
rect 185261 40066 185327 40069
rect 187886 40066 187946 40376
rect 142389 40064 145074 40066
rect 142389 40008 142394 40064
rect 142450 40008 145074 40064
rect 142389 40006 145074 40008
rect 142389 40003 142455 40006
rect 18097 39386 18163 39389
rect 19894 39386 19954 39560
rect 47862 39522 47922 39696
rect 58301 39658 58367 39661
rect 58301 39656 60956 39658
rect 58301 39600 58306 39656
rect 58362 39600 60956 39656
rect 58301 39598 60956 39600
rect 58301 39595 58367 39598
rect 51217 39522 51283 39525
rect 47862 39520 51283 39522
rect 47862 39464 51222 39520
rect 51278 39464 51283 39520
rect 47862 39462 51283 39464
rect 51217 39459 51283 39462
rect 18097 39384 19954 39386
rect 18097 39328 18102 39384
rect 18158 39328 19954 39384
rect 18097 39326 19954 39328
rect 100989 39386 101055 39389
rect 103982 39386 104042 39832
rect 131766 39522 131826 39832
rect 145014 39696 145074 40006
rect 185261 40064 187946 40066
rect 185261 40008 185266 40064
rect 185322 40008 187946 40064
rect 185261 40006 187946 40008
rect 185261 40003 185327 40006
rect 177257 39658 177323 39661
rect 174852 39656 177323 39658
rect 174852 39600 177262 39656
rect 177318 39600 177323 39656
rect 174852 39598 177323 39600
rect 177257 39595 177323 39598
rect 134661 39522 134727 39525
rect 131766 39520 134727 39522
rect 131766 39464 134666 39520
rect 134722 39464 134727 39520
rect 131766 39462 134727 39464
rect 134661 39459 134727 39462
rect 100989 39384 104042 39386
rect 100989 39328 100994 39384
rect 101050 39328 104042 39384
rect 100989 39326 104042 39328
rect 185169 39386 185235 39389
rect 187886 39386 187946 39832
rect 185169 39384 187946 39386
rect 185169 39328 185174 39384
rect 185230 39328 187946 39384
rect 185169 39326 187946 39328
rect 18097 39323 18163 39326
rect 100989 39323 101055 39326
rect 185169 39323 185235 39326
rect 47862 38842 47922 39152
rect 58209 39114 58275 39117
rect 93997 39114 94063 39117
rect 58209 39112 60956 39114
rect 58209 39056 58214 39112
rect 58270 39056 60956 39112
rect 58209 39054 60956 39056
rect 90764 39112 94063 39114
rect 90764 39056 94002 39112
rect 94058 39056 94063 39112
rect 90764 39054 94063 39056
rect 58209 39051 58275 39054
rect 93997 39051 94063 39054
rect 51217 38842 51283 38845
rect 47862 38840 51283 38842
rect 47862 38784 51222 38840
rect 51278 38784 51283 38840
rect 47862 38782 51283 38784
rect 51217 38779 51283 38782
rect 101081 38842 101147 38845
rect 103982 38842 104042 39152
rect 101081 38840 104042 38842
rect 101081 38784 101086 38840
rect 101142 38784 104042 38840
rect 101081 38782 104042 38784
rect 131766 38842 131826 39152
rect 142481 39114 142547 39117
rect 177717 39114 177783 39117
rect 142481 39112 145044 39114
rect 142481 39056 142486 39112
rect 142542 39056 145044 39112
rect 142481 39054 145044 39056
rect 174852 39112 177783 39114
rect 174852 39056 177722 39112
rect 177778 39056 177783 39112
rect 174852 39054 177783 39056
rect 142481 39051 142547 39054
rect 177717 39051 177783 39054
rect 142389 38978 142455 38981
rect 142389 38976 145074 38978
rect 142389 38920 142394 38976
rect 142450 38920 145074 38976
rect 142389 38918 145074 38920
rect 142389 38915 142455 38918
rect 134109 38842 134175 38845
rect 131766 38840 134175 38842
rect 131766 38784 134114 38840
rect 134170 38784 134175 38840
rect 131766 38782 134175 38784
rect 101081 38779 101147 38782
rect 134109 38779 134175 38782
rect 93905 38706 93971 38709
rect 90734 38704 93971 38706
rect 90734 38648 93910 38704
rect 93966 38648 93971 38704
rect 90734 38646 93971 38648
rect 90734 38472 90794 38646
rect 93905 38643 93971 38646
rect 47862 38162 47922 38472
rect 58393 38434 58459 38437
rect 58393 38432 60956 38434
rect 58393 38376 58398 38432
rect 58454 38376 60956 38432
rect 58393 38374 60956 38376
rect 58393 38371 58459 38374
rect 92893 38298 92959 38301
rect 90734 38296 92959 38298
rect 90734 38240 92898 38296
rect 92954 38240 92959 38296
rect 90734 38238 92959 38240
rect 51125 38162 51191 38165
rect 47862 38160 51191 38162
rect 47862 38104 51130 38160
rect 51186 38104 51191 38160
rect 47862 38102 51191 38104
rect 51125 38099 51191 38102
rect 90734 37928 90794 38238
rect 92893 38235 92959 38238
rect 100989 38298 101055 38301
rect 103982 38298 104042 38608
rect 100989 38296 104042 38298
rect 100989 38240 100994 38296
rect 101050 38240 104042 38296
rect 100989 38238 104042 38240
rect 131766 38298 131826 38608
rect 145014 38472 145074 38918
rect 185261 38842 185327 38845
rect 187886 38842 187946 39152
rect 185261 38840 187946 38842
rect 185261 38784 185266 38840
rect 185322 38784 187946 38840
rect 185261 38782 187946 38784
rect 185261 38779 185327 38782
rect 177441 38434 177507 38437
rect 174852 38432 177507 38434
rect 174852 38376 177446 38432
rect 177502 38376 177507 38432
rect 174852 38374 177507 38376
rect 177441 38371 177507 38374
rect 134293 38298 134359 38301
rect 131766 38296 134359 38298
rect 131766 38240 134298 38296
rect 134354 38240 134359 38296
rect 131766 38238 134359 38240
rect 100989 38235 101055 38238
rect 134293 38235 134359 38238
rect 142573 38298 142639 38301
rect 142573 38296 145074 38298
rect 142573 38240 142578 38296
rect 142634 38240 145074 38296
rect 142573 38238 145074 38240
rect 142573 38235 142639 38238
rect 134661 38026 134727 38029
rect 131766 38024 134727 38026
rect 131766 37968 134666 38024
rect 134722 37968 134727 38024
rect 131766 37966 134727 37968
rect 131766 37928 131826 37966
rect 134661 37963 134727 37966
rect 145014 37928 145074 38238
rect 185169 38162 185235 38165
rect 187886 38162 187946 38608
rect 185169 38160 187946 38162
rect 185169 38104 185174 38160
rect 185230 38104 187946 38160
rect 185169 38102 187946 38104
rect 185169 38099 185235 38102
rect 47862 37890 47922 37928
rect 51217 37890 51283 37893
rect 47862 37888 51283 37890
rect 47862 37832 51222 37888
rect 51278 37832 51283 37888
rect 47862 37830 51283 37832
rect 51217 37827 51283 37830
rect 58301 37890 58367 37893
rect 100805 37890 100871 37893
rect 103982 37890 104042 37928
rect 177349 37890 177415 37893
rect 58301 37888 60956 37890
rect 58301 37832 58306 37888
rect 58362 37832 60956 37888
rect 58301 37830 60956 37832
rect 100805 37888 104042 37890
rect 100805 37832 100810 37888
rect 100866 37832 104042 37888
rect 100805 37830 104042 37832
rect 174852 37888 177415 37890
rect 174852 37832 177354 37888
rect 177410 37832 177415 37888
rect 174852 37830 177415 37832
rect 58301 37827 58367 37830
rect 100805 37827 100871 37830
rect 177349 37827 177415 37830
rect 184985 37890 185051 37893
rect 187886 37890 187946 37928
rect 184985 37888 187946 37890
rect 184985 37832 184990 37888
rect 185046 37832 187946 37888
rect 184985 37830 187946 37832
rect 184985 37827 185051 37830
rect 142389 37754 142455 37757
rect 142389 37752 145074 37754
rect 142389 37696 142394 37752
rect 142450 37696 145074 37752
rect 142389 37694 145074 37696
rect 142389 37691 142455 37694
rect 93997 37618 94063 37621
rect 90734 37616 94063 37618
rect 90734 37560 94002 37616
rect 94058 37560 94063 37616
rect 90734 37558 94063 37560
rect 90734 37248 90794 37558
rect 93997 37555 94063 37558
rect 47862 36938 47922 37248
rect 58393 37210 58459 37213
rect 58393 37208 60956 37210
rect 58393 37152 58398 37208
rect 58454 37152 60956 37208
rect 58393 37150 60956 37152
rect 58393 37147 58459 37150
rect 93997 37074 94063 37077
rect 90734 37072 94063 37074
rect 90734 37016 94002 37072
rect 94058 37016 94063 37072
rect 90734 37014 94063 37016
rect 51125 36938 51191 36941
rect 47862 36936 51191 36938
rect 47862 36880 51130 36936
rect 51186 36880 51191 36936
rect 47862 36878 51191 36880
rect 51125 36875 51191 36878
rect 90734 36704 90794 37014
rect 93997 37011 94063 37014
rect 100989 36938 101055 36941
rect 103982 36938 104042 37384
rect 100989 36936 104042 36938
rect 100989 36880 100994 36936
rect 101050 36880 104042 36936
rect 100989 36878 104042 36880
rect 131766 36938 131826 37384
rect 145014 37248 145074 37694
rect 177441 37210 177507 37213
rect 174852 37208 177507 37210
rect 174852 37152 177446 37208
rect 177502 37152 177507 37208
rect 174852 37150 177507 37152
rect 177441 37147 177507 37150
rect 142481 37074 142547 37077
rect 142481 37072 145074 37074
rect 142481 37016 142486 37072
rect 142542 37016 145074 37072
rect 142481 37014 145074 37016
rect 142481 37011 142547 37014
rect 134661 36938 134727 36941
rect 131766 36936 134727 36938
rect 131766 36880 134666 36936
rect 134722 36880 134727 36936
rect 131766 36878 134727 36880
rect 100989 36875 101055 36878
rect 134661 36875 134727 36878
rect 145014 36704 145074 37014
rect 185169 36938 185235 36941
rect 187886 36938 187946 37384
rect 185169 36936 187946 36938
rect 185169 36880 185174 36936
rect 185230 36880 187946 36936
rect 185169 36878 187946 36880
rect 185169 36875 185235 36878
rect 47862 36666 47922 36704
rect 51217 36666 51283 36669
rect 47862 36664 51283 36666
rect 47862 36608 51222 36664
rect 51278 36608 51283 36664
rect 47862 36606 51283 36608
rect 51217 36603 51283 36606
rect 58209 36666 58275 36669
rect 58209 36664 60956 36666
rect 58209 36608 58214 36664
rect 58270 36608 60956 36664
rect 58209 36606 60956 36608
rect 58209 36603 58275 36606
rect 100897 36530 100963 36533
rect 103982 36530 104042 36704
rect 131766 36666 131826 36704
rect 134385 36666 134451 36669
rect 177717 36666 177783 36669
rect 131766 36664 134451 36666
rect 131766 36608 134390 36664
rect 134446 36608 134451 36664
rect 131766 36606 134451 36608
rect 174852 36664 177783 36666
rect 174852 36608 177722 36664
rect 177778 36608 177783 36664
rect 174852 36606 177783 36608
rect 134385 36603 134451 36606
rect 177717 36603 177783 36606
rect 100897 36528 104042 36530
rect 100897 36472 100902 36528
rect 100958 36472 104042 36528
rect 100897 36470 104042 36472
rect 185077 36530 185143 36533
rect 187886 36530 187946 36704
rect 185077 36528 187946 36530
rect 185077 36472 185082 36528
rect 185138 36472 187946 36528
rect 185077 36470 187946 36472
rect 100897 36467 100963 36470
rect 185077 36467 185143 36470
rect 142573 36394 142639 36397
rect 142573 36392 145074 36394
rect 142573 36336 142578 36392
rect 142634 36336 145074 36392
rect 142573 36334 145074 36336
rect 142573 36331 142639 36334
rect 145014 36160 145074 36334
rect 47862 35714 47922 36160
rect 58209 36122 58275 36125
rect 93997 36122 94063 36125
rect 58209 36120 60956 36122
rect 58209 36064 58214 36120
rect 58270 36064 60956 36120
rect 58209 36062 60956 36064
rect 90764 36120 94063 36122
rect 90764 36064 94002 36120
rect 94058 36064 94063 36120
rect 90764 36062 94063 36064
rect 58209 36059 58275 36062
rect 93997 36059 94063 36062
rect 92893 35986 92959 35989
rect 90734 35984 92959 35986
rect 90734 35928 92898 35984
rect 92954 35928 92959 35984
rect 90734 35926 92959 35928
rect 50021 35714 50087 35717
rect 47862 35712 50087 35714
rect 47862 35656 50026 35712
rect 50082 35656 50087 35712
rect 47862 35654 50087 35656
rect 50021 35651 50087 35654
rect 90734 35480 90794 35926
rect 92893 35923 92959 35926
rect 100989 35714 101055 35717
rect 103982 35714 104042 36160
rect 131766 35986 131826 36160
rect 177717 36122 177783 36125
rect 174852 36120 177783 36122
rect 174852 36064 177722 36120
rect 177778 36064 177783 36120
rect 174852 36062 177783 36064
rect 177717 36059 177783 36062
rect 134661 35986 134727 35989
rect 131766 35984 134727 35986
rect 131766 35928 134666 35984
rect 134722 35928 134727 35984
rect 131766 35926 134727 35928
rect 134661 35923 134727 35926
rect 142389 35986 142455 35989
rect 142389 35984 145074 35986
rect 142389 35928 142394 35984
rect 142450 35928 145074 35984
rect 142389 35926 145074 35928
rect 142389 35923 142455 35926
rect 100989 35712 104042 35714
rect 100989 35656 100994 35712
rect 101050 35656 104042 35712
rect 100989 35654 104042 35656
rect 100989 35651 101055 35654
rect 145014 35480 145074 35926
rect 185445 35714 185511 35717
rect 187886 35714 187946 36160
rect 185445 35712 187946 35714
rect 185445 35656 185450 35712
rect 185506 35656 187946 35712
rect 185445 35654 187946 35656
rect 185445 35651 185511 35654
rect 47862 35306 47922 35480
rect 58301 35442 58367 35445
rect 58301 35440 60956 35442
rect 58301 35384 58306 35440
rect 58362 35384 60956 35440
rect 58301 35382 60956 35384
rect 58301 35379 58367 35382
rect 51217 35306 51283 35309
rect 47862 35304 51283 35306
rect 47862 35248 51222 35304
rect 51278 35248 51283 35304
rect 47862 35246 51283 35248
rect 51217 35243 51283 35246
rect 100713 35170 100779 35173
rect 103982 35170 104042 35480
rect 131766 35306 131826 35480
rect 177349 35442 177415 35445
rect 174852 35440 177415 35442
rect 174852 35384 177354 35440
rect 177410 35384 177415 35440
rect 174852 35382 177415 35384
rect 177349 35379 177415 35382
rect 134109 35306 134175 35309
rect 131766 35304 134175 35306
rect 131766 35248 134114 35304
rect 134170 35248 134175 35304
rect 131766 35246 134175 35248
rect 134109 35243 134175 35246
rect 184893 35306 184959 35309
rect 187886 35306 187946 35480
rect 184893 35304 187946 35306
rect 184893 35248 184898 35304
rect 184954 35248 187946 35304
rect 184893 35246 187946 35248
rect 184893 35243 184959 35246
rect 100713 35168 104042 35170
rect 100713 35112 100718 35168
rect 100774 35112 104042 35168
rect 100713 35110 104042 35112
rect 100713 35107 100779 35110
rect 47862 34490 47922 34936
rect 58209 34898 58275 34901
rect 93997 34898 94063 34901
rect 58209 34896 60956 34898
rect 58209 34840 58214 34896
rect 58270 34840 60956 34896
rect 58209 34838 60956 34840
rect 90764 34896 94063 34898
rect 90764 34840 94002 34896
rect 94058 34840 94063 34896
rect 90764 34838 94063 34840
rect 58209 34835 58275 34838
rect 93997 34835 94063 34838
rect 93445 34626 93511 34629
rect 90734 34624 93511 34626
rect 90734 34568 93450 34624
rect 93506 34568 93511 34624
rect 90734 34566 93511 34568
rect 50205 34490 50271 34493
rect 47862 34488 50271 34490
rect 47862 34432 50210 34488
rect 50266 34432 50271 34488
rect 47862 34430 50271 34432
rect 50205 34427 50271 34430
rect 90734 34256 90794 34566
rect 93445 34563 93511 34566
rect 101081 34490 101147 34493
rect 103982 34490 104042 34936
rect 101081 34488 104042 34490
rect 101081 34432 101086 34488
rect 101142 34432 104042 34488
rect 101081 34430 104042 34432
rect 131766 34490 131826 34936
rect 142573 34898 142639 34901
rect 177717 34898 177783 34901
rect 142573 34896 145044 34898
rect 142573 34840 142578 34896
rect 142634 34840 145044 34896
rect 142573 34838 145044 34840
rect 174852 34896 177783 34898
rect 174852 34840 177722 34896
rect 177778 34840 177783 34896
rect 174852 34838 177783 34840
rect 142573 34835 142639 34838
rect 177717 34835 177783 34838
rect 142389 34762 142455 34765
rect 142389 34760 145074 34762
rect 142389 34704 142394 34760
rect 142450 34704 145074 34760
rect 142389 34702 145074 34704
rect 142389 34699 142455 34702
rect 134569 34490 134635 34493
rect 131766 34488 134635 34490
rect 131766 34432 134574 34488
rect 134630 34432 134635 34488
rect 131766 34430 134635 34432
rect 101081 34427 101147 34430
rect 134569 34427 134635 34430
rect 145014 34256 145074 34702
rect 185261 34490 185327 34493
rect 187886 34490 187946 34936
rect 185261 34488 187946 34490
rect 185261 34432 185266 34488
rect 185322 34432 187946 34488
rect 185261 34430 187946 34432
rect 185261 34427 185327 34430
rect 47862 34218 47922 34256
rect 51217 34218 51283 34221
rect 47862 34216 51283 34218
rect 47862 34160 51222 34216
rect 51278 34160 51283 34216
rect 47862 34158 51283 34160
rect 51217 34155 51283 34158
rect 58301 34218 58367 34221
rect 58301 34216 60956 34218
rect 58301 34160 58306 34216
rect 58362 34160 60956 34216
rect 58301 34158 60956 34160
rect 58301 34155 58367 34158
rect 100989 33946 101055 33949
rect 103982 33946 104042 34256
rect 131766 34218 131826 34256
rect 134661 34218 134727 34221
rect 177625 34218 177691 34221
rect 131766 34216 134727 34218
rect 131766 34160 134666 34216
rect 134722 34160 134727 34216
rect 131766 34158 134727 34160
rect 174852 34216 177691 34218
rect 174852 34160 177630 34216
rect 177686 34160 177691 34216
rect 174852 34158 177691 34160
rect 134661 34155 134727 34158
rect 177625 34155 177691 34158
rect 100989 33944 104042 33946
rect 100989 33888 100994 33944
rect 101050 33888 104042 33944
rect 100989 33886 104042 33888
rect 185169 33946 185235 33949
rect 187886 33946 187946 34256
rect 185169 33944 187946 33946
rect 185169 33888 185174 33944
rect 185230 33888 187946 33944
rect 185169 33886 187946 33888
rect 100989 33883 101055 33886
rect 185169 33883 185235 33886
rect 51217 33810 51283 33813
rect 47862 33808 51283 33810
rect 47862 33752 51222 33808
rect 51278 33752 51283 33808
rect 47862 33750 51283 33752
rect 47862 33712 47922 33750
rect 51217 33747 51283 33750
rect 100805 33810 100871 33813
rect 134661 33810 134727 33813
rect 100805 33808 104042 33810
rect 100805 33752 100810 33808
rect 100866 33752 104042 33808
rect 100805 33750 104042 33752
rect 100805 33747 100871 33750
rect 103982 33716 104042 33750
rect 131766 33808 134727 33810
rect 131766 33752 134666 33808
rect 134722 33752 134727 33808
rect 131766 33750 134727 33752
rect 131766 33712 131826 33750
rect 134661 33747 134727 33750
rect 184985 33810 185051 33813
rect 184985 33808 187946 33810
rect 184985 33752 184990 33808
rect 185046 33752 187946 33808
rect 184985 33750 187946 33752
rect 184985 33747 185051 33750
rect 187886 33712 187946 33750
rect 58209 33674 58275 33677
rect 93905 33674 93971 33677
rect 58209 33672 60956 33674
rect 58209 33616 58214 33672
rect 58270 33616 60956 33672
rect 58209 33614 60956 33616
rect 90764 33672 93971 33674
rect 90764 33616 93910 33672
rect 93966 33616 93971 33672
rect 90764 33614 93971 33616
rect 58209 33611 58275 33614
rect 93905 33611 93971 33614
rect 142481 33674 142547 33677
rect 177625 33674 177691 33677
rect 142481 33672 145044 33674
rect 142481 33616 142486 33672
rect 142542 33616 145044 33672
rect 142481 33614 145044 33616
rect 174852 33672 177691 33674
rect 174852 33616 177630 33672
rect 177686 33616 177691 33672
rect 174852 33614 177691 33616
rect 142481 33611 142547 33614
rect 177625 33611 177691 33614
rect 93997 33402 94063 33405
rect 90734 33400 94063 33402
rect 90734 33344 94002 33400
rect 94058 33344 94063 33400
rect 90734 33342 94063 33344
rect 90734 33168 90794 33342
rect 93997 33339 94063 33342
rect 142389 33402 142455 33405
rect 215713 33402 215779 33405
rect 142389 33400 145074 33402
rect 142389 33344 142394 33400
rect 142450 33344 145074 33400
rect 142389 33342 145074 33344
rect 142389 33339 142455 33342
rect 145014 33168 145074 33342
rect 215670 33400 215779 33402
rect 215670 33344 215718 33400
rect 215774 33344 215779 33400
rect 215670 33339 215779 33344
rect 47862 32722 47922 33168
rect 58209 33130 58275 33133
rect 58209 33128 60956 33130
rect 58209 33072 58214 33128
rect 58270 33072 60956 33128
rect 58209 33070 60956 33072
rect 58209 33067 58275 33070
rect 93813 32994 93879 32997
rect 90734 32992 93879 32994
rect 90734 32936 93818 32992
rect 93874 32936 93879 32992
rect 90734 32934 93879 32936
rect 50021 32722 50087 32725
rect 47862 32720 50087 32722
rect 47862 32664 50026 32720
rect 50082 32664 50087 32720
rect 47862 32662 50087 32664
rect 50021 32659 50087 32662
rect 90734 32488 90794 32934
rect 93813 32931 93879 32934
rect 100989 32722 101055 32725
rect 103982 32722 104042 33168
rect 100989 32720 104042 32722
rect 100989 32664 100994 32720
rect 101050 32664 104042 32720
rect 100989 32662 104042 32664
rect 131766 32722 131826 33168
rect 177717 33130 177783 33133
rect 174852 33128 177783 33130
rect 174852 33072 177722 33128
rect 177778 33072 177783 33128
rect 174852 33070 177783 33072
rect 177717 33067 177783 33070
rect 142389 32994 142455 32997
rect 142389 32992 145074 32994
rect 142389 32936 142394 32992
rect 142450 32936 145074 32992
rect 142389 32934 145074 32936
rect 142389 32931 142455 32934
rect 134293 32722 134359 32725
rect 131766 32720 134359 32722
rect 131766 32664 134298 32720
rect 134354 32664 134359 32720
rect 131766 32662 134359 32664
rect 100989 32659 101055 32662
rect 134293 32659 134359 32662
rect 145014 32488 145074 32934
rect 185169 32722 185235 32725
rect 187886 32722 187946 33168
rect 215670 32896 215730 33339
rect 185169 32720 187946 32722
rect 185169 32664 185174 32720
rect 185230 32664 187946 32720
rect 185169 32662 187946 32664
rect 185169 32659 185235 32662
rect 47862 32450 47922 32488
rect 51217 32450 51283 32453
rect 47862 32448 51283 32450
rect 47862 32392 51222 32448
rect 51278 32392 51283 32448
rect 47862 32390 51283 32392
rect 51217 32387 51283 32390
rect 58209 32450 58275 32453
rect 58209 32448 60956 32450
rect 58209 32392 58214 32448
rect 58270 32392 60956 32448
rect 58209 32390 60956 32392
rect 58209 32387 58275 32390
rect 100897 32314 100963 32317
rect 103982 32314 104042 32488
rect 131766 32450 131826 32488
rect 134385 32450 134451 32453
rect 177809 32450 177875 32453
rect 131766 32448 134451 32450
rect 131766 32392 134390 32448
rect 134446 32392 134451 32448
rect 131766 32390 134451 32392
rect 174852 32448 177875 32450
rect 174852 32392 177814 32448
rect 177870 32392 177875 32448
rect 174852 32390 177875 32392
rect 134385 32387 134451 32390
rect 177809 32387 177875 32390
rect 100897 32312 104042 32314
rect 100897 32256 100902 32312
rect 100958 32256 104042 32312
rect 100897 32254 104042 32256
rect 185077 32314 185143 32317
rect 187886 32314 187946 32488
rect 185077 32312 187946 32314
rect 185077 32256 185082 32312
rect 185138 32256 187946 32312
rect 185077 32254 187946 32256
rect 100897 32251 100963 32254
rect 185077 32251 185143 32254
rect 142481 32178 142547 32181
rect 142481 32176 145074 32178
rect 142481 32120 142486 32176
rect 142542 32120 145074 32176
rect 142481 32118 145074 32120
rect 142481 32115 142547 32118
rect 145014 31944 145074 32118
rect 47862 31634 47922 31944
rect 58209 31906 58275 31909
rect 93997 31906 94063 31909
rect 58209 31904 60956 31906
rect 58209 31848 58214 31904
rect 58270 31848 60956 31904
rect 58209 31846 60956 31848
rect 90764 31904 94063 31906
rect 90764 31848 94002 31904
rect 94058 31848 94063 31904
rect 90764 31846 94063 31848
rect 58209 31843 58275 31846
rect 93997 31843 94063 31846
rect 93905 31770 93971 31773
rect 90734 31768 93971 31770
rect 90734 31712 93910 31768
rect 93966 31712 93971 31768
rect 90734 31710 93971 31712
rect 51125 31634 51191 31637
rect 47862 31632 51191 31634
rect 47862 31576 51130 31632
rect 51186 31576 51191 31632
rect 47862 31574 51191 31576
rect 51125 31571 51191 31574
rect 47862 31226 47922 31400
rect 90734 31264 90794 31710
rect 93905 31707 93971 31710
rect 100989 31498 101055 31501
rect 103982 31498 104042 31944
rect 131766 31634 131826 31944
rect 176981 31906 177047 31909
rect 174852 31904 177047 31906
rect 174852 31848 176986 31904
rect 177042 31848 177047 31904
rect 174852 31846 177047 31848
rect 176981 31843 177047 31846
rect 142389 31770 142455 31773
rect 142389 31768 145074 31770
rect 142389 31712 142394 31768
rect 142450 31712 145074 31768
rect 142389 31710 145074 31712
rect 142389 31707 142455 31710
rect 134661 31634 134727 31637
rect 131766 31632 134727 31634
rect 131766 31576 134666 31632
rect 134722 31576 134727 31632
rect 131766 31574 134727 31576
rect 134661 31571 134727 31574
rect 100989 31496 104042 31498
rect 100989 31440 100994 31496
rect 101050 31440 104042 31496
rect 100989 31438 104042 31440
rect 100989 31435 101055 31438
rect 145014 31264 145074 31710
rect 185169 31498 185235 31501
rect 187886 31498 187946 31944
rect 185169 31496 187946 31498
rect 185169 31440 185174 31496
rect 185230 31440 187946 31496
rect 185169 31438 187946 31440
rect 185169 31435 185235 31438
rect 51217 31226 51283 31229
rect 47862 31224 51283 31226
rect 47862 31168 51222 31224
rect 51278 31168 51283 31224
rect 47862 31166 51283 31168
rect 51217 31163 51283 31166
rect 58301 31226 58367 31229
rect 58301 31224 60956 31226
rect 58301 31168 58306 31224
rect 58362 31168 60956 31224
rect 58301 31166 60956 31168
rect 58301 31163 58367 31166
rect 100805 30954 100871 30957
rect 103982 30954 104042 31264
rect 131766 31090 131826 31264
rect 177717 31226 177783 31229
rect 174852 31224 177783 31226
rect 174852 31168 177722 31224
rect 177778 31168 177783 31224
rect 174852 31166 177783 31168
rect 177717 31163 177783 31166
rect 134661 31090 134727 31093
rect 131766 31088 134727 31090
rect 131766 31032 134666 31088
rect 134722 31032 134727 31088
rect 131766 31030 134727 31032
rect 134661 31027 134727 31030
rect 100805 30952 104042 30954
rect 100805 30896 100810 30952
rect 100866 30896 104042 30952
rect 100805 30894 104042 30896
rect 184985 30954 185051 30957
rect 187886 30954 187946 31264
rect 184985 30952 187946 30954
rect 184985 30896 184990 30952
rect 185046 30896 187946 30952
rect 184985 30894 187946 30896
rect 100805 30891 100871 30894
rect 184985 30891 185051 30894
rect 47862 30410 47922 30720
rect 58209 30682 58275 30685
rect 93997 30682 94063 30685
rect 58209 30680 60956 30682
rect 58209 30624 58214 30680
rect 58270 30624 60956 30680
rect 58209 30622 60956 30624
rect 90764 30680 94063 30682
rect 90764 30624 94002 30680
rect 94058 30624 94063 30680
rect 90764 30622 94063 30624
rect 58209 30619 58275 30622
rect 93997 30619 94063 30622
rect 92709 30546 92775 30549
rect 90734 30544 92775 30546
rect 90734 30488 92714 30544
rect 92770 30488 92775 30544
rect 90734 30486 92775 30488
rect 51125 30410 51191 30413
rect 47862 30408 51191 30410
rect 47862 30352 51130 30408
rect 51186 30352 51191 30408
rect 47862 30350 51191 30352
rect 51125 30347 51191 30350
rect 90734 30176 90794 30486
rect 92709 30483 92775 30486
rect 101081 30274 101147 30277
rect 103982 30274 104042 30720
rect 101081 30272 104042 30274
rect 101081 30216 101086 30272
rect 101142 30216 104042 30272
rect 101081 30214 104042 30216
rect 131766 30274 131826 30720
rect 142389 30682 142455 30685
rect 177441 30682 177507 30685
rect 142389 30680 145044 30682
rect 142389 30624 142394 30680
rect 142450 30624 145044 30680
rect 142389 30622 145044 30624
rect 174852 30680 177507 30682
rect 174852 30624 177446 30680
rect 177502 30624 177507 30680
rect 174852 30622 177507 30624
rect 142389 30619 142455 30622
rect 177441 30619 177507 30622
rect 142389 30546 142455 30549
rect 142389 30544 145074 30546
rect 142389 30488 142394 30544
rect 142450 30488 145074 30544
rect 142389 30486 145074 30488
rect 142389 30483 142455 30486
rect 134753 30274 134819 30277
rect 131766 30272 134819 30274
rect 131766 30216 134758 30272
rect 134814 30216 134819 30272
rect 131766 30214 134819 30216
rect 101081 30211 101147 30214
rect 134753 30211 134819 30214
rect 145014 30176 145074 30486
rect 185261 30274 185327 30277
rect 187886 30274 187946 30720
rect 185261 30272 187946 30274
rect 185261 30216 185266 30272
rect 185322 30216 187946 30272
rect 185261 30214 187946 30216
rect 185261 30211 185327 30214
rect 47862 29866 47922 30176
rect 58301 30138 58367 30141
rect 177165 30138 177231 30141
rect 58301 30136 60956 30138
rect 58301 30080 58306 30136
rect 58362 30080 60956 30136
rect 58301 30078 60956 30080
rect 174852 30136 177231 30138
rect 174852 30080 177170 30136
rect 177226 30080 177231 30136
rect 174852 30078 177231 30080
rect 58301 30075 58367 30078
rect 177165 30075 177231 30078
rect 51217 29866 51283 29869
rect 47862 29864 51283 29866
rect 47862 29808 51222 29864
rect 51278 29808 51283 29864
rect 47862 29806 51283 29808
rect 51217 29803 51283 29806
rect 100989 29730 101055 29733
rect 103982 29730 104042 30040
rect 131766 29866 131826 30040
rect 134201 29866 134267 29869
rect 131766 29864 134267 29866
rect 131766 29808 134206 29864
rect 134262 29808 134267 29864
rect 131766 29806 134267 29808
rect 134201 29803 134267 29806
rect 100989 29728 104042 29730
rect 100989 29672 100994 29728
rect 101050 29672 104042 29728
rect 100989 29670 104042 29672
rect 185169 29730 185235 29733
rect 187886 29730 187946 30040
rect 185169 29728 187946 29730
rect 185169 29672 185174 29728
rect 185230 29672 187946 29728
rect 185169 29670 187946 29672
rect 100989 29667 101055 29670
rect 185169 29667 185235 29670
rect 47862 29186 47922 29496
rect 58209 29458 58275 29461
rect 93997 29458 94063 29461
rect 58209 29456 60956 29458
rect 58209 29400 58214 29456
rect 58270 29400 60956 29456
rect 58209 29398 60956 29400
rect 90764 29456 94063 29458
rect 90764 29400 94002 29456
rect 94058 29400 94063 29456
rect 90764 29398 94063 29400
rect 58209 29395 58275 29398
rect 93997 29395 94063 29398
rect 51125 29186 51191 29189
rect 93905 29186 93971 29189
rect 47862 29184 51191 29186
rect 47862 29128 51130 29184
rect 51186 29128 51191 29184
rect 47862 29126 51191 29128
rect 51125 29123 51191 29126
rect 90734 29184 93971 29186
rect 90734 29128 93910 29184
rect 93966 29128 93971 29184
rect 90734 29126 93971 29128
rect 90734 28952 90794 29126
rect 93905 29123 93971 29126
rect 101173 29050 101239 29053
rect 103982 29050 104042 29496
rect 101173 29048 104042 29050
rect 101173 28992 101178 29048
rect 101234 28992 104042 29048
rect 101173 28990 104042 28992
rect 131766 29050 131826 29496
rect 143585 29458 143651 29461
rect 177717 29458 177783 29461
rect 143585 29456 145044 29458
rect 143585 29400 143590 29456
rect 143646 29400 145044 29456
rect 143585 29398 145044 29400
rect 174852 29456 177783 29458
rect 174852 29400 177722 29456
rect 177778 29400 177783 29456
rect 174852 29398 177783 29400
rect 143585 29395 143651 29398
rect 177717 29395 177783 29398
rect 142389 29322 142455 29325
rect 142389 29320 145074 29322
rect 142389 29264 142394 29320
rect 142450 29264 145074 29320
rect 142389 29262 145074 29264
rect 142389 29259 142455 29262
rect 134569 29050 134635 29053
rect 131766 29048 134635 29050
rect 131766 28992 134574 29048
rect 134630 28992 134635 29048
rect 131766 28990 134635 28992
rect 101173 28987 101239 28990
rect 134569 28987 134635 28990
rect 145014 28952 145074 29262
rect 185353 29050 185419 29053
rect 187886 29050 187946 29496
rect 185353 29048 187946 29050
rect 185353 28992 185358 29048
rect 185414 28992 187946 29048
rect 185353 28990 187946 28992
rect 185353 28987 185419 28990
rect 47862 28778 47922 28952
rect 58209 28914 58275 28917
rect 177809 28914 177875 28917
rect 58209 28912 60956 28914
rect 58209 28856 58214 28912
rect 58270 28856 60956 28912
rect 58209 28854 60956 28856
rect 174852 28912 177875 28914
rect 174852 28856 177814 28912
rect 177870 28856 177875 28912
rect 174852 28854 177875 28856
rect 58209 28851 58275 28854
rect 177809 28851 177875 28854
rect 51217 28778 51283 28781
rect 92709 28778 92775 28781
rect 47862 28776 51283 28778
rect 47862 28720 51222 28776
rect 51278 28720 51283 28776
rect 47862 28718 51283 28720
rect 51217 28715 51283 28718
rect 90734 28776 92775 28778
rect 90734 28720 92714 28776
rect 92770 28720 92775 28776
rect 90734 28718 92775 28720
rect 47862 28370 47922 28408
rect 51217 28370 51283 28373
rect 47862 28368 51283 28370
rect 47862 28312 51222 28368
rect 51278 28312 51283 28368
rect 47862 28310 51283 28312
rect 51217 28307 51283 28310
rect 90734 28272 90794 28718
rect 92709 28715 92775 28718
rect 101081 28506 101147 28509
rect 103982 28506 104042 28816
rect 131766 28642 131826 28816
rect 142481 28778 142547 28781
rect 142481 28776 145074 28778
rect 142481 28720 142486 28776
rect 142542 28720 145074 28776
rect 142481 28718 145074 28720
rect 142481 28715 142547 28718
rect 134753 28642 134819 28645
rect 131766 28640 134819 28642
rect 131766 28584 134758 28640
rect 134814 28584 134819 28640
rect 131766 28582 134819 28584
rect 134753 28579 134819 28582
rect 101081 28504 104042 28506
rect 101081 28448 101086 28504
rect 101142 28448 104042 28504
rect 101081 28446 104042 28448
rect 101081 28443 101147 28446
rect 145014 28272 145074 28718
rect 185261 28506 185327 28509
rect 187886 28506 187946 28816
rect 185261 28504 187946 28506
rect 185261 28448 185266 28504
rect 185322 28448 187946 28504
rect 185261 28446 187946 28448
rect 185261 28443 185327 28446
rect 58209 28234 58275 28237
rect 100989 28234 101055 28237
rect 103982 28234 104042 28272
rect 58209 28232 60956 28234
rect 58209 28176 58214 28232
rect 58270 28176 60956 28232
rect 58209 28174 60956 28176
rect 100989 28232 104042 28234
rect 100989 28176 100994 28232
rect 101050 28176 104042 28232
rect 100989 28174 104042 28176
rect 131766 28234 131826 28272
rect 134753 28234 134819 28237
rect 177625 28234 177691 28237
rect 131766 28232 134819 28234
rect 131766 28176 134758 28232
rect 134814 28176 134819 28232
rect 131766 28174 134819 28176
rect 174852 28232 177691 28234
rect 174852 28176 177630 28232
rect 177686 28176 177691 28232
rect 174852 28174 177691 28176
rect 58209 28171 58275 28174
rect 100989 28171 101055 28174
rect 134753 28171 134819 28174
rect 177625 28171 177691 28174
rect 185169 28234 185235 28237
rect 187886 28234 187946 28272
rect 185169 28232 187946 28234
rect 185169 28176 185174 28232
rect 185230 28176 187946 28232
rect 185169 28174 187946 28176
rect 185169 28171 185235 28174
rect 93997 27962 94063 27965
rect 90734 27960 94063 27962
rect 90734 27904 94002 27960
rect 94058 27904 94063 27960
rect 90734 27902 94063 27904
rect 90734 27728 90794 27902
rect 93997 27899 94063 27902
rect 142389 27962 142455 27965
rect 142389 27960 145074 27962
rect 142389 27904 142394 27960
rect 142450 27904 145074 27960
rect 142389 27902 145074 27904
rect 142389 27899 142455 27902
rect 145014 27728 145074 27902
rect 47862 27418 47922 27728
rect 58209 27690 58275 27693
rect 177717 27690 177783 27693
rect 58209 27688 60956 27690
rect 58209 27632 58214 27688
rect 58270 27632 60956 27688
rect 58209 27630 60956 27632
rect 174852 27688 177783 27690
rect 174852 27632 177722 27688
rect 177778 27632 177783 27688
rect 174852 27630 177783 27632
rect 58209 27627 58275 27630
rect 177717 27627 177783 27630
rect 92709 27554 92775 27557
rect 90734 27552 92775 27554
rect 90734 27496 92714 27552
rect 92770 27496 92775 27552
rect 90734 27494 92775 27496
rect 51125 27418 51191 27421
rect 47862 27416 51191 27418
rect 47862 27360 51130 27416
rect 51186 27360 51191 27416
rect 47862 27358 51191 27360
rect 51125 27355 51191 27358
rect 90734 27184 90794 27494
rect 92709 27491 92775 27494
rect 100989 27282 101055 27285
rect 103982 27282 104042 27592
rect 100989 27280 104042 27282
rect 100989 27224 100994 27280
rect 101050 27224 104042 27280
rect 100989 27222 104042 27224
rect 131766 27282 131826 27592
rect 142389 27554 142455 27557
rect 142389 27552 145074 27554
rect 142389 27496 142394 27552
rect 142450 27496 145074 27552
rect 142389 27494 145074 27496
rect 142389 27491 142455 27494
rect 134569 27282 134635 27285
rect 131766 27280 134635 27282
rect 131766 27224 134574 27280
rect 134630 27224 134635 27280
rect 131766 27222 134635 27224
rect 100989 27219 101055 27222
rect 134569 27219 134635 27222
rect 145014 27184 145074 27494
rect 185169 27282 185235 27285
rect 187886 27282 187946 27592
rect 185169 27280 187946 27282
rect 185169 27224 185174 27280
rect 185230 27224 187946 27280
rect 185169 27222 187946 27224
rect 185169 27219 185235 27222
rect 47862 27010 47922 27184
rect 58301 27146 58367 27149
rect 177257 27146 177323 27149
rect 58301 27144 60956 27146
rect 58301 27088 58306 27144
rect 58362 27088 60956 27144
rect 58301 27086 60956 27088
rect 174852 27144 177323 27146
rect 174852 27088 177262 27144
rect 177318 27088 177323 27144
rect 174852 27086 177323 27088
rect 58301 27083 58367 27086
rect 177257 27083 177323 27086
rect 51217 27010 51283 27013
rect 47862 27008 51283 27010
rect 47862 26952 51222 27008
rect 51278 26952 51283 27008
rect 47862 26950 51283 26952
rect 51217 26947 51283 26950
rect 101173 26874 101239 26877
rect 103982 26874 104042 27048
rect 131766 27010 131826 27048
rect 134753 27010 134819 27013
rect 131766 27008 134819 27010
rect 131766 26952 134758 27008
rect 134814 26952 134819 27008
rect 131766 26950 134819 26952
rect 134753 26947 134819 26950
rect 101173 26872 104042 26874
rect 101173 26816 101178 26872
rect 101234 26816 104042 26872
rect 101173 26814 104042 26816
rect 185353 26874 185419 26877
rect 187886 26874 187946 27048
rect 185353 26872 187946 26874
rect 185353 26816 185358 26872
rect 185414 26816 187946 26872
rect 185353 26814 187946 26816
rect 101173 26811 101239 26814
rect 185353 26811 185419 26814
rect 93905 26738 93971 26741
rect 90734 26736 93971 26738
rect 90734 26680 93910 26736
rect 93966 26680 93971 26736
rect 90734 26678 93971 26680
rect 90734 26504 90794 26678
rect 93905 26675 93971 26678
rect 142481 26738 142547 26741
rect 142481 26736 145074 26738
rect 142481 26680 142486 26736
rect 142542 26680 145074 26736
rect 142481 26678 145074 26680
rect 142481 26675 142547 26678
rect 145014 26504 145074 26678
rect 47862 26194 47922 26504
rect 58209 26466 58275 26469
rect 177441 26466 177507 26469
rect 58209 26464 60956 26466
rect 58209 26408 58214 26464
rect 58270 26408 60956 26464
rect 58209 26406 60956 26408
rect 174852 26464 177507 26466
rect 174852 26408 177446 26464
rect 177502 26408 177507 26464
rect 174852 26406 177507 26408
rect 58209 26403 58275 26406
rect 177441 26403 177507 26406
rect 93997 26330 94063 26333
rect 90734 26328 94063 26330
rect 90734 26272 94002 26328
rect 94058 26272 94063 26328
rect 90734 26270 94063 26272
rect 50481 26194 50547 26197
rect 47862 26192 50547 26194
rect 47862 26136 50486 26192
rect 50542 26136 50547 26192
rect 47862 26134 50547 26136
rect 50481 26131 50547 26134
rect 90734 25960 90794 26270
rect 93997 26267 94063 26270
rect 101081 26058 101147 26061
rect 103982 26058 104042 26368
rect 101081 26056 104042 26058
rect 101081 26000 101086 26056
rect 101142 26000 104042 26056
rect 101081 25998 104042 26000
rect 131766 26058 131826 26368
rect 142389 26330 142455 26333
rect 142389 26328 145074 26330
rect 142389 26272 142394 26328
rect 142450 26272 145074 26328
rect 142389 26270 145074 26272
rect 142389 26267 142455 26270
rect 134569 26058 134635 26061
rect 131766 26056 134635 26058
rect 131766 26000 134574 26056
rect 134630 26000 134635 26056
rect 131766 25998 134635 26000
rect 101081 25995 101147 25998
rect 134569 25995 134635 25998
rect 145014 25960 145074 26270
rect 185537 26058 185603 26061
rect 187886 26058 187946 26368
rect 185537 26056 187946 26058
rect 185537 26000 185542 26056
rect 185598 26000 187946 26056
rect 185537 25998 187946 26000
rect 185537 25995 185603 25998
rect 47862 25786 47922 25960
rect 58301 25922 58367 25925
rect 177717 25922 177783 25925
rect 58301 25920 60956 25922
rect 58301 25864 58306 25920
rect 58362 25864 60956 25920
rect 58301 25862 60956 25864
rect 174852 25920 177783 25922
rect 174852 25864 177722 25920
rect 177778 25864 177783 25920
rect 174852 25862 177783 25864
rect 58301 25859 58367 25862
rect 177717 25859 177783 25862
rect 51217 25786 51283 25789
rect 47862 25784 51283 25786
rect 47862 25728 51222 25784
rect 51278 25728 51283 25784
rect 47862 25726 51283 25728
rect 51217 25723 51283 25726
rect 100989 25650 101055 25653
rect 103982 25650 104042 25824
rect 100989 25648 104042 25650
rect 100989 25592 100994 25648
rect 101050 25592 104042 25648
rect 100989 25590 104042 25592
rect 131766 25650 131826 25824
rect 134753 25650 134819 25653
rect 131766 25648 134819 25650
rect 131766 25592 134758 25648
rect 134814 25592 134819 25648
rect 131766 25590 134819 25592
rect 100989 25587 101055 25590
rect 134753 25587 134819 25590
rect 185445 25650 185511 25653
rect 187886 25650 187946 25824
rect 185445 25648 187946 25650
rect 185445 25592 185450 25648
rect 185506 25592 187946 25648
rect 185445 25590 187946 25592
rect 185445 25587 185511 25590
rect 18097 25514 18163 25517
rect 19894 25514 19954 25552
rect 51125 25514 51191 25517
rect 18097 25512 19954 25514
rect 18097 25456 18102 25512
rect 18158 25456 19954 25512
rect 18097 25454 19954 25456
rect 47862 25512 51191 25514
rect 47862 25456 51130 25512
rect 51186 25456 51191 25512
rect 47862 25454 51191 25456
rect 18097 25451 18163 25454
rect 47862 25416 47922 25454
rect 51125 25451 51191 25454
rect 59497 25242 59563 25245
rect 93997 25242 94063 25245
rect 59497 25240 60956 25242
rect 59497 25184 59502 25240
rect 59558 25184 60956 25240
rect 59497 25182 60956 25184
rect 90764 25240 94063 25242
rect 90764 25184 94002 25240
rect 94058 25184 94063 25240
rect 90764 25182 94063 25184
rect 59497 25179 59563 25182
rect 93997 25179 94063 25182
rect 142573 25242 142639 25245
rect 177717 25242 177783 25245
rect 142573 25240 145044 25242
rect 142573 25184 142578 25240
rect 142634 25184 145044 25240
rect 142573 25182 145044 25184
rect 174852 25240 177783 25242
rect 174852 25184 177722 25240
rect 177778 25184 177783 25240
rect 174852 25182 177783 25184
rect 142573 25179 142639 25182
rect 177717 25179 177783 25182
rect 93905 24970 93971 24973
rect 90734 24968 93971 24970
rect 90734 24912 93910 24968
rect 93966 24912 93971 24968
rect 90734 24910 93971 24912
rect 90734 24736 90794 24910
rect 93905 24907 93971 24910
rect 101081 24834 101147 24837
rect 103982 24834 104042 25144
rect 101081 24832 104042 24834
rect 101081 24776 101086 24832
rect 101142 24776 104042 24832
rect 101081 24774 104042 24776
rect 131766 24834 131826 25144
rect 142389 25106 142455 25109
rect 142389 25104 145074 25106
rect 142389 25048 142394 25104
rect 142450 25048 145074 25104
rect 142389 25046 145074 25048
rect 142389 25043 142455 25046
rect 134569 24834 134635 24837
rect 131766 24832 134635 24834
rect 131766 24776 134574 24832
rect 134630 24776 134635 24832
rect 131766 24774 134635 24776
rect 101081 24771 101147 24774
rect 134569 24771 134635 24774
rect 145014 24736 145074 25046
rect 185261 24834 185327 24837
rect 187886 24834 187946 25144
rect 185261 24832 187946 24834
rect 185261 24776 185266 24832
rect 185322 24776 187946 24832
rect 185261 24774 187946 24776
rect 185261 24771 185327 24774
rect 47862 24426 47922 24736
rect 59405 24698 59471 24701
rect 177625 24698 177691 24701
rect 59405 24696 60956 24698
rect 59405 24640 59410 24696
rect 59466 24640 60956 24696
rect 59405 24638 60956 24640
rect 174852 24696 177691 24698
rect 174852 24640 177630 24696
rect 177686 24640 177691 24696
rect 174852 24638 177691 24640
rect 59405 24635 59471 24638
rect 177625 24635 177691 24638
rect 93813 24562 93879 24565
rect 90734 24560 93879 24562
rect 90734 24504 93818 24560
rect 93874 24504 93879 24560
rect 90734 24502 93879 24504
rect 51125 24426 51191 24429
rect 47862 24424 51191 24426
rect 47862 24368 51130 24424
rect 51186 24368 51191 24424
rect 47862 24366 51191 24368
rect 51125 24363 51191 24366
rect 90734 24192 90794 24502
rect 93813 24499 93879 24502
rect 47862 24154 47922 24192
rect 51217 24154 51283 24157
rect 47862 24152 51283 24154
rect 47862 24096 51222 24152
rect 51278 24096 51283 24152
rect 47862 24094 51283 24096
rect 51217 24091 51283 24094
rect 59313 24154 59379 24157
rect 100989 24154 101055 24157
rect 103982 24154 104042 24600
rect 131766 24290 131826 24600
rect 142481 24562 142547 24565
rect 142481 24560 145074 24562
rect 142481 24504 142486 24560
rect 142542 24504 145074 24560
rect 142481 24502 145074 24504
rect 142481 24499 142547 24502
rect 134753 24290 134819 24293
rect 131766 24288 134819 24290
rect 131766 24232 134758 24288
rect 134814 24232 134819 24288
rect 131766 24230 134819 24232
rect 134753 24227 134819 24230
rect 145014 24192 145074 24502
rect 177349 24154 177415 24157
rect 59313 24152 60956 24154
rect 59313 24096 59318 24152
rect 59374 24096 60956 24152
rect 59313 24094 60956 24096
rect 100989 24152 104042 24154
rect 100989 24096 100994 24152
rect 101050 24096 104042 24152
rect 100989 24094 104042 24096
rect 174852 24152 177415 24154
rect 174852 24096 177354 24152
rect 177410 24096 177415 24152
rect 174852 24094 177415 24096
rect 59313 24091 59379 24094
rect 100989 24091 101055 24094
rect 177349 24091 177415 24094
rect 185169 24154 185235 24157
rect 187886 24154 187946 24600
rect 185169 24152 187946 24154
rect 185169 24096 185174 24152
rect 185230 24096 187946 24152
rect 185169 24094 187946 24096
rect 185169 24091 185235 24094
rect 93997 23746 94063 23749
rect 90734 23744 94063 23746
rect 90734 23688 94002 23744
rect 94058 23688 94063 23744
rect 90734 23686 94063 23688
rect 47862 23202 47922 23648
rect 90734 23512 90794 23686
rect 93997 23683 94063 23686
rect 100989 23610 101055 23613
rect 103982 23610 104042 23920
rect 100989 23608 104042 23610
rect 100989 23552 100994 23608
rect 101050 23552 104042 23608
rect 100989 23550 104042 23552
rect 131766 23610 131826 23920
rect 142389 23882 142455 23885
rect 142389 23880 145074 23882
rect 142389 23824 142394 23880
rect 142450 23824 145074 23880
rect 142389 23822 145074 23824
rect 142389 23819 142455 23822
rect 134569 23610 134635 23613
rect 131766 23608 134635 23610
rect 131766 23552 134574 23608
rect 134630 23552 134635 23608
rect 131766 23550 134635 23552
rect 100989 23547 101055 23550
rect 134569 23547 134635 23550
rect 145014 23512 145074 23822
rect 185261 23610 185327 23613
rect 187886 23610 187946 23920
rect 185261 23608 187946 23610
rect 185261 23552 185266 23608
rect 185322 23552 187946 23608
rect 185261 23550 187946 23552
rect 185261 23547 185327 23550
rect 58209 23474 58275 23477
rect 177717 23474 177783 23477
rect 58209 23472 60956 23474
rect 58209 23416 58214 23472
rect 58270 23416 60956 23472
rect 58209 23414 60956 23416
rect 174852 23472 177783 23474
rect 174852 23416 177722 23472
rect 177778 23416 177783 23472
rect 174852 23414 177783 23416
rect 58209 23411 58275 23414
rect 177717 23411 177783 23414
rect 92893 23338 92959 23341
rect 90734 23336 92959 23338
rect 90734 23280 92898 23336
rect 92954 23280 92959 23336
rect 90734 23278 92959 23280
rect 50205 23202 50271 23205
rect 47862 23200 50271 23202
rect 47862 23144 50210 23200
rect 50266 23144 50271 23200
rect 47862 23142 50271 23144
rect 50205 23139 50271 23142
rect 90734 22968 90794 23278
rect 92893 23275 92959 23278
rect 47862 22930 47922 22968
rect 51217 22930 51283 22933
rect 47862 22928 51283 22930
rect 47862 22872 51222 22928
rect 51278 22872 51283 22928
rect 47862 22870 51283 22872
rect 51217 22867 51283 22870
rect 58301 22930 58367 22933
rect 101081 22930 101147 22933
rect 103982 22930 104042 23376
rect 131766 23202 131826 23376
rect 142481 23338 142547 23341
rect 142481 23336 145074 23338
rect 142481 23280 142486 23336
rect 142542 23280 145074 23336
rect 142481 23278 145074 23280
rect 142481 23275 142547 23278
rect 134753 23202 134819 23205
rect 131766 23200 134819 23202
rect 131766 23144 134758 23200
rect 134814 23144 134819 23200
rect 131766 23142 134819 23144
rect 134753 23139 134819 23142
rect 145014 22968 145074 23278
rect 177533 22930 177599 22933
rect 58301 22928 60956 22930
rect 58301 22872 58306 22928
rect 58362 22872 60956 22928
rect 58301 22870 60956 22872
rect 101081 22928 104042 22930
rect 101081 22872 101086 22928
rect 101142 22872 104042 22928
rect 101081 22870 104042 22872
rect 174852 22928 177599 22930
rect 174852 22872 177538 22928
rect 177594 22872 177599 22928
rect 174852 22870 177599 22872
rect 58301 22867 58367 22870
rect 101081 22867 101147 22870
rect 177533 22867 177599 22870
rect 185169 22930 185235 22933
rect 187886 22930 187946 23376
rect 185169 22928 187946 22930
rect 185169 22872 185174 22928
rect 185230 22872 187946 22928
rect 185169 22870 187946 22872
rect 185169 22867 185235 22870
rect 134753 22794 134819 22797
rect 131766 22792 134819 22794
rect 131766 22736 134758 22792
rect 134814 22736 134819 22792
rect 131766 22734 134819 22736
rect 131766 22696 131826 22734
rect 134753 22731 134819 22734
rect 101173 22658 101239 22661
rect 103982 22658 104042 22696
rect 101173 22656 104042 22658
rect 101173 22600 101178 22656
rect 101234 22600 104042 22656
rect 101173 22598 104042 22600
rect 185261 22658 185327 22661
rect 187886 22658 187946 22696
rect 185261 22656 187946 22658
rect 185261 22600 185266 22656
rect 185322 22600 187946 22656
rect 185261 22598 187946 22600
rect 101173 22595 101239 22598
rect 185261 22595 185327 22598
rect 93997 22522 94063 22525
rect 135305 22522 135371 22525
rect 90734 22520 94063 22522
rect 90734 22464 94002 22520
rect 94058 22464 94063 22520
rect 90734 22462 94063 22464
rect 47862 21978 47922 22424
rect 90734 22288 90794 22462
rect 93997 22459 94063 22462
rect 131766 22520 135371 22522
rect 131766 22464 135310 22520
rect 135366 22464 135371 22520
rect 131766 22462 135371 22464
rect 100989 22386 101055 22389
rect 100989 22384 104042 22386
rect 100989 22328 100994 22384
rect 101050 22328 104042 22384
rect 100989 22326 104042 22328
rect 100989 22323 101055 22326
rect 58209 22250 58275 22253
rect 58209 22248 60956 22250
rect 58209 22192 58214 22248
rect 58270 22192 60956 22248
rect 58209 22190 60956 22192
rect 58209 22187 58275 22190
rect 103982 22156 104042 22326
rect 131766 22152 131826 22462
rect 135305 22459 135371 22462
rect 142389 22522 142455 22525
rect 142389 22520 145074 22522
rect 142389 22464 142394 22520
rect 142450 22464 145074 22520
rect 142389 22462 145074 22464
rect 142389 22459 142455 22462
rect 145014 22288 145074 22462
rect 185169 22386 185235 22389
rect 185169 22384 187946 22386
rect 185169 22328 185174 22384
rect 185230 22328 187946 22384
rect 185169 22326 187946 22328
rect 185169 22323 185235 22326
rect 177625 22250 177691 22253
rect 174852 22248 177691 22250
rect 174852 22192 177630 22248
rect 177686 22192 177691 22248
rect 174852 22190 177691 22192
rect 177625 22187 177691 22190
rect 187886 22152 187946 22326
rect 93905 22114 93971 22117
rect 90734 22112 93971 22114
rect 90734 22056 93910 22112
rect 93966 22056 93971 22112
rect 90734 22054 93971 22056
rect 51217 21978 51283 21981
rect 47862 21976 51283 21978
rect 47862 21920 51222 21976
rect 51278 21920 51283 21976
rect 47862 21918 51283 21920
rect 51217 21915 51283 21918
rect 50941 21842 51007 21845
rect 47862 21840 51007 21842
rect 47862 21784 50946 21840
rect 51002 21784 51007 21840
rect 47862 21782 51007 21784
rect 47862 21744 47922 21782
rect 50941 21779 51007 21782
rect 90734 21744 90794 22054
rect 93905 22051 93971 22054
rect 142481 22114 142547 22117
rect 142481 22112 145074 22114
rect 142481 22056 142486 22112
rect 142542 22056 145074 22112
rect 142481 22054 145074 22056
rect 142481 22051 142547 22054
rect 101081 21978 101147 21981
rect 135121 21978 135187 21981
rect 101081 21976 104042 21978
rect 101081 21920 101086 21976
rect 101142 21920 104042 21976
rect 101081 21918 104042 21920
rect 101081 21915 101147 21918
rect 58301 21706 58367 21709
rect 58301 21704 60956 21706
rect 58301 21648 58306 21704
rect 58362 21648 60956 21704
rect 58301 21646 60956 21648
rect 58301 21643 58367 21646
rect 103982 21476 104042 21918
rect 131766 21976 135187 21978
rect 131766 21920 135126 21976
rect 135182 21920 135187 21976
rect 131766 21918 135187 21920
rect 131766 21472 131826 21918
rect 135121 21915 135187 21918
rect 145014 21744 145074 22054
rect 185118 21916 185124 21980
rect 185188 21978 185194 21980
rect 185188 21918 187946 21978
rect 185188 21916 185194 21918
rect 177717 21706 177783 21709
rect 174852 21704 177783 21706
rect 174852 21648 177722 21704
rect 177778 21648 177783 21704
rect 174852 21646 177783 21648
rect 177717 21643 177783 21646
rect 187886 21472 187946 21918
rect 222286 21916 222292 21980
rect 222356 21978 222362 21980
rect 225416 21978 225896 22008
rect 222356 21918 225896 21978
rect 222356 21916 222362 21918
rect 225416 21888 225896 21918
rect 47862 21162 47922 21200
rect 50665 21162 50731 21165
rect 47862 21160 50731 21162
rect 47862 21104 50670 21160
rect 50726 21104 50731 21160
rect 47862 21102 50731 21104
rect 50665 21099 50731 21102
rect 58209 21162 58275 21165
rect 93997 21162 94063 21165
rect 134753 21162 134819 21165
rect 58209 21160 60956 21162
rect 58209 21104 58214 21160
rect 58270 21104 60956 21160
rect 58209 21102 60956 21104
rect 90764 21160 94063 21162
rect 90764 21104 94002 21160
rect 94058 21104 94063 21160
rect 90764 21102 94063 21104
rect 58209 21099 58275 21102
rect 93997 21099 94063 21102
rect 131766 21160 134819 21162
rect 131766 21104 134758 21160
rect 134814 21104 134819 21160
rect 131766 21102 134819 21104
rect 51033 21026 51099 21029
rect 47862 21024 51099 21026
rect 47862 20968 51038 21024
rect 51094 20968 51099 21024
rect 47862 20966 51099 20968
rect 47862 20656 47922 20966
rect 51033 20963 51099 20966
rect 61705 21026 61771 21029
rect 63177 21028 63243 21029
rect 62206 21026 62212 21028
rect 61705 21024 62212 21026
rect 61705 20968 61710 21024
rect 61766 20968 62212 21024
rect 61705 20966 62212 20968
rect 61705 20963 61771 20966
rect 62206 20964 62212 20966
rect 62276 20964 62282 21028
rect 63126 20964 63132 21028
rect 63196 21026 63243 21028
rect 64741 21028 64807 21029
rect 64741 21026 64788 21028
rect 63196 21024 63288 21026
rect 63238 20968 63288 21024
rect 63196 20966 63288 20968
rect 64696 21024 64788 21026
rect 64696 20968 64746 21024
rect 64696 20966 64788 20968
rect 63196 20964 63243 20966
rect 63177 20963 63243 20964
rect 64741 20964 64788 20966
rect 64852 20964 64858 21028
rect 64966 20964 64972 21028
rect 65036 21026 65042 21028
rect 65109 21026 65175 21029
rect 65036 21024 65175 21026
rect 65036 20968 65114 21024
rect 65170 20968 65175 21024
rect 65036 20966 65175 20968
rect 65036 20964 65042 20966
rect 64741 20963 64807 20964
rect 65109 20963 65175 20966
rect 131766 20928 131826 21102
rect 134753 21099 134819 21102
rect 143677 21162 143743 21165
rect 177717 21162 177783 21165
rect 143677 21160 145044 21162
rect 143677 21104 143682 21160
rect 143738 21104 145044 21160
rect 143677 21102 145044 21104
rect 174852 21160 177783 21162
rect 174852 21104 177722 21160
rect 177778 21104 177783 21160
rect 174852 21102 177783 21104
rect 143677 21099 143743 21102
rect 177717 21099 177783 21102
rect 146253 21028 146319 21029
rect 147725 21028 147791 21029
rect 146253 21026 146300 21028
rect 146208 21024 146300 21026
rect 146208 20968 146258 21024
rect 146208 20966 146300 20968
rect 146253 20964 146300 20966
rect 146364 20964 146370 21028
rect 147725 21026 147772 21028
rect 147680 21024 147772 21026
rect 147680 20968 147730 21024
rect 147680 20966 147772 20968
rect 147725 20964 147772 20966
rect 147836 20964 147842 21028
rect 148737 21026 148803 21029
rect 149054 21026 149060 21028
rect 148737 21024 149060 21026
rect 148737 20968 148742 21024
rect 148798 20968 149060 21024
rect 148737 20966 149060 20968
rect 146253 20963 146319 20964
rect 147725 20963 147791 20964
rect 148737 20963 148803 20966
rect 149054 20964 149060 20966
rect 149124 20964 149130 21028
rect 150853 21026 150919 21029
rect 156046 21026 156052 21028
rect 150853 21024 156052 21026
rect 150853 20968 150858 21024
rect 150914 20968 156052 21024
rect 150853 20966 156052 20968
rect 150853 20963 150919 20966
rect 156046 20964 156052 20966
rect 156116 20964 156122 21028
rect 62717 20890 62783 20893
rect 63310 20890 63316 20892
rect 62717 20888 63316 20890
rect 62717 20832 62722 20888
rect 62778 20832 63316 20888
rect 62717 20830 63316 20832
rect 62717 20827 62783 20830
rect 63310 20828 63316 20830
rect 63380 20828 63386 20892
rect 101582 20692 101588 20756
rect 101652 20754 101658 20756
rect 103982 20754 104042 20928
rect 145701 20890 145767 20893
rect 146110 20890 146116 20892
rect 145701 20888 146116 20890
rect 145701 20832 145706 20888
rect 145762 20832 146116 20888
rect 145701 20830 146116 20832
rect 145701 20827 145767 20830
rect 146110 20828 146116 20830
rect 146180 20828 146186 20892
rect 185486 20828 185492 20892
rect 185556 20890 185562 20892
rect 187886 20890 187946 20928
rect 185556 20830 187946 20890
rect 185556 20828 185562 20830
rect 135029 20754 135095 20757
rect 101652 20694 104042 20754
rect 131766 20752 135095 20754
rect 131766 20696 135034 20752
rect 135090 20696 135095 20752
rect 131766 20694 135095 20696
rect 101652 20692 101658 20694
rect 9896 20618 10376 20648
rect 13313 20618 13379 20621
rect 9896 20616 13379 20618
rect 9896 20560 13318 20616
rect 13374 20560 13379 20616
rect 9896 20558 13379 20560
rect 9896 20528 10376 20558
rect 13313 20555 13379 20558
rect 50849 20482 50915 20485
rect 47862 20480 50915 20482
rect 47862 20424 50854 20480
rect 50910 20424 50915 20480
rect 47862 20422 50915 20424
rect 47862 19976 47922 20422
rect 50849 20419 50915 20422
rect 131766 20248 131826 20694
rect 135029 20691 135095 20694
rect 185118 20692 185124 20756
rect 185188 20754 185194 20756
rect 185188 20694 187946 20754
rect 185188 20692 185194 20694
rect 187886 20248 187946 20694
rect 101582 20012 101588 20076
rect 101652 20074 101658 20076
rect 103982 20074 104042 20248
rect 101652 20014 104042 20074
rect 101652 20012 101658 20014
rect 50757 19802 50823 19805
rect 47862 19800 50823 19802
rect 47862 19744 50762 19800
rect 50818 19744 50823 19800
rect 47862 19742 50823 19744
rect 47862 19432 47922 19742
rect 50757 19739 50823 19742
rect 101541 19802 101607 19805
rect 134937 19802 135003 19805
rect 101541 19800 104042 19802
rect 101541 19744 101546 19800
rect 101602 19744 104042 19800
rect 101541 19742 104042 19744
rect 101541 19739 101607 19742
rect 103982 19708 104042 19742
rect 131766 19800 135003 19802
rect 131766 19744 134942 19800
rect 134998 19744 135003 19800
rect 131766 19742 135003 19744
rect 131766 19704 131826 19742
rect 134937 19739 135003 19742
rect 185169 19802 185235 19805
rect 185169 19800 187946 19802
rect 185169 19744 185174 19800
rect 185230 19744 187946 19800
rect 185169 19742 187946 19744
rect 185169 19739 185235 19742
rect 187886 19704 187946 19742
rect 101817 19530 101883 19533
rect 134477 19530 134543 19533
rect 101817 19528 104042 19530
rect 101817 19472 101822 19528
rect 101878 19472 104042 19528
rect 101817 19470 104042 19472
rect 101817 19467 101883 19470
rect 50573 19258 50639 19261
rect 47862 19256 50639 19258
rect 47862 19200 50578 19256
rect 50634 19200 50639 19256
rect 47862 19198 50639 19200
rect 47862 18888 47922 19198
rect 50573 19195 50639 19198
rect 103982 19164 104042 19470
rect 131766 19528 134543 19530
rect 131766 19472 134482 19528
rect 134538 19472 134543 19528
rect 131766 19470 134543 19472
rect 131766 19160 131826 19470
rect 134477 19467 134543 19470
rect 185261 19530 185327 19533
rect 185261 19528 187946 19530
rect 185261 19472 185266 19528
rect 185322 19472 187946 19528
rect 185261 19470 187946 19472
rect 185261 19467 185327 19470
rect 187886 19160 187946 19470
rect 212493 18444 212559 18445
rect 212493 18440 212540 18444
rect 212604 18442 212610 18444
rect 212493 18384 212498 18440
rect 212493 18380 212540 18384
rect 212604 18382 212650 18442
rect 212604 18380 212610 18382
rect 212493 18379 212559 18380
rect 63494 18244 63500 18308
rect 63564 18306 63570 18308
rect 66489 18306 66555 18309
rect 63564 18304 66555 18306
rect 63564 18248 66494 18304
rect 66550 18248 66555 18304
rect 63564 18246 66555 18248
rect 63564 18244 63570 18246
rect 66489 18243 66555 18246
rect 149749 18306 149815 18309
rect 151630 18306 151636 18308
rect 149749 18304 151636 18306
rect 149749 18248 149754 18304
rect 149810 18248 151636 18304
rect 149749 18246 151636 18248
rect 149749 18243 149815 18246
rect 151630 18244 151636 18246
rect 151700 18244 151706 18308
rect 129049 17082 129115 17085
rect 147030 17082 147036 17084
rect 129049 17080 147036 17082
rect 129049 17024 129054 17080
rect 129110 17024 147036 17080
rect 129049 17022 147036 17024
rect 129049 17019 129115 17022
rect 147030 17020 147036 17022
rect 147100 17020 147106 17084
<< via3 >>
rect 189172 236524 189236 236588
rect 88524 235164 88588 235228
rect 171140 232580 171204 232644
rect 171140 208916 171204 208980
rect 88524 207420 88588 207484
rect 189172 206876 189236 206940
rect 140228 195180 140292 195244
rect 209964 190752 210028 190756
rect 209964 190696 209978 190752
rect 209978 190696 210028 190752
rect 209964 190692 210028 190696
rect 193956 190556 194020 190620
rect 138020 156692 138084 156756
rect 209780 156692 209844 156756
rect 193772 96852 193836 96916
rect 209780 96716 209844 96780
rect 13268 67748 13332 67812
rect 212356 63124 212420 63188
rect 140228 58364 140292 58428
rect 55956 58228 56020 58292
rect 64972 46804 65036 46868
rect 159548 46804 159612 46868
rect 63500 46668 63564 46732
rect 149060 46668 149124 46732
rect 62212 46532 62276 46596
rect 146300 46532 146364 46596
rect 63132 46396 63196 46460
rect 63316 46260 63380 46324
rect 89812 46260 89876 46324
rect 64788 46124 64852 46188
rect 89076 46124 89140 46188
rect 147772 46396 147836 46460
rect 146116 46260 146180 46324
rect 147036 46124 147100 46188
rect 154948 45988 155012 46052
rect 173164 46260 173228 46324
rect 173532 46124 173596 46188
rect 173900 44628 173964 44692
rect 185124 21916 185188 21980
rect 222292 21916 222356 21980
rect 62212 20964 62276 21028
rect 63132 21024 63196 21028
rect 63132 20968 63182 21024
rect 63182 20968 63196 21024
rect 63132 20964 63196 20968
rect 64788 21024 64852 21028
rect 64788 20968 64802 21024
rect 64802 20968 64852 21024
rect 64788 20964 64852 20968
rect 64972 20964 65036 21028
rect 146300 21024 146364 21028
rect 146300 20968 146314 21024
rect 146314 20968 146364 21024
rect 146300 20964 146364 20968
rect 147772 21024 147836 21028
rect 147772 20968 147786 21024
rect 147786 20968 147836 21024
rect 147772 20964 147836 20968
rect 149060 20964 149124 21028
rect 156052 20964 156116 21028
rect 63316 20828 63380 20892
rect 101588 20692 101652 20756
rect 146116 20828 146180 20892
rect 185492 20828 185556 20892
rect 185124 20692 185188 20756
rect 101588 20012 101652 20076
rect 212540 18440 212604 18444
rect 212540 18384 212554 18440
rect 212554 18384 212604 18440
rect 212540 18380 212604 18384
rect 63500 18244 63564 18308
rect 151636 18244 151700 18308
rect 147036 17020 147100 17084
<< metal4 >>
rect 0 253078 4000 253200
rect 0 252842 122 253078
rect 358 252842 442 253078
rect 678 252842 762 253078
rect 998 252842 1082 253078
rect 1318 252842 1402 253078
rect 1638 252842 1722 253078
rect 1958 252842 2042 253078
rect 2278 252842 2362 253078
rect 2598 252842 2682 253078
rect 2918 252842 3002 253078
rect 3238 252842 3322 253078
rect 3558 252842 3642 253078
rect 3878 252842 4000 253078
rect 0 252758 4000 252842
rect 0 252522 122 252758
rect 358 252522 442 252758
rect 678 252522 762 252758
rect 998 252522 1082 252758
rect 1318 252522 1402 252758
rect 1638 252522 1722 252758
rect 1958 252522 2042 252758
rect 2278 252522 2362 252758
rect 2598 252522 2682 252758
rect 2918 252522 3002 252758
rect 3238 252522 3322 252758
rect 3558 252522 3642 252758
rect 3878 252522 4000 252758
rect 0 252438 4000 252522
rect 0 252202 122 252438
rect 358 252202 442 252438
rect 678 252202 762 252438
rect 998 252202 1082 252438
rect 1318 252202 1402 252438
rect 1638 252202 1722 252438
rect 1958 252202 2042 252438
rect 2278 252202 2362 252438
rect 2598 252202 2682 252438
rect 2918 252202 3002 252438
rect 3238 252202 3322 252438
rect 3558 252202 3642 252438
rect 3878 252202 4000 252438
rect 0 252118 4000 252202
rect 0 251882 122 252118
rect 358 251882 442 252118
rect 678 251882 762 252118
rect 998 251882 1082 252118
rect 1318 251882 1402 252118
rect 1638 251882 1722 252118
rect 1958 251882 2042 252118
rect 2278 251882 2362 252118
rect 2598 251882 2682 252118
rect 2918 251882 3002 252118
rect 3238 251882 3322 252118
rect 3558 251882 3642 252118
rect 3878 251882 4000 252118
rect 0 251798 4000 251882
rect 0 251562 122 251798
rect 358 251562 442 251798
rect 678 251562 762 251798
rect 998 251562 1082 251798
rect 1318 251562 1402 251798
rect 1638 251562 1722 251798
rect 1958 251562 2042 251798
rect 2278 251562 2362 251798
rect 2598 251562 2682 251798
rect 2918 251562 3002 251798
rect 3238 251562 3322 251798
rect 3558 251562 3642 251798
rect 3878 251562 4000 251798
rect 0 251478 4000 251562
rect 0 251242 122 251478
rect 358 251242 442 251478
rect 678 251242 762 251478
rect 998 251242 1082 251478
rect 1318 251242 1402 251478
rect 1638 251242 1722 251478
rect 1958 251242 2042 251478
rect 2278 251242 2362 251478
rect 2598 251242 2682 251478
rect 2918 251242 3002 251478
rect 3238 251242 3322 251478
rect 3558 251242 3642 251478
rect 3878 251242 4000 251478
rect 0 251158 4000 251242
rect 0 250922 122 251158
rect 358 250922 442 251158
rect 678 250922 762 251158
rect 998 250922 1082 251158
rect 1318 250922 1402 251158
rect 1638 250922 1722 251158
rect 1958 250922 2042 251158
rect 2278 250922 2362 251158
rect 2598 250922 2682 251158
rect 2918 250922 3002 251158
rect 3238 250922 3322 251158
rect 3558 250922 3642 251158
rect 3878 250922 4000 251158
rect 0 250838 4000 250922
rect 0 250602 122 250838
rect 358 250602 442 250838
rect 678 250602 762 250838
rect 998 250602 1082 250838
rect 1318 250602 1402 250838
rect 1638 250602 1722 250838
rect 1958 250602 2042 250838
rect 2278 250602 2362 250838
rect 2598 250602 2682 250838
rect 2918 250602 3002 250838
rect 3238 250602 3322 250838
rect 3558 250602 3642 250838
rect 3878 250602 4000 250838
rect 0 250518 4000 250602
rect 0 250282 122 250518
rect 358 250282 442 250518
rect 678 250282 762 250518
rect 998 250282 1082 250518
rect 1318 250282 1402 250518
rect 1638 250282 1722 250518
rect 1958 250282 2042 250518
rect 2278 250282 2362 250518
rect 2598 250282 2682 250518
rect 2918 250282 3002 250518
rect 3238 250282 3322 250518
rect 3558 250282 3642 250518
rect 3878 250282 4000 250518
rect 0 250198 4000 250282
rect 0 249962 122 250198
rect 358 249962 442 250198
rect 678 249962 762 250198
rect 998 249962 1082 250198
rect 1318 249962 1402 250198
rect 1638 249962 1722 250198
rect 1958 249962 2042 250198
rect 2278 249962 2362 250198
rect 2598 249962 2682 250198
rect 2918 249962 3002 250198
rect 3238 249962 3322 250198
rect 3558 249962 3642 250198
rect 3878 249962 4000 250198
rect 0 249878 4000 249962
rect 0 249642 122 249878
rect 358 249642 442 249878
rect 678 249642 762 249878
rect 998 249642 1082 249878
rect 1318 249642 1402 249878
rect 1638 249642 1722 249878
rect 1958 249642 2042 249878
rect 2278 249642 2362 249878
rect 2598 249642 2682 249878
rect 2918 249642 3002 249878
rect 3238 249642 3322 249878
rect 3558 249642 3642 249878
rect 3878 249642 4000 249878
rect 0 249558 4000 249642
rect 0 249322 122 249558
rect 358 249322 442 249558
rect 678 249322 762 249558
rect 998 249322 1082 249558
rect 1318 249322 1402 249558
rect 1638 249322 1722 249558
rect 1958 249322 2042 249558
rect 2278 249322 2362 249558
rect 2598 249322 2682 249558
rect 2918 249322 3002 249558
rect 3238 249322 3322 249558
rect 3558 249322 3642 249558
rect 3878 249322 4000 249558
rect 0 228918 4000 249322
rect 231716 253078 235716 253200
rect 231716 252842 231838 253078
rect 232074 252842 232158 253078
rect 232394 252842 232478 253078
rect 232714 252842 232798 253078
rect 233034 252842 233118 253078
rect 233354 252842 233438 253078
rect 233674 252842 233758 253078
rect 233994 252842 234078 253078
rect 234314 252842 234398 253078
rect 234634 252842 234718 253078
rect 234954 252842 235038 253078
rect 235274 252842 235358 253078
rect 235594 252842 235716 253078
rect 231716 252758 235716 252842
rect 231716 252522 231838 252758
rect 232074 252522 232158 252758
rect 232394 252522 232478 252758
rect 232714 252522 232798 252758
rect 233034 252522 233118 252758
rect 233354 252522 233438 252758
rect 233674 252522 233758 252758
rect 233994 252522 234078 252758
rect 234314 252522 234398 252758
rect 234634 252522 234718 252758
rect 234954 252522 235038 252758
rect 235274 252522 235358 252758
rect 235594 252522 235716 252758
rect 231716 252438 235716 252522
rect 231716 252202 231838 252438
rect 232074 252202 232158 252438
rect 232394 252202 232478 252438
rect 232714 252202 232798 252438
rect 233034 252202 233118 252438
rect 233354 252202 233438 252438
rect 233674 252202 233758 252438
rect 233994 252202 234078 252438
rect 234314 252202 234398 252438
rect 234634 252202 234718 252438
rect 234954 252202 235038 252438
rect 235274 252202 235358 252438
rect 235594 252202 235716 252438
rect 231716 252118 235716 252202
rect 231716 251882 231838 252118
rect 232074 251882 232158 252118
rect 232394 251882 232478 252118
rect 232714 251882 232798 252118
rect 233034 251882 233118 252118
rect 233354 251882 233438 252118
rect 233674 251882 233758 252118
rect 233994 251882 234078 252118
rect 234314 251882 234398 252118
rect 234634 251882 234718 252118
rect 234954 251882 235038 252118
rect 235274 251882 235358 252118
rect 235594 251882 235716 252118
rect 231716 251798 235716 251882
rect 231716 251562 231838 251798
rect 232074 251562 232158 251798
rect 232394 251562 232478 251798
rect 232714 251562 232798 251798
rect 233034 251562 233118 251798
rect 233354 251562 233438 251798
rect 233674 251562 233758 251798
rect 233994 251562 234078 251798
rect 234314 251562 234398 251798
rect 234634 251562 234718 251798
rect 234954 251562 235038 251798
rect 235274 251562 235358 251798
rect 235594 251562 235716 251798
rect 231716 251478 235716 251562
rect 231716 251242 231838 251478
rect 232074 251242 232158 251478
rect 232394 251242 232478 251478
rect 232714 251242 232798 251478
rect 233034 251242 233118 251478
rect 233354 251242 233438 251478
rect 233674 251242 233758 251478
rect 233994 251242 234078 251478
rect 234314 251242 234398 251478
rect 234634 251242 234718 251478
rect 234954 251242 235038 251478
rect 235274 251242 235358 251478
rect 235594 251242 235716 251478
rect 231716 251158 235716 251242
rect 231716 250922 231838 251158
rect 232074 250922 232158 251158
rect 232394 250922 232478 251158
rect 232714 250922 232798 251158
rect 233034 250922 233118 251158
rect 233354 250922 233438 251158
rect 233674 250922 233758 251158
rect 233994 250922 234078 251158
rect 234314 250922 234398 251158
rect 234634 250922 234718 251158
rect 234954 250922 235038 251158
rect 235274 250922 235358 251158
rect 235594 250922 235716 251158
rect 231716 250838 235716 250922
rect 231716 250602 231838 250838
rect 232074 250602 232158 250838
rect 232394 250602 232478 250838
rect 232714 250602 232798 250838
rect 233034 250602 233118 250838
rect 233354 250602 233438 250838
rect 233674 250602 233758 250838
rect 233994 250602 234078 250838
rect 234314 250602 234398 250838
rect 234634 250602 234718 250838
rect 234954 250602 235038 250838
rect 235274 250602 235358 250838
rect 235594 250602 235716 250838
rect 231716 250518 235716 250602
rect 231716 250282 231838 250518
rect 232074 250282 232158 250518
rect 232394 250282 232478 250518
rect 232714 250282 232798 250518
rect 233034 250282 233118 250518
rect 233354 250282 233438 250518
rect 233674 250282 233758 250518
rect 233994 250282 234078 250518
rect 234314 250282 234398 250518
rect 234634 250282 234718 250518
rect 234954 250282 235038 250518
rect 235274 250282 235358 250518
rect 235594 250282 235716 250518
rect 231716 250198 235716 250282
rect 231716 249962 231838 250198
rect 232074 249962 232158 250198
rect 232394 249962 232478 250198
rect 232714 249962 232798 250198
rect 233034 249962 233118 250198
rect 233354 249962 233438 250198
rect 233674 249962 233758 250198
rect 233994 249962 234078 250198
rect 234314 249962 234398 250198
rect 234634 249962 234718 250198
rect 234954 249962 235038 250198
rect 235274 249962 235358 250198
rect 235594 249962 235716 250198
rect 231716 249878 235716 249962
rect 231716 249642 231838 249878
rect 232074 249642 232158 249878
rect 232394 249642 232478 249878
rect 232714 249642 232798 249878
rect 233034 249642 233118 249878
rect 233354 249642 233438 249878
rect 233674 249642 233758 249878
rect 233994 249642 234078 249878
rect 234314 249642 234398 249878
rect 234634 249642 234718 249878
rect 234954 249642 235038 249878
rect 235274 249642 235358 249878
rect 235594 249642 235716 249878
rect 231716 249558 235716 249642
rect 231716 249322 231838 249558
rect 232074 249322 232158 249558
rect 232394 249322 232478 249558
rect 232714 249322 232798 249558
rect 233034 249322 233118 249558
rect 233354 249322 233438 249558
rect 233674 249322 233758 249558
rect 233994 249322 234078 249558
rect 234314 249322 234398 249558
rect 234634 249322 234718 249558
rect 234954 249322 235038 249558
rect 235274 249322 235358 249558
rect 235594 249322 235716 249558
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 4000 228918
rect 0 206518 4000 228682
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 4000 206518
rect 0 184118 4000 206282
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 4000 184118
rect 0 161718 4000 183882
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 4000 161718
rect 0 139318 4000 161482
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 4000 139318
rect 0 116918 4000 139082
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 4000 116918
rect 0 94518 4000 116682
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 4000 94518
rect 0 72118 4000 94282
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 4000 72118
rect 0 49718 4000 71882
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 4000 49718
rect 0 27318 4000 49482
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 4000 27318
rect 0 3878 4000 27082
rect 5000 248078 9000 248200
rect 5000 247842 5122 248078
rect 5358 247842 5442 248078
rect 5678 247842 5762 248078
rect 5998 247842 6082 248078
rect 6318 247842 6402 248078
rect 6638 247842 6722 248078
rect 6958 247842 7042 248078
rect 7278 247842 7362 248078
rect 7598 247842 7682 248078
rect 7918 247842 8002 248078
rect 8238 247842 8322 248078
rect 8558 247842 8642 248078
rect 8878 247842 9000 248078
rect 5000 247758 9000 247842
rect 5000 247522 5122 247758
rect 5358 247522 5442 247758
rect 5678 247522 5762 247758
rect 5998 247522 6082 247758
rect 6318 247522 6402 247758
rect 6638 247522 6722 247758
rect 6958 247522 7042 247758
rect 7278 247522 7362 247758
rect 7598 247522 7682 247758
rect 7918 247522 8002 247758
rect 8238 247522 8322 247758
rect 8558 247522 8642 247758
rect 8878 247522 9000 247758
rect 5000 247438 9000 247522
rect 5000 247202 5122 247438
rect 5358 247202 5442 247438
rect 5678 247202 5762 247438
rect 5998 247202 6082 247438
rect 6318 247202 6402 247438
rect 6638 247202 6722 247438
rect 6958 247202 7042 247438
rect 7278 247202 7362 247438
rect 7598 247202 7682 247438
rect 7918 247202 8002 247438
rect 8238 247202 8322 247438
rect 8558 247202 8642 247438
rect 8878 247202 9000 247438
rect 5000 247118 9000 247202
rect 5000 246882 5122 247118
rect 5358 246882 5442 247118
rect 5678 246882 5762 247118
rect 5998 246882 6082 247118
rect 6318 246882 6402 247118
rect 6638 246882 6722 247118
rect 6958 246882 7042 247118
rect 7278 246882 7362 247118
rect 7598 246882 7682 247118
rect 7918 246882 8002 247118
rect 8238 246882 8322 247118
rect 8558 246882 8642 247118
rect 8878 246882 9000 247118
rect 5000 246798 9000 246882
rect 5000 246562 5122 246798
rect 5358 246562 5442 246798
rect 5678 246562 5762 246798
rect 5998 246562 6082 246798
rect 6318 246562 6402 246798
rect 6638 246562 6722 246798
rect 6958 246562 7042 246798
rect 7278 246562 7362 246798
rect 7598 246562 7682 246798
rect 7918 246562 8002 246798
rect 8238 246562 8322 246798
rect 8558 246562 8642 246798
rect 8878 246562 9000 246798
rect 5000 246478 9000 246562
rect 5000 246242 5122 246478
rect 5358 246242 5442 246478
rect 5678 246242 5762 246478
rect 5998 246242 6082 246478
rect 6318 246242 6402 246478
rect 6638 246242 6722 246478
rect 6958 246242 7042 246478
rect 7278 246242 7362 246478
rect 7598 246242 7682 246478
rect 7918 246242 8002 246478
rect 8238 246242 8322 246478
rect 8558 246242 8642 246478
rect 8878 246242 9000 246478
rect 5000 246158 9000 246242
rect 5000 245922 5122 246158
rect 5358 245922 5442 246158
rect 5678 245922 5762 246158
rect 5998 245922 6082 246158
rect 6318 245922 6402 246158
rect 6638 245922 6722 246158
rect 6958 245922 7042 246158
rect 7278 245922 7362 246158
rect 7598 245922 7682 246158
rect 7918 245922 8002 246158
rect 8238 245922 8322 246158
rect 8558 245922 8642 246158
rect 8878 245922 9000 246158
rect 5000 245838 9000 245922
rect 5000 245602 5122 245838
rect 5358 245602 5442 245838
rect 5678 245602 5762 245838
rect 5998 245602 6082 245838
rect 6318 245602 6402 245838
rect 6638 245602 6722 245838
rect 6958 245602 7042 245838
rect 7278 245602 7362 245838
rect 7598 245602 7682 245838
rect 7918 245602 8002 245838
rect 8238 245602 8322 245838
rect 8558 245602 8642 245838
rect 8878 245602 9000 245838
rect 5000 245518 9000 245602
rect 5000 245282 5122 245518
rect 5358 245282 5442 245518
rect 5678 245282 5762 245518
rect 5998 245282 6082 245518
rect 6318 245282 6402 245518
rect 6638 245282 6722 245518
rect 6958 245282 7042 245518
rect 7278 245282 7362 245518
rect 7598 245282 7682 245518
rect 7918 245282 8002 245518
rect 8238 245282 8322 245518
rect 8558 245282 8642 245518
rect 8878 245282 9000 245518
rect 5000 245198 9000 245282
rect 5000 244962 5122 245198
rect 5358 244962 5442 245198
rect 5678 244962 5762 245198
rect 5998 244962 6082 245198
rect 6318 244962 6402 245198
rect 6638 244962 6722 245198
rect 6958 244962 7042 245198
rect 7278 244962 7362 245198
rect 7598 244962 7682 245198
rect 7918 244962 8002 245198
rect 8238 244962 8322 245198
rect 8558 244962 8642 245198
rect 8878 244962 9000 245198
rect 5000 244878 9000 244962
rect 5000 244642 5122 244878
rect 5358 244642 5442 244878
rect 5678 244642 5762 244878
rect 5998 244642 6082 244878
rect 6318 244642 6402 244878
rect 6638 244642 6722 244878
rect 6958 244642 7042 244878
rect 7278 244642 7362 244878
rect 7598 244642 7682 244878
rect 7918 244642 8002 244878
rect 8238 244642 8322 244878
rect 8558 244642 8642 244878
rect 8878 244642 9000 244878
rect 5000 244558 9000 244642
rect 5000 244322 5122 244558
rect 5358 244322 5442 244558
rect 5678 244322 5762 244558
rect 5998 244322 6082 244558
rect 6318 244322 6402 244558
rect 6638 244322 6722 244558
rect 6958 244322 7042 244558
rect 7278 244322 7362 244558
rect 7598 244322 7682 244558
rect 7918 244322 8002 244558
rect 8238 244322 8322 244558
rect 8558 244322 8642 244558
rect 8878 244322 9000 244558
rect 5000 240118 9000 244322
rect 5000 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 9000 240118
rect 5000 217718 9000 239882
rect 226716 248078 230716 248200
rect 226716 247842 226838 248078
rect 227074 247842 227158 248078
rect 227394 247842 227478 248078
rect 227714 247842 227798 248078
rect 228034 247842 228118 248078
rect 228354 247842 228438 248078
rect 228674 247842 228758 248078
rect 228994 247842 229078 248078
rect 229314 247842 229398 248078
rect 229634 247842 229718 248078
rect 229954 247842 230038 248078
rect 230274 247842 230358 248078
rect 230594 247842 230716 248078
rect 226716 247758 230716 247842
rect 226716 247522 226838 247758
rect 227074 247522 227158 247758
rect 227394 247522 227478 247758
rect 227714 247522 227798 247758
rect 228034 247522 228118 247758
rect 228354 247522 228438 247758
rect 228674 247522 228758 247758
rect 228994 247522 229078 247758
rect 229314 247522 229398 247758
rect 229634 247522 229718 247758
rect 229954 247522 230038 247758
rect 230274 247522 230358 247758
rect 230594 247522 230716 247758
rect 226716 247438 230716 247522
rect 226716 247202 226838 247438
rect 227074 247202 227158 247438
rect 227394 247202 227478 247438
rect 227714 247202 227798 247438
rect 228034 247202 228118 247438
rect 228354 247202 228438 247438
rect 228674 247202 228758 247438
rect 228994 247202 229078 247438
rect 229314 247202 229398 247438
rect 229634 247202 229718 247438
rect 229954 247202 230038 247438
rect 230274 247202 230358 247438
rect 230594 247202 230716 247438
rect 226716 247118 230716 247202
rect 226716 246882 226838 247118
rect 227074 246882 227158 247118
rect 227394 246882 227478 247118
rect 227714 246882 227798 247118
rect 228034 246882 228118 247118
rect 228354 246882 228438 247118
rect 228674 246882 228758 247118
rect 228994 246882 229078 247118
rect 229314 246882 229398 247118
rect 229634 246882 229718 247118
rect 229954 246882 230038 247118
rect 230274 246882 230358 247118
rect 230594 246882 230716 247118
rect 226716 246798 230716 246882
rect 226716 246562 226838 246798
rect 227074 246562 227158 246798
rect 227394 246562 227478 246798
rect 227714 246562 227798 246798
rect 228034 246562 228118 246798
rect 228354 246562 228438 246798
rect 228674 246562 228758 246798
rect 228994 246562 229078 246798
rect 229314 246562 229398 246798
rect 229634 246562 229718 246798
rect 229954 246562 230038 246798
rect 230274 246562 230358 246798
rect 230594 246562 230716 246798
rect 226716 246478 230716 246562
rect 226716 246242 226838 246478
rect 227074 246242 227158 246478
rect 227394 246242 227478 246478
rect 227714 246242 227798 246478
rect 228034 246242 228118 246478
rect 228354 246242 228438 246478
rect 228674 246242 228758 246478
rect 228994 246242 229078 246478
rect 229314 246242 229398 246478
rect 229634 246242 229718 246478
rect 229954 246242 230038 246478
rect 230274 246242 230358 246478
rect 230594 246242 230716 246478
rect 226716 246158 230716 246242
rect 226716 245922 226838 246158
rect 227074 245922 227158 246158
rect 227394 245922 227478 246158
rect 227714 245922 227798 246158
rect 228034 245922 228118 246158
rect 228354 245922 228438 246158
rect 228674 245922 228758 246158
rect 228994 245922 229078 246158
rect 229314 245922 229398 246158
rect 229634 245922 229718 246158
rect 229954 245922 230038 246158
rect 230274 245922 230358 246158
rect 230594 245922 230716 246158
rect 226716 245838 230716 245922
rect 226716 245602 226838 245838
rect 227074 245602 227158 245838
rect 227394 245602 227478 245838
rect 227714 245602 227798 245838
rect 228034 245602 228118 245838
rect 228354 245602 228438 245838
rect 228674 245602 228758 245838
rect 228994 245602 229078 245838
rect 229314 245602 229398 245838
rect 229634 245602 229718 245838
rect 229954 245602 230038 245838
rect 230274 245602 230358 245838
rect 230594 245602 230716 245838
rect 226716 245518 230716 245602
rect 226716 245282 226838 245518
rect 227074 245282 227158 245518
rect 227394 245282 227478 245518
rect 227714 245282 227798 245518
rect 228034 245282 228118 245518
rect 228354 245282 228438 245518
rect 228674 245282 228758 245518
rect 228994 245282 229078 245518
rect 229314 245282 229398 245518
rect 229634 245282 229718 245518
rect 229954 245282 230038 245518
rect 230274 245282 230358 245518
rect 230594 245282 230716 245518
rect 226716 245198 230716 245282
rect 226716 244962 226838 245198
rect 227074 244962 227158 245198
rect 227394 244962 227478 245198
rect 227714 244962 227798 245198
rect 228034 244962 228118 245198
rect 228354 244962 228438 245198
rect 228674 244962 228758 245198
rect 228994 244962 229078 245198
rect 229314 244962 229398 245198
rect 229634 244962 229718 245198
rect 229954 244962 230038 245198
rect 230274 244962 230358 245198
rect 230594 244962 230716 245198
rect 226716 244878 230716 244962
rect 226716 244642 226838 244878
rect 227074 244642 227158 244878
rect 227394 244642 227478 244878
rect 227714 244642 227798 244878
rect 228034 244642 228118 244878
rect 228354 244642 228438 244878
rect 228674 244642 228758 244878
rect 228994 244642 229078 244878
rect 229314 244642 229398 244878
rect 229634 244642 229718 244878
rect 229954 244642 230038 244878
rect 230274 244642 230358 244878
rect 230594 244642 230716 244878
rect 226716 244558 230716 244642
rect 226716 244322 226838 244558
rect 227074 244322 227158 244558
rect 227394 244322 227478 244558
rect 227714 244322 227798 244558
rect 228034 244322 228118 244558
rect 228354 244322 228438 244558
rect 228674 244322 228758 244558
rect 228994 244322 229078 244558
rect 229314 244322 229398 244558
rect 229634 244322 229718 244558
rect 229954 244322 230038 244558
rect 230274 244322 230358 244558
rect 230594 244322 230716 244558
rect 226716 240118 230716 244322
rect 226716 239882 226838 240118
rect 227074 239882 227158 240118
rect 227394 239882 227478 240118
rect 227714 239882 227798 240118
rect 228034 239882 228118 240118
rect 228354 239882 228438 240118
rect 228674 239882 228758 240118
rect 228994 239882 229078 240118
rect 229314 239882 229398 240118
rect 229634 239882 229718 240118
rect 229954 239882 230038 240118
rect 230274 239882 230358 240118
rect 230594 239882 230716 240118
rect 189171 236588 189237 236589
rect 189171 236524 189172 236588
rect 189236 236524 189237 236588
rect 189171 236523 189237 236524
rect 88523 235228 88589 235229
rect 88523 235164 88524 235228
rect 88588 235164 88589 235228
rect 88523 235163 88589 235164
rect 30173 228918 30493 228960
rect 30173 228682 30215 228918
rect 30451 228682 30493 228918
rect 30173 228640 30493 228682
rect 71840 228918 72160 228960
rect 71840 228682 71882 228918
rect 72118 228682 72160 228918
rect 71840 228640 72160 228682
rect 5000 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 9000 217718
rect 5000 195318 9000 217482
rect 25507 217718 25827 217760
rect 25507 217482 25549 217718
rect 25785 217482 25827 217718
rect 25507 217440 25827 217482
rect 66840 217718 67160 217760
rect 66840 217482 66882 217718
rect 67118 217482 67160 217718
rect 66840 217440 67160 217482
rect 88526 207485 88586 235163
rect 171139 232644 171205 232645
rect 171139 232580 171140 232644
rect 171204 232580 171205 232644
rect 171139 232579 171205 232580
rect 171142 230874 171202 232579
rect 171142 230814 171570 230874
rect 114173 228918 114493 228960
rect 114173 228682 114215 228918
rect 114451 228682 114493 228918
rect 114173 228640 114493 228682
rect 155840 228918 156160 228960
rect 155840 228682 155882 228918
rect 156118 228682 156160 228918
rect 155840 228640 156160 228682
rect 109507 217718 109827 217760
rect 109507 217482 109549 217718
rect 109785 217482 109827 217718
rect 109507 217440 109827 217482
rect 150840 217718 151160 217760
rect 150840 217482 150882 217718
rect 151118 217482 151160 217718
rect 150840 217440 151160 217482
rect 171510 213874 171570 230814
rect 171326 213814 171570 213874
rect 171326 210474 171386 213814
rect 171142 210414 171386 210474
rect 171142 208981 171202 210414
rect 171139 208980 171205 208981
rect 171139 208916 171140 208980
rect 171204 208916 171205 208980
rect 171139 208915 171205 208916
rect 88523 207484 88589 207485
rect 88523 207420 88524 207484
rect 88588 207420 88589 207484
rect 88523 207419 88589 207420
rect 189174 206941 189234 236523
rect 198173 228918 198493 228960
rect 198173 228682 198215 228918
rect 198451 228682 198493 228918
rect 198173 228640 198493 228682
rect 193507 217718 193827 217760
rect 193507 217482 193549 217718
rect 193785 217482 193827 217718
rect 193507 217440 193827 217482
rect 226716 217718 230716 239882
rect 226716 217482 226838 217718
rect 227074 217482 227158 217718
rect 227394 217482 227478 217718
rect 227714 217482 227798 217718
rect 228034 217482 228118 217718
rect 228354 217482 228438 217718
rect 228674 217482 228758 217718
rect 228994 217482 229078 217718
rect 229314 217482 229398 217718
rect 229634 217482 229718 217718
rect 229954 217482 230038 217718
rect 230274 217482 230358 217718
rect 230594 217482 230716 217718
rect 189171 206940 189237 206941
rect 189171 206876 189172 206940
rect 189236 206876 189237 206940
rect 189171 206875 189237 206876
rect 5000 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 9000 195318
rect 226716 195318 230716 217482
rect 140227 195244 140293 195245
rect 140227 195180 140228 195244
rect 140292 195180 140293 195244
rect 140227 195179 140293 195180
rect 5000 172918 9000 195082
rect 32173 184118 32493 184160
rect 32173 183882 32215 184118
rect 32451 183882 32493 184118
rect 32173 183840 32493 183882
rect 75464 184118 75784 184160
rect 75464 183882 75506 184118
rect 75742 183882 75784 184118
rect 75464 183840 75784 183882
rect 116173 184118 116493 184160
rect 116173 183882 116215 184118
rect 116451 183882 116493 184118
rect 116173 183840 116493 183882
rect 5000 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 9000 172918
rect 5000 150518 9000 172682
rect 29507 172918 29827 172960
rect 29507 172682 29549 172918
rect 29785 172682 29827 172918
rect 29507 172640 29827 172682
rect 60104 172918 60424 172960
rect 60104 172682 60146 172918
rect 60382 172682 60424 172918
rect 60104 172640 60424 172682
rect 113507 172918 113827 172960
rect 113507 172682 113549 172918
rect 113785 172682 113827 172918
rect 113507 172640 113827 172682
rect 32173 161718 32493 161760
rect 32173 161482 32215 161718
rect 32451 161482 32493 161718
rect 32173 161440 32493 161482
rect 75464 161718 75784 161760
rect 75464 161482 75506 161718
rect 75742 161482 75784 161718
rect 75464 161440 75784 161482
rect 116173 161718 116493 161760
rect 116173 161482 116215 161718
rect 116451 161482 116493 161718
rect 116173 161440 116493 161482
rect 5000 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 9000 150518
rect 5000 128118 9000 150282
rect 5000 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 9000 128118
rect 5000 105718 9000 127882
rect 25507 128118 25827 128160
rect 25507 127882 25549 128118
rect 25785 127882 25827 128118
rect 25507 127840 25827 127882
rect 66840 128118 67160 128160
rect 66840 127882 66882 128118
rect 67118 127882 67160 128118
rect 66840 127840 67160 127882
rect 109507 128118 109827 128160
rect 109507 127882 109549 128118
rect 109785 127882 109827 128118
rect 109507 127840 109827 127882
rect 30173 116918 30493 116960
rect 30173 116682 30215 116918
rect 30451 116682 30493 116918
rect 30173 116640 30493 116682
rect 114173 116918 114493 116960
rect 114173 116682 114215 116918
rect 114451 116682 114493 116918
rect 114173 116640 114493 116682
rect 5000 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 9000 105718
rect 5000 83318 9000 105482
rect 32173 94518 32493 94560
rect 32173 94282 32215 94518
rect 32451 94282 32493 94518
rect 32173 94240 32493 94282
rect 75464 94518 75784 94560
rect 75464 94282 75506 94518
rect 75742 94282 75784 94518
rect 75464 94240 75784 94282
rect 116173 94518 116493 94560
rect 116173 94282 116215 94518
rect 116451 94282 116493 94518
rect 116173 94240 116493 94282
rect 5000 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 9000 83318
rect 5000 60918 9000 83082
rect 29507 83318 29827 83360
rect 29507 83082 29549 83318
rect 29785 83082 29827 83318
rect 29507 83040 29827 83082
rect 60104 83318 60424 83360
rect 60104 83082 60146 83318
rect 60382 83082 60424 83318
rect 60104 83040 60424 83082
rect 113507 83318 113827 83360
rect 113507 83082 113549 83318
rect 113785 83082 113827 83318
rect 113507 83040 113827 83082
rect 32173 72118 32493 72160
rect 32173 71882 32215 72118
rect 32451 71882 32493 72118
rect 32173 71840 32493 71882
rect 75464 72118 75784 72160
rect 75464 71882 75506 72118
rect 75742 71882 75784 72118
rect 75464 71840 75784 71882
rect 116173 72118 116493 72160
rect 116173 71882 116215 72118
rect 116451 71882 116493 72118
rect 116173 71840 116493 71882
rect 13267 67812 13333 67813
rect 13267 67748 13268 67812
rect 13332 67748 13333 67812
rect 13267 67747 13333 67748
rect 13270 67082 13330 67747
rect 5000 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 9000 60918
rect 5000 38518 9000 60682
rect 55958 58293 56018 66846
rect 140230 58429 140290 195179
rect 226716 195082 226838 195318
rect 227074 195082 227158 195318
rect 227394 195082 227478 195318
rect 227714 195082 227798 195318
rect 228034 195082 228118 195318
rect 228354 195082 228438 195318
rect 228674 195082 228758 195318
rect 228994 195082 229078 195318
rect 229314 195082 229398 195318
rect 229634 195082 229718 195318
rect 229954 195082 230038 195318
rect 230274 195082 230358 195318
rect 230594 195082 230716 195318
rect 193955 190556 193956 190606
rect 194020 190556 194021 190606
rect 193955 190555 194021 190556
rect 159464 184118 159784 184160
rect 159464 183882 159506 184118
rect 159742 183882 159784 184118
rect 159464 183840 159784 183882
rect 200173 184118 200493 184160
rect 200173 183882 200215 184118
rect 200451 183882 200493 184118
rect 200173 183840 200493 183882
rect 144104 172918 144424 172960
rect 144104 172682 144146 172918
rect 144382 172682 144424 172918
rect 144104 172640 144424 172682
rect 197507 172918 197827 172960
rect 197507 172682 197549 172918
rect 197785 172682 197827 172918
rect 197507 172640 197827 172682
rect 226716 172918 230716 195082
rect 226716 172682 226838 172918
rect 227074 172682 227158 172918
rect 227394 172682 227478 172918
rect 227714 172682 227798 172918
rect 228034 172682 228118 172918
rect 228354 172682 228438 172918
rect 228674 172682 228758 172918
rect 228994 172682 229078 172918
rect 229314 172682 229398 172918
rect 229634 172682 229718 172918
rect 229954 172682 230038 172918
rect 230274 172682 230358 172918
rect 230594 172682 230716 172918
rect 159464 161718 159784 161760
rect 159464 161482 159506 161718
rect 159742 161482 159784 161718
rect 159464 161440 159784 161482
rect 200173 161718 200493 161760
rect 200173 161482 200215 161718
rect 200451 161482 200493 161718
rect 200173 161440 200493 161482
rect 226716 150518 230716 172682
rect 226716 150282 226838 150518
rect 227074 150282 227158 150518
rect 227394 150282 227478 150518
rect 227714 150282 227798 150518
rect 228034 150282 228118 150518
rect 228354 150282 228438 150518
rect 228674 150282 228758 150518
rect 228994 150282 229078 150518
rect 229314 150282 229398 150518
rect 229634 150282 229718 150518
rect 229954 150282 230038 150518
rect 230274 150282 230358 150518
rect 230594 150282 230716 150518
rect 150840 128118 151160 128160
rect 150840 127882 150882 128118
rect 151118 127882 151160 128118
rect 150840 127840 151160 127882
rect 193507 128118 193827 128160
rect 193507 127882 193549 128118
rect 193785 127882 193827 128118
rect 193507 127840 193827 127882
rect 226716 128118 230716 150282
rect 226716 127882 226838 128118
rect 227074 127882 227158 128118
rect 227394 127882 227478 128118
rect 227714 127882 227798 128118
rect 228034 127882 228118 128118
rect 228354 127882 228438 128118
rect 228674 127882 228758 128118
rect 228994 127882 229078 128118
rect 229314 127882 229398 128118
rect 229634 127882 229718 128118
rect 229954 127882 230038 128118
rect 230274 127882 230358 128118
rect 230594 127882 230716 128118
rect 198173 116918 198493 116960
rect 198173 116682 198215 116918
rect 198451 116682 198493 116918
rect 198173 116640 198493 116682
rect 226716 105718 230716 127882
rect 226716 105482 226838 105718
rect 227074 105482 227158 105718
rect 227394 105482 227478 105718
rect 227714 105482 227798 105718
rect 228034 105482 228118 105718
rect 228354 105482 228438 105718
rect 228674 105482 228758 105718
rect 228994 105482 229078 105718
rect 229314 105482 229398 105718
rect 229634 105482 229718 105718
rect 229954 105482 230038 105718
rect 230274 105482 230358 105718
rect 230594 105482 230716 105718
rect 209779 96716 209780 96766
rect 209844 96716 209845 96766
rect 209779 96715 209845 96716
rect 159464 94518 159784 94560
rect 159464 94282 159506 94518
rect 159742 94282 159784 94518
rect 159464 94240 159784 94282
rect 200173 94518 200493 94560
rect 200173 94282 200215 94518
rect 200451 94282 200493 94518
rect 200173 94240 200493 94282
rect 144104 83318 144424 83360
rect 144104 83082 144146 83318
rect 144382 83082 144424 83318
rect 144104 83040 144424 83082
rect 197507 83318 197827 83360
rect 197507 83082 197549 83318
rect 197785 83082 197827 83318
rect 197507 83040 197827 83082
rect 226716 83318 230716 105482
rect 226716 83082 226838 83318
rect 227074 83082 227158 83318
rect 227394 83082 227478 83318
rect 227714 83082 227798 83318
rect 228034 83082 228118 83318
rect 228354 83082 228438 83318
rect 228674 83082 228758 83318
rect 228994 83082 229078 83318
rect 229314 83082 229398 83318
rect 229634 83082 229718 83318
rect 229954 83082 230038 83318
rect 230274 83082 230358 83318
rect 230594 83082 230716 83318
rect 159464 72118 159784 72160
rect 159464 71882 159506 72118
rect 159742 71882 159784 72118
rect 159464 71840 159784 71882
rect 200173 72118 200493 72160
rect 200173 71882 200215 72118
rect 200451 71882 200493 72118
rect 200173 71840 200493 71882
rect 212355 63188 212421 63189
rect 212355 63124 212356 63188
rect 212420 63124 212421 63188
rect 212355 63123 212421 63124
rect 140227 58428 140293 58429
rect 140227 58364 140228 58428
rect 140292 58364 140293 58428
rect 140227 58363 140293 58364
rect 55955 58292 56021 58293
rect 55955 58228 55956 58292
rect 56020 58228 56021 58292
rect 55955 58227 56021 58228
rect 212358 54074 212418 63123
rect 226716 60918 230716 83082
rect 226716 60682 226838 60918
rect 227074 60682 227158 60918
rect 227394 60682 227478 60918
rect 227714 60682 227798 60918
rect 228034 60682 228118 60918
rect 228354 60682 228438 60918
rect 228674 60682 228758 60918
rect 228994 60682 229078 60918
rect 229314 60682 229398 60918
rect 229634 60682 229718 60918
rect 229954 60682 230038 60918
rect 230274 60682 230358 60918
rect 230594 60682 230716 60918
rect 212358 54014 212602 54074
rect 64971 46868 65037 46869
rect 64971 46804 64972 46868
rect 65036 46804 65037 46868
rect 64971 46803 65037 46804
rect 159547 46868 159613 46869
rect 159547 46804 159548 46868
rect 159612 46804 159613 46868
rect 159547 46803 159613 46804
rect 63499 46732 63565 46733
rect 63499 46668 63500 46732
rect 63564 46668 63565 46732
rect 63499 46667 63565 46668
rect 62211 46596 62277 46597
rect 62211 46532 62212 46596
rect 62276 46532 62277 46596
rect 62211 46531 62277 46532
rect 5000 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 9000 38518
rect 5000 16118 9000 38282
rect 25507 38518 25827 38560
rect 25507 38282 25549 38518
rect 25785 38282 25827 38518
rect 25507 38240 25827 38282
rect 30173 27318 30493 27360
rect 30173 27082 30215 27318
rect 30451 27082 30493 27318
rect 30173 27040 30493 27082
rect 62214 21029 62274 46531
rect 63131 46460 63197 46461
rect 63131 46396 63132 46460
rect 63196 46396 63197 46460
rect 63131 46395 63197 46396
rect 63134 21029 63194 46395
rect 63315 46324 63381 46325
rect 63315 46260 63316 46324
rect 63380 46260 63381 46324
rect 63315 46259 63381 46260
rect 62211 21028 62277 21029
rect 62211 20964 62212 21028
rect 62276 20964 62277 21028
rect 62211 20963 62277 20964
rect 63131 21028 63197 21029
rect 63131 20964 63132 21028
rect 63196 20964 63197 21028
rect 63131 20963 63197 20964
rect 63318 20893 63378 46259
rect 63315 20892 63381 20893
rect 63315 20828 63316 20892
rect 63380 20828 63381 20892
rect 63315 20827 63381 20828
rect 63502 18309 63562 46667
rect 64787 46188 64853 46189
rect 64787 46124 64788 46188
rect 64852 46124 64853 46188
rect 64787 46123 64853 46124
rect 64790 21029 64850 46123
rect 64974 21029 65034 46803
rect 149059 46732 149125 46733
rect 149059 46668 149060 46732
rect 149124 46668 149125 46732
rect 149059 46667 149125 46668
rect 146299 46596 146365 46597
rect 146299 46532 146300 46596
rect 146364 46532 146365 46596
rect 146299 46531 146365 46532
rect 89811 46324 89877 46325
rect 89811 46260 89812 46324
rect 89876 46260 89877 46324
rect 89811 46259 89877 46260
rect 146115 46324 146181 46325
rect 146115 46260 146116 46324
rect 146180 46260 146181 46324
rect 146115 46259 146181 46260
rect 89075 46188 89141 46189
rect 89075 46124 89076 46188
rect 89140 46124 89141 46188
rect 89075 46123 89141 46124
rect 66840 38518 67160 38560
rect 66840 38282 66882 38518
rect 67118 38282 67160 38518
rect 66840 38240 67160 38282
rect 71840 27318 72160 27360
rect 71840 27082 71882 27318
rect 72118 27082 72160 27318
rect 71840 27040 72160 27082
rect 64787 21028 64853 21029
rect 64787 20964 64788 21028
rect 64852 20964 64853 21028
rect 64787 20963 64853 20964
rect 64971 21028 65037 21029
rect 64971 20964 64972 21028
rect 65036 20964 65037 21028
rect 64971 20963 65037 20964
rect 89078 20842 89138 46123
rect 89814 20162 89874 46259
rect 109507 38518 109827 38560
rect 109507 38282 109549 38518
rect 109785 38282 109827 38518
rect 109507 38240 109827 38282
rect 114173 27318 114493 27360
rect 114173 27082 114215 27318
rect 114451 27082 114493 27318
rect 114173 27040 114493 27082
rect 146118 20893 146178 46259
rect 146302 21029 146362 46531
rect 147771 46460 147837 46461
rect 147771 46396 147772 46460
rect 147836 46396 147837 46460
rect 147771 46395 147837 46396
rect 147035 46188 147101 46189
rect 147035 46124 147036 46188
rect 147100 46124 147101 46188
rect 147035 46123 147101 46124
rect 146299 21028 146365 21029
rect 146299 20964 146300 21028
rect 146364 20964 146365 21028
rect 146299 20963 146365 20964
rect 146115 20892 146181 20893
rect 146115 20828 146116 20892
rect 146180 20828 146181 20892
rect 146115 20827 146181 20828
rect 63499 18308 63565 18309
rect 63499 18244 63500 18308
rect 63564 18244 63565 18308
rect 63499 18243 63565 18244
rect 147038 17085 147098 46123
rect 147774 21029 147834 46395
rect 149062 21029 149122 46667
rect 154947 46052 155013 46053
rect 154947 45988 154948 46052
rect 155012 45988 155013 46052
rect 154947 45987 155013 45988
rect 154950 43282 155010 45987
rect 159550 43282 159610 46803
rect 173163 46324 173229 46325
rect 173163 46260 173164 46324
rect 173228 46260 173229 46324
rect 173163 46259 173229 46260
rect 150534 22202 150594 39646
rect 150840 38518 151160 38560
rect 150840 38282 150882 38518
rect 151118 38282 151160 38518
rect 150840 38240 151160 38282
rect 147771 21028 147837 21029
rect 147771 20964 147772 21028
rect 147836 20964 147837 21028
rect 147771 20963 147837 20964
rect 149059 21028 149125 21029
rect 149059 20964 149060 21028
rect 149124 20964 149125 21028
rect 149059 20963 149125 20964
rect 151638 18309 151698 40326
rect 155840 27318 156160 27360
rect 155840 27082 155882 27318
rect 156118 27082 156160 27318
rect 155840 27040 156160 27082
rect 156054 21029 156114 21966
rect 156051 21028 156117 21029
rect 156051 20964 156052 21028
rect 156116 20964 156117 21028
rect 156051 20963 156117 20964
rect 173166 20842 173226 46259
rect 173531 46188 173597 46189
rect 173531 46124 173532 46188
rect 173596 46124 173597 46188
rect 173531 46123 173597 46124
rect 173534 20162 173594 46123
rect 173899 44692 173965 44693
rect 173899 44628 173900 44692
rect 173964 44628 173965 44692
rect 173899 44627 173965 44628
rect 173902 22202 173962 44627
rect 212542 44554 212602 54014
rect 212542 44494 212786 44554
rect 193507 38518 193827 38560
rect 193507 38282 193549 38518
rect 193785 38282 193827 38518
rect 193507 38240 193827 38282
rect 212726 35802 212786 44494
rect 226716 38518 230716 60682
rect 226716 38282 226838 38518
rect 227074 38282 227158 38518
rect 227394 38282 227478 38518
rect 227714 38282 227798 38518
rect 228034 38282 228118 38518
rect 228354 38282 228438 38518
rect 228674 38282 228758 38518
rect 228994 38282 229078 38518
rect 229314 38282 229398 38518
rect 229634 38282 229718 38518
rect 229954 38282 230038 38518
rect 230274 38282 230358 38518
rect 230594 38282 230716 38518
rect 198173 27318 198493 27360
rect 198173 27082 198215 27318
rect 198451 27082 198493 27318
rect 198173 27040 198493 27082
rect 212726 25602 212786 34886
rect 185123 21916 185124 21966
rect 185188 21916 185189 21966
rect 185123 21915 185189 21916
rect 212726 21522 212786 24686
rect 222291 21980 222357 21981
rect 222291 21916 222292 21980
rect 222356 21916 222357 21980
rect 222291 21915 222357 21916
rect 222294 21522 222354 21915
rect 185491 20892 185557 20893
rect 185491 20828 185492 20892
rect 185556 20828 185557 20892
rect 185491 20827 185557 20828
rect 185494 20162 185554 20827
rect 212726 20754 212786 21286
rect 212542 20694 212786 20754
rect 212542 18445 212602 20694
rect 212539 18444 212605 18445
rect 212539 18380 212540 18444
rect 212604 18380 212605 18444
rect 212539 18379 212605 18380
rect 151635 18308 151701 18309
rect 151635 18244 151636 18308
rect 151700 18244 151701 18308
rect 151635 18243 151701 18244
rect 147035 17084 147101 17085
rect 147035 17020 147036 17084
rect 147100 17020 147101 17084
rect 147035 17019 147101 17020
rect 5000 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 9000 16118
rect 5000 8878 9000 15882
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 226716 16118 230716 38282
rect 226716 15882 226838 16118
rect 227074 15882 227158 16118
rect 227394 15882 227478 16118
rect 227714 15882 227798 16118
rect 228034 15882 228118 16118
rect 228354 15882 228438 16118
rect 228674 15882 228758 16118
rect 228994 15882 229078 16118
rect 229314 15882 229398 16118
rect 229634 15882 229718 16118
rect 229954 15882 230038 16118
rect 230274 15882 230358 16118
rect 230594 15882 230716 16118
rect 226716 8878 230716 15882
rect 226716 8642 226838 8878
rect 227074 8642 227158 8878
rect 227394 8642 227478 8878
rect 227714 8642 227798 8878
rect 228034 8642 228118 8878
rect 228354 8642 228438 8878
rect 228674 8642 228758 8878
rect 228994 8642 229078 8878
rect 229314 8642 229398 8878
rect 229634 8642 229718 8878
rect 229954 8642 230038 8878
rect 230274 8642 230358 8878
rect 230594 8642 230716 8878
rect 226716 8558 230716 8642
rect 226716 8322 226838 8558
rect 227074 8322 227158 8558
rect 227394 8322 227478 8558
rect 227714 8322 227798 8558
rect 228034 8322 228118 8558
rect 228354 8322 228438 8558
rect 228674 8322 228758 8558
rect 228994 8322 229078 8558
rect 229314 8322 229398 8558
rect 229634 8322 229718 8558
rect 229954 8322 230038 8558
rect 230274 8322 230358 8558
rect 230594 8322 230716 8558
rect 226716 8238 230716 8322
rect 226716 8002 226838 8238
rect 227074 8002 227158 8238
rect 227394 8002 227478 8238
rect 227714 8002 227798 8238
rect 228034 8002 228118 8238
rect 228354 8002 228438 8238
rect 228674 8002 228758 8238
rect 228994 8002 229078 8238
rect 229314 8002 229398 8238
rect 229634 8002 229718 8238
rect 229954 8002 230038 8238
rect 230274 8002 230358 8238
rect 230594 8002 230716 8238
rect 226716 7918 230716 8002
rect 226716 7682 226838 7918
rect 227074 7682 227158 7918
rect 227394 7682 227478 7918
rect 227714 7682 227798 7918
rect 228034 7682 228118 7918
rect 228354 7682 228438 7918
rect 228674 7682 228758 7918
rect 228994 7682 229078 7918
rect 229314 7682 229398 7918
rect 229634 7682 229718 7918
rect 229954 7682 230038 7918
rect 230274 7682 230358 7918
rect 230594 7682 230716 7918
rect 226716 7598 230716 7682
rect 226716 7362 226838 7598
rect 227074 7362 227158 7598
rect 227394 7362 227478 7598
rect 227714 7362 227798 7598
rect 228034 7362 228118 7598
rect 228354 7362 228438 7598
rect 228674 7362 228758 7598
rect 228994 7362 229078 7598
rect 229314 7362 229398 7598
rect 229634 7362 229718 7598
rect 229954 7362 230038 7598
rect 230274 7362 230358 7598
rect 230594 7362 230716 7598
rect 226716 7278 230716 7362
rect 226716 7042 226838 7278
rect 227074 7042 227158 7278
rect 227394 7042 227478 7278
rect 227714 7042 227798 7278
rect 228034 7042 228118 7278
rect 228354 7042 228438 7278
rect 228674 7042 228758 7278
rect 228994 7042 229078 7278
rect 229314 7042 229398 7278
rect 229634 7042 229718 7278
rect 229954 7042 230038 7278
rect 230274 7042 230358 7278
rect 230594 7042 230716 7278
rect 226716 6958 230716 7042
rect 226716 6722 226838 6958
rect 227074 6722 227158 6958
rect 227394 6722 227478 6958
rect 227714 6722 227798 6958
rect 228034 6722 228118 6958
rect 228354 6722 228438 6958
rect 228674 6722 228758 6958
rect 228994 6722 229078 6958
rect 229314 6722 229398 6958
rect 229634 6722 229718 6958
rect 229954 6722 230038 6958
rect 230274 6722 230358 6958
rect 230594 6722 230716 6958
rect 226716 6638 230716 6722
rect 226716 6402 226838 6638
rect 227074 6402 227158 6638
rect 227394 6402 227478 6638
rect 227714 6402 227798 6638
rect 228034 6402 228118 6638
rect 228354 6402 228438 6638
rect 228674 6402 228758 6638
rect 228994 6402 229078 6638
rect 229314 6402 229398 6638
rect 229634 6402 229718 6638
rect 229954 6402 230038 6638
rect 230274 6402 230358 6638
rect 230594 6402 230716 6638
rect 226716 6318 230716 6402
rect 226716 6082 226838 6318
rect 227074 6082 227158 6318
rect 227394 6082 227478 6318
rect 227714 6082 227798 6318
rect 228034 6082 228118 6318
rect 228354 6082 228438 6318
rect 228674 6082 228758 6318
rect 228994 6082 229078 6318
rect 229314 6082 229398 6318
rect 229634 6082 229718 6318
rect 229954 6082 230038 6318
rect 230274 6082 230358 6318
rect 230594 6082 230716 6318
rect 226716 5998 230716 6082
rect 226716 5762 226838 5998
rect 227074 5762 227158 5998
rect 227394 5762 227478 5998
rect 227714 5762 227798 5998
rect 228034 5762 228118 5998
rect 228354 5762 228438 5998
rect 228674 5762 228758 5998
rect 228994 5762 229078 5998
rect 229314 5762 229398 5998
rect 229634 5762 229718 5998
rect 229954 5762 230038 5998
rect 230274 5762 230358 5998
rect 230594 5762 230716 5998
rect 226716 5678 230716 5762
rect 226716 5442 226838 5678
rect 227074 5442 227158 5678
rect 227394 5442 227478 5678
rect 227714 5442 227798 5678
rect 228034 5442 228118 5678
rect 228354 5442 228438 5678
rect 228674 5442 228758 5678
rect 228994 5442 229078 5678
rect 229314 5442 229398 5678
rect 229634 5442 229718 5678
rect 229954 5442 230038 5678
rect 230274 5442 230358 5678
rect 230594 5442 230716 5678
rect 226716 5358 230716 5442
rect 226716 5122 226838 5358
rect 227074 5122 227158 5358
rect 227394 5122 227478 5358
rect 227714 5122 227798 5358
rect 228034 5122 228118 5358
rect 228354 5122 228438 5358
rect 228674 5122 228758 5358
rect 228994 5122 229078 5358
rect 229314 5122 229398 5358
rect 229634 5122 229718 5358
rect 229954 5122 230038 5358
rect 230274 5122 230358 5358
rect 230594 5122 230716 5358
rect 226716 5000 230716 5122
rect 231716 228918 235716 249322
rect 231716 228682 231838 228918
rect 232074 228682 232158 228918
rect 232394 228682 232478 228918
rect 232714 228682 232798 228918
rect 233034 228682 233118 228918
rect 233354 228682 233438 228918
rect 233674 228682 233758 228918
rect 233994 228682 234078 228918
rect 234314 228682 234398 228918
rect 234634 228682 234718 228918
rect 234954 228682 235038 228918
rect 235274 228682 235358 228918
rect 235594 228682 235716 228918
rect 231716 206518 235716 228682
rect 231716 206282 231838 206518
rect 232074 206282 232158 206518
rect 232394 206282 232478 206518
rect 232714 206282 232798 206518
rect 233034 206282 233118 206518
rect 233354 206282 233438 206518
rect 233674 206282 233758 206518
rect 233994 206282 234078 206518
rect 234314 206282 234398 206518
rect 234634 206282 234718 206518
rect 234954 206282 235038 206518
rect 235274 206282 235358 206518
rect 235594 206282 235716 206518
rect 231716 184118 235716 206282
rect 231716 183882 231838 184118
rect 232074 183882 232158 184118
rect 232394 183882 232478 184118
rect 232714 183882 232798 184118
rect 233034 183882 233118 184118
rect 233354 183882 233438 184118
rect 233674 183882 233758 184118
rect 233994 183882 234078 184118
rect 234314 183882 234398 184118
rect 234634 183882 234718 184118
rect 234954 183882 235038 184118
rect 235274 183882 235358 184118
rect 235594 183882 235716 184118
rect 231716 161718 235716 183882
rect 231716 161482 231838 161718
rect 232074 161482 232158 161718
rect 232394 161482 232478 161718
rect 232714 161482 232798 161718
rect 233034 161482 233118 161718
rect 233354 161482 233438 161718
rect 233674 161482 233758 161718
rect 233994 161482 234078 161718
rect 234314 161482 234398 161718
rect 234634 161482 234718 161718
rect 234954 161482 235038 161718
rect 235274 161482 235358 161718
rect 235594 161482 235716 161718
rect 231716 139318 235716 161482
rect 231716 139082 231838 139318
rect 232074 139082 232158 139318
rect 232394 139082 232478 139318
rect 232714 139082 232798 139318
rect 233034 139082 233118 139318
rect 233354 139082 233438 139318
rect 233674 139082 233758 139318
rect 233994 139082 234078 139318
rect 234314 139082 234398 139318
rect 234634 139082 234718 139318
rect 234954 139082 235038 139318
rect 235274 139082 235358 139318
rect 235594 139082 235716 139318
rect 231716 116918 235716 139082
rect 231716 116682 231838 116918
rect 232074 116682 232158 116918
rect 232394 116682 232478 116918
rect 232714 116682 232798 116918
rect 233034 116682 233118 116918
rect 233354 116682 233438 116918
rect 233674 116682 233758 116918
rect 233994 116682 234078 116918
rect 234314 116682 234398 116918
rect 234634 116682 234718 116918
rect 234954 116682 235038 116918
rect 235274 116682 235358 116918
rect 235594 116682 235716 116918
rect 231716 94518 235716 116682
rect 231716 94282 231838 94518
rect 232074 94282 232158 94518
rect 232394 94282 232478 94518
rect 232714 94282 232798 94518
rect 233034 94282 233118 94518
rect 233354 94282 233438 94518
rect 233674 94282 233758 94518
rect 233994 94282 234078 94518
rect 234314 94282 234398 94518
rect 234634 94282 234718 94518
rect 234954 94282 235038 94518
rect 235274 94282 235358 94518
rect 235594 94282 235716 94518
rect 231716 72118 235716 94282
rect 231716 71882 231838 72118
rect 232074 71882 232158 72118
rect 232394 71882 232478 72118
rect 232714 71882 232798 72118
rect 233034 71882 233118 72118
rect 233354 71882 233438 72118
rect 233674 71882 233758 72118
rect 233994 71882 234078 72118
rect 234314 71882 234398 72118
rect 234634 71882 234718 72118
rect 234954 71882 235038 72118
rect 235274 71882 235358 72118
rect 235594 71882 235716 72118
rect 231716 49718 235716 71882
rect 231716 49482 231838 49718
rect 232074 49482 232158 49718
rect 232394 49482 232478 49718
rect 232714 49482 232798 49718
rect 233034 49482 233118 49718
rect 233354 49482 233438 49718
rect 233674 49482 233758 49718
rect 233994 49482 234078 49718
rect 234314 49482 234398 49718
rect 234634 49482 234718 49718
rect 234954 49482 235038 49718
rect 235274 49482 235358 49718
rect 235594 49482 235716 49718
rect 231716 27318 235716 49482
rect 231716 27082 231838 27318
rect 232074 27082 232158 27318
rect 232394 27082 232478 27318
rect 232714 27082 232798 27318
rect 233034 27082 233118 27318
rect 233354 27082 233438 27318
rect 233674 27082 233758 27318
rect 233994 27082 234078 27318
rect 234314 27082 234398 27318
rect 234634 27082 234718 27318
rect 234954 27082 235038 27318
rect 235274 27082 235358 27318
rect 235594 27082 235716 27318
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 231716 3878 235716 27082
rect 231716 3642 231838 3878
rect 232074 3642 232158 3878
rect 232394 3642 232478 3878
rect 232714 3642 232798 3878
rect 233034 3642 233118 3878
rect 233354 3642 233438 3878
rect 233674 3642 233758 3878
rect 233994 3642 234078 3878
rect 234314 3642 234398 3878
rect 234634 3642 234718 3878
rect 234954 3642 235038 3878
rect 235274 3642 235358 3878
rect 235594 3642 235716 3878
rect 231716 3558 235716 3642
rect 231716 3322 231838 3558
rect 232074 3322 232158 3558
rect 232394 3322 232478 3558
rect 232714 3322 232798 3558
rect 233034 3322 233118 3558
rect 233354 3322 233438 3558
rect 233674 3322 233758 3558
rect 233994 3322 234078 3558
rect 234314 3322 234398 3558
rect 234634 3322 234718 3558
rect 234954 3322 235038 3558
rect 235274 3322 235358 3558
rect 235594 3322 235716 3558
rect 231716 3238 235716 3322
rect 231716 3002 231838 3238
rect 232074 3002 232158 3238
rect 232394 3002 232478 3238
rect 232714 3002 232798 3238
rect 233034 3002 233118 3238
rect 233354 3002 233438 3238
rect 233674 3002 233758 3238
rect 233994 3002 234078 3238
rect 234314 3002 234398 3238
rect 234634 3002 234718 3238
rect 234954 3002 235038 3238
rect 235274 3002 235358 3238
rect 235594 3002 235716 3238
rect 231716 2918 235716 3002
rect 231716 2682 231838 2918
rect 232074 2682 232158 2918
rect 232394 2682 232478 2918
rect 232714 2682 232798 2918
rect 233034 2682 233118 2918
rect 233354 2682 233438 2918
rect 233674 2682 233758 2918
rect 233994 2682 234078 2918
rect 234314 2682 234398 2918
rect 234634 2682 234718 2918
rect 234954 2682 235038 2918
rect 235274 2682 235358 2918
rect 235594 2682 235716 2918
rect 231716 2598 235716 2682
rect 231716 2362 231838 2598
rect 232074 2362 232158 2598
rect 232394 2362 232478 2598
rect 232714 2362 232798 2598
rect 233034 2362 233118 2598
rect 233354 2362 233438 2598
rect 233674 2362 233758 2598
rect 233994 2362 234078 2598
rect 234314 2362 234398 2598
rect 234634 2362 234718 2598
rect 234954 2362 235038 2598
rect 235274 2362 235358 2598
rect 235594 2362 235716 2598
rect 231716 2278 235716 2362
rect 231716 2042 231838 2278
rect 232074 2042 232158 2278
rect 232394 2042 232478 2278
rect 232714 2042 232798 2278
rect 233034 2042 233118 2278
rect 233354 2042 233438 2278
rect 233674 2042 233758 2278
rect 233994 2042 234078 2278
rect 234314 2042 234398 2278
rect 234634 2042 234718 2278
rect 234954 2042 235038 2278
rect 235274 2042 235358 2278
rect 235594 2042 235716 2278
rect 231716 1958 235716 2042
rect 231716 1722 231838 1958
rect 232074 1722 232158 1958
rect 232394 1722 232478 1958
rect 232714 1722 232798 1958
rect 233034 1722 233118 1958
rect 233354 1722 233438 1958
rect 233674 1722 233758 1958
rect 233994 1722 234078 1958
rect 234314 1722 234398 1958
rect 234634 1722 234718 1958
rect 234954 1722 235038 1958
rect 235274 1722 235358 1958
rect 235594 1722 235716 1958
rect 231716 1638 235716 1722
rect 231716 1402 231838 1638
rect 232074 1402 232158 1638
rect 232394 1402 232478 1638
rect 232714 1402 232798 1638
rect 233034 1402 233118 1638
rect 233354 1402 233438 1638
rect 233674 1402 233758 1638
rect 233994 1402 234078 1638
rect 234314 1402 234398 1638
rect 234634 1402 234718 1638
rect 234954 1402 235038 1638
rect 235274 1402 235358 1638
rect 235594 1402 235716 1638
rect 231716 1318 235716 1402
rect 231716 1082 231838 1318
rect 232074 1082 232158 1318
rect 232394 1082 232478 1318
rect 232714 1082 232798 1318
rect 233034 1082 233118 1318
rect 233354 1082 233438 1318
rect 233674 1082 233758 1318
rect 233994 1082 234078 1318
rect 234314 1082 234398 1318
rect 234634 1082 234718 1318
rect 234954 1082 235038 1318
rect 235274 1082 235358 1318
rect 235594 1082 235716 1318
rect 231716 998 235716 1082
rect 231716 762 231838 998
rect 232074 762 232158 998
rect 232394 762 232478 998
rect 232714 762 232798 998
rect 233034 762 233118 998
rect 233354 762 233438 998
rect 233674 762 233758 998
rect 233994 762 234078 998
rect 234314 762 234398 998
rect 234634 762 234718 998
rect 234954 762 235038 998
rect 235274 762 235358 998
rect 235594 762 235716 998
rect 231716 678 235716 762
rect 231716 442 231838 678
rect 232074 442 232158 678
rect 232394 442 232478 678
rect 232714 442 232798 678
rect 233034 442 233118 678
rect 233354 442 233438 678
rect 233674 442 233758 678
rect 233994 442 234078 678
rect 234314 442 234398 678
rect 234634 442 234718 678
rect 234954 442 235038 678
rect 235274 442 235358 678
rect 235594 442 235716 678
rect 231716 358 235716 442
rect 231716 122 231838 358
rect 232074 122 232158 358
rect 232394 122 232478 358
rect 232714 122 232798 358
rect 233034 122 233118 358
rect 233354 122 233438 358
rect 233674 122 233758 358
rect 233994 122 234078 358
rect 234314 122 234398 358
rect 234634 122 234718 358
rect 234954 122 235038 358
rect 235274 122 235358 358
rect 235594 122 235716 358
rect 231716 0 235716 122
<< via4 >>
rect 122 252842 358 253078
rect 442 252842 678 253078
rect 762 252842 998 253078
rect 1082 252842 1318 253078
rect 1402 252842 1638 253078
rect 1722 252842 1958 253078
rect 2042 252842 2278 253078
rect 2362 252842 2598 253078
rect 2682 252842 2918 253078
rect 3002 252842 3238 253078
rect 3322 252842 3558 253078
rect 3642 252842 3878 253078
rect 122 252522 358 252758
rect 442 252522 678 252758
rect 762 252522 998 252758
rect 1082 252522 1318 252758
rect 1402 252522 1638 252758
rect 1722 252522 1958 252758
rect 2042 252522 2278 252758
rect 2362 252522 2598 252758
rect 2682 252522 2918 252758
rect 3002 252522 3238 252758
rect 3322 252522 3558 252758
rect 3642 252522 3878 252758
rect 122 252202 358 252438
rect 442 252202 678 252438
rect 762 252202 998 252438
rect 1082 252202 1318 252438
rect 1402 252202 1638 252438
rect 1722 252202 1958 252438
rect 2042 252202 2278 252438
rect 2362 252202 2598 252438
rect 2682 252202 2918 252438
rect 3002 252202 3238 252438
rect 3322 252202 3558 252438
rect 3642 252202 3878 252438
rect 122 251882 358 252118
rect 442 251882 678 252118
rect 762 251882 998 252118
rect 1082 251882 1318 252118
rect 1402 251882 1638 252118
rect 1722 251882 1958 252118
rect 2042 251882 2278 252118
rect 2362 251882 2598 252118
rect 2682 251882 2918 252118
rect 3002 251882 3238 252118
rect 3322 251882 3558 252118
rect 3642 251882 3878 252118
rect 122 251562 358 251798
rect 442 251562 678 251798
rect 762 251562 998 251798
rect 1082 251562 1318 251798
rect 1402 251562 1638 251798
rect 1722 251562 1958 251798
rect 2042 251562 2278 251798
rect 2362 251562 2598 251798
rect 2682 251562 2918 251798
rect 3002 251562 3238 251798
rect 3322 251562 3558 251798
rect 3642 251562 3878 251798
rect 122 251242 358 251478
rect 442 251242 678 251478
rect 762 251242 998 251478
rect 1082 251242 1318 251478
rect 1402 251242 1638 251478
rect 1722 251242 1958 251478
rect 2042 251242 2278 251478
rect 2362 251242 2598 251478
rect 2682 251242 2918 251478
rect 3002 251242 3238 251478
rect 3322 251242 3558 251478
rect 3642 251242 3878 251478
rect 122 250922 358 251158
rect 442 250922 678 251158
rect 762 250922 998 251158
rect 1082 250922 1318 251158
rect 1402 250922 1638 251158
rect 1722 250922 1958 251158
rect 2042 250922 2278 251158
rect 2362 250922 2598 251158
rect 2682 250922 2918 251158
rect 3002 250922 3238 251158
rect 3322 250922 3558 251158
rect 3642 250922 3878 251158
rect 122 250602 358 250838
rect 442 250602 678 250838
rect 762 250602 998 250838
rect 1082 250602 1318 250838
rect 1402 250602 1638 250838
rect 1722 250602 1958 250838
rect 2042 250602 2278 250838
rect 2362 250602 2598 250838
rect 2682 250602 2918 250838
rect 3002 250602 3238 250838
rect 3322 250602 3558 250838
rect 3642 250602 3878 250838
rect 122 250282 358 250518
rect 442 250282 678 250518
rect 762 250282 998 250518
rect 1082 250282 1318 250518
rect 1402 250282 1638 250518
rect 1722 250282 1958 250518
rect 2042 250282 2278 250518
rect 2362 250282 2598 250518
rect 2682 250282 2918 250518
rect 3002 250282 3238 250518
rect 3322 250282 3558 250518
rect 3642 250282 3878 250518
rect 122 249962 358 250198
rect 442 249962 678 250198
rect 762 249962 998 250198
rect 1082 249962 1318 250198
rect 1402 249962 1638 250198
rect 1722 249962 1958 250198
rect 2042 249962 2278 250198
rect 2362 249962 2598 250198
rect 2682 249962 2918 250198
rect 3002 249962 3238 250198
rect 3322 249962 3558 250198
rect 3642 249962 3878 250198
rect 122 249642 358 249878
rect 442 249642 678 249878
rect 762 249642 998 249878
rect 1082 249642 1318 249878
rect 1402 249642 1638 249878
rect 1722 249642 1958 249878
rect 2042 249642 2278 249878
rect 2362 249642 2598 249878
rect 2682 249642 2918 249878
rect 3002 249642 3238 249878
rect 3322 249642 3558 249878
rect 3642 249642 3878 249878
rect 122 249322 358 249558
rect 442 249322 678 249558
rect 762 249322 998 249558
rect 1082 249322 1318 249558
rect 1402 249322 1638 249558
rect 1722 249322 1958 249558
rect 2042 249322 2278 249558
rect 2362 249322 2598 249558
rect 2682 249322 2918 249558
rect 3002 249322 3238 249558
rect 3322 249322 3558 249558
rect 3642 249322 3878 249558
rect 231838 252842 232074 253078
rect 232158 252842 232394 253078
rect 232478 252842 232714 253078
rect 232798 252842 233034 253078
rect 233118 252842 233354 253078
rect 233438 252842 233674 253078
rect 233758 252842 233994 253078
rect 234078 252842 234314 253078
rect 234398 252842 234634 253078
rect 234718 252842 234954 253078
rect 235038 252842 235274 253078
rect 235358 252842 235594 253078
rect 231838 252522 232074 252758
rect 232158 252522 232394 252758
rect 232478 252522 232714 252758
rect 232798 252522 233034 252758
rect 233118 252522 233354 252758
rect 233438 252522 233674 252758
rect 233758 252522 233994 252758
rect 234078 252522 234314 252758
rect 234398 252522 234634 252758
rect 234718 252522 234954 252758
rect 235038 252522 235274 252758
rect 235358 252522 235594 252758
rect 231838 252202 232074 252438
rect 232158 252202 232394 252438
rect 232478 252202 232714 252438
rect 232798 252202 233034 252438
rect 233118 252202 233354 252438
rect 233438 252202 233674 252438
rect 233758 252202 233994 252438
rect 234078 252202 234314 252438
rect 234398 252202 234634 252438
rect 234718 252202 234954 252438
rect 235038 252202 235274 252438
rect 235358 252202 235594 252438
rect 231838 251882 232074 252118
rect 232158 251882 232394 252118
rect 232478 251882 232714 252118
rect 232798 251882 233034 252118
rect 233118 251882 233354 252118
rect 233438 251882 233674 252118
rect 233758 251882 233994 252118
rect 234078 251882 234314 252118
rect 234398 251882 234634 252118
rect 234718 251882 234954 252118
rect 235038 251882 235274 252118
rect 235358 251882 235594 252118
rect 231838 251562 232074 251798
rect 232158 251562 232394 251798
rect 232478 251562 232714 251798
rect 232798 251562 233034 251798
rect 233118 251562 233354 251798
rect 233438 251562 233674 251798
rect 233758 251562 233994 251798
rect 234078 251562 234314 251798
rect 234398 251562 234634 251798
rect 234718 251562 234954 251798
rect 235038 251562 235274 251798
rect 235358 251562 235594 251798
rect 231838 251242 232074 251478
rect 232158 251242 232394 251478
rect 232478 251242 232714 251478
rect 232798 251242 233034 251478
rect 233118 251242 233354 251478
rect 233438 251242 233674 251478
rect 233758 251242 233994 251478
rect 234078 251242 234314 251478
rect 234398 251242 234634 251478
rect 234718 251242 234954 251478
rect 235038 251242 235274 251478
rect 235358 251242 235594 251478
rect 231838 250922 232074 251158
rect 232158 250922 232394 251158
rect 232478 250922 232714 251158
rect 232798 250922 233034 251158
rect 233118 250922 233354 251158
rect 233438 250922 233674 251158
rect 233758 250922 233994 251158
rect 234078 250922 234314 251158
rect 234398 250922 234634 251158
rect 234718 250922 234954 251158
rect 235038 250922 235274 251158
rect 235358 250922 235594 251158
rect 231838 250602 232074 250838
rect 232158 250602 232394 250838
rect 232478 250602 232714 250838
rect 232798 250602 233034 250838
rect 233118 250602 233354 250838
rect 233438 250602 233674 250838
rect 233758 250602 233994 250838
rect 234078 250602 234314 250838
rect 234398 250602 234634 250838
rect 234718 250602 234954 250838
rect 235038 250602 235274 250838
rect 235358 250602 235594 250838
rect 231838 250282 232074 250518
rect 232158 250282 232394 250518
rect 232478 250282 232714 250518
rect 232798 250282 233034 250518
rect 233118 250282 233354 250518
rect 233438 250282 233674 250518
rect 233758 250282 233994 250518
rect 234078 250282 234314 250518
rect 234398 250282 234634 250518
rect 234718 250282 234954 250518
rect 235038 250282 235274 250518
rect 235358 250282 235594 250518
rect 231838 249962 232074 250198
rect 232158 249962 232394 250198
rect 232478 249962 232714 250198
rect 232798 249962 233034 250198
rect 233118 249962 233354 250198
rect 233438 249962 233674 250198
rect 233758 249962 233994 250198
rect 234078 249962 234314 250198
rect 234398 249962 234634 250198
rect 234718 249962 234954 250198
rect 235038 249962 235274 250198
rect 235358 249962 235594 250198
rect 231838 249642 232074 249878
rect 232158 249642 232394 249878
rect 232478 249642 232714 249878
rect 232798 249642 233034 249878
rect 233118 249642 233354 249878
rect 233438 249642 233674 249878
rect 233758 249642 233994 249878
rect 234078 249642 234314 249878
rect 234398 249642 234634 249878
rect 234718 249642 234954 249878
rect 235038 249642 235274 249878
rect 235358 249642 235594 249878
rect 231838 249322 232074 249558
rect 232158 249322 232394 249558
rect 232478 249322 232714 249558
rect 232798 249322 233034 249558
rect 233118 249322 233354 249558
rect 233438 249322 233674 249558
rect 233758 249322 233994 249558
rect 234078 249322 234314 249558
rect 234398 249322 234634 249558
rect 234718 249322 234954 249558
rect 235038 249322 235274 249558
rect 235358 249322 235594 249558
rect 122 228682 358 228918
rect 442 228682 678 228918
rect 762 228682 998 228918
rect 1082 228682 1318 228918
rect 1402 228682 1638 228918
rect 1722 228682 1958 228918
rect 2042 228682 2278 228918
rect 2362 228682 2598 228918
rect 2682 228682 2918 228918
rect 3002 228682 3238 228918
rect 3322 228682 3558 228918
rect 3642 228682 3878 228918
rect 122 206282 358 206518
rect 442 206282 678 206518
rect 762 206282 998 206518
rect 1082 206282 1318 206518
rect 1402 206282 1638 206518
rect 1722 206282 1958 206518
rect 2042 206282 2278 206518
rect 2362 206282 2598 206518
rect 2682 206282 2918 206518
rect 3002 206282 3238 206518
rect 3322 206282 3558 206518
rect 3642 206282 3878 206518
rect 122 183882 358 184118
rect 442 183882 678 184118
rect 762 183882 998 184118
rect 1082 183882 1318 184118
rect 1402 183882 1638 184118
rect 1722 183882 1958 184118
rect 2042 183882 2278 184118
rect 2362 183882 2598 184118
rect 2682 183882 2918 184118
rect 3002 183882 3238 184118
rect 3322 183882 3558 184118
rect 3642 183882 3878 184118
rect 122 161482 358 161718
rect 442 161482 678 161718
rect 762 161482 998 161718
rect 1082 161482 1318 161718
rect 1402 161482 1638 161718
rect 1722 161482 1958 161718
rect 2042 161482 2278 161718
rect 2362 161482 2598 161718
rect 2682 161482 2918 161718
rect 3002 161482 3238 161718
rect 3322 161482 3558 161718
rect 3642 161482 3878 161718
rect 122 139082 358 139318
rect 442 139082 678 139318
rect 762 139082 998 139318
rect 1082 139082 1318 139318
rect 1402 139082 1638 139318
rect 1722 139082 1958 139318
rect 2042 139082 2278 139318
rect 2362 139082 2598 139318
rect 2682 139082 2918 139318
rect 3002 139082 3238 139318
rect 3322 139082 3558 139318
rect 3642 139082 3878 139318
rect 122 116682 358 116918
rect 442 116682 678 116918
rect 762 116682 998 116918
rect 1082 116682 1318 116918
rect 1402 116682 1638 116918
rect 1722 116682 1958 116918
rect 2042 116682 2278 116918
rect 2362 116682 2598 116918
rect 2682 116682 2918 116918
rect 3002 116682 3238 116918
rect 3322 116682 3558 116918
rect 3642 116682 3878 116918
rect 122 94282 358 94518
rect 442 94282 678 94518
rect 762 94282 998 94518
rect 1082 94282 1318 94518
rect 1402 94282 1638 94518
rect 1722 94282 1958 94518
rect 2042 94282 2278 94518
rect 2362 94282 2598 94518
rect 2682 94282 2918 94518
rect 3002 94282 3238 94518
rect 3322 94282 3558 94518
rect 3642 94282 3878 94518
rect 122 71882 358 72118
rect 442 71882 678 72118
rect 762 71882 998 72118
rect 1082 71882 1318 72118
rect 1402 71882 1638 72118
rect 1722 71882 1958 72118
rect 2042 71882 2278 72118
rect 2362 71882 2598 72118
rect 2682 71882 2918 72118
rect 3002 71882 3238 72118
rect 3322 71882 3558 72118
rect 3642 71882 3878 72118
rect 122 49482 358 49718
rect 442 49482 678 49718
rect 762 49482 998 49718
rect 1082 49482 1318 49718
rect 1402 49482 1638 49718
rect 1722 49482 1958 49718
rect 2042 49482 2278 49718
rect 2362 49482 2598 49718
rect 2682 49482 2918 49718
rect 3002 49482 3238 49718
rect 3322 49482 3558 49718
rect 3642 49482 3878 49718
rect 122 27082 358 27318
rect 442 27082 678 27318
rect 762 27082 998 27318
rect 1082 27082 1318 27318
rect 1402 27082 1638 27318
rect 1722 27082 1958 27318
rect 2042 27082 2278 27318
rect 2362 27082 2598 27318
rect 2682 27082 2918 27318
rect 3002 27082 3238 27318
rect 3322 27082 3558 27318
rect 3642 27082 3878 27318
rect 5122 247842 5358 248078
rect 5442 247842 5678 248078
rect 5762 247842 5998 248078
rect 6082 247842 6318 248078
rect 6402 247842 6638 248078
rect 6722 247842 6958 248078
rect 7042 247842 7278 248078
rect 7362 247842 7598 248078
rect 7682 247842 7918 248078
rect 8002 247842 8238 248078
rect 8322 247842 8558 248078
rect 8642 247842 8878 248078
rect 5122 247522 5358 247758
rect 5442 247522 5678 247758
rect 5762 247522 5998 247758
rect 6082 247522 6318 247758
rect 6402 247522 6638 247758
rect 6722 247522 6958 247758
rect 7042 247522 7278 247758
rect 7362 247522 7598 247758
rect 7682 247522 7918 247758
rect 8002 247522 8238 247758
rect 8322 247522 8558 247758
rect 8642 247522 8878 247758
rect 5122 247202 5358 247438
rect 5442 247202 5678 247438
rect 5762 247202 5998 247438
rect 6082 247202 6318 247438
rect 6402 247202 6638 247438
rect 6722 247202 6958 247438
rect 7042 247202 7278 247438
rect 7362 247202 7598 247438
rect 7682 247202 7918 247438
rect 8002 247202 8238 247438
rect 8322 247202 8558 247438
rect 8642 247202 8878 247438
rect 5122 246882 5358 247118
rect 5442 246882 5678 247118
rect 5762 246882 5998 247118
rect 6082 246882 6318 247118
rect 6402 246882 6638 247118
rect 6722 246882 6958 247118
rect 7042 246882 7278 247118
rect 7362 246882 7598 247118
rect 7682 246882 7918 247118
rect 8002 246882 8238 247118
rect 8322 246882 8558 247118
rect 8642 246882 8878 247118
rect 5122 246562 5358 246798
rect 5442 246562 5678 246798
rect 5762 246562 5998 246798
rect 6082 246562 6318 246798
rect 6402 246562 6638 246798
rect 6722 246562 6958 246798
rect 7042 246562 7278 246798
rect 7362 246562 7598 246798
rect 7682 246562 7918 246798
rect 8002 246562 8238 246798
rect 8322 246562 8558 246798
rect 8642 246562 8878 246798
rect 5122 246242 5358 246478
rect 5442 246242 5678 246478
rect 5762 246242 5998 246478
rect 6082 246242 6318 246478
rect 6402 246242 6638 246478
rect 6722 246242 6958 246478
rect 7042 246242 7278 246478
rect 7362 246242 7598 246478
rect 7682 246242 7918 246478
rect 8002 246242 8238 246478
rect 8322 246242 8558 246478
rect 8642 246242 8878 246478
rect 5122 245922 5358 246158
rect 5442 245922 5678 246158
rect 5762 245922 5998 246158
rect 6082 245922 6318 246158
rect 6402 245922 6638 246158
rect 6722 245922 6958 246158
rect 7042 245922 7278 246158
rect 7362 245922 7598 246158
rect 7682 245922 7918 246158
rect 8002 245922 8238 246158
rect 8322 245922 8558 246158
rect 8642 245922 8878 246158
rect 5122 245602 5358 245838
rect 5442 245602 5678 245838
rect 5762 245602 5998 245838
rect 6082 245602 6318 245838
rect 6402 245602 6638 245838
rect 6722 245602 6958 245838
rect 7042 245602 7278 245838
rect 7362 245602 7598 245838
rect 7682 245602 7918 245838
rect 8002 245602 8238 245838
rect 8322 245602 8558 245838
rect 8642 245602 8878 245838
rect 5122 245282 5358 245518
rect 5442 245282 5678 245518
rect 5762 245282 5998 245518
rect 6082 245282 6318 245518
rect 6402 245282 6638 245518
rect 6722 245282 6958 245518
rect 7042 245282 7278 245518
rect 7362 245282 7598 245518
rect 7682 245282 7918 245518
rect 8002 245282 8238 245518
rect 8322 245282 8558 245518
rect 8642 245282 8878 245518
rect 5122 244962 5358 245198
rect 5442 244962 5678 245198
rect 5762 244962 5998 245198
rect 6082 244962 6318 245198
rect 6402 244962 6638 245198
rect 6722 244962 6958 245198
rect 7042 244962 7278 245198
rect 7362 244962 7598 245198
rect 7682 244962 7918 245198
rect 8002 244962 8238 245198
rect 8322 244962 8558 245198
rect 8642 244962 8878 245198
rect 5122 244642 5358 244878
rect 5442 244642 5678 244878
rect 5762 244642 5998 244878
rect 6082 244642 6318 244878
rect 6402 244642 6638 244878
rect 6722 244642 6958 244878
rect 7042 244642 7278 244878
rect 7362 244642 7598 244878
rect 7682 244642 7918 244878
rect 8002 244642 8238 244878
rect 8322 244642 8558 244878
rect 8642 244642 8878 244878
rect 5122 244322 5358 244558
rect 5442 244322 5678 244558
rect 5762 244322 5998 244558
rect 6082 244322 6318 244558
rect 6402 244322 6638 244558
rect 6722 244322 6958 244558
rect 7042 244322 7278 244558
rect 7362 244322 7598 244558
rect 7682 244322 7918 244558
rect 8002 244322 8238 244558
rect 8322 244322 8558 244558
rect 8642 244322 8878 244558
rect 5122 239882 5358 240118
rect 5442 239882 5678 240118
rect 5762 239882 5998 240118
rect 6082 239882 6318 240118
rect 6402 239882 6638 240118
rect 6722 239882 6958 240118
rect 7042 239882 7278 240118
rect 7362 239882 7598 240118
rect 7682 239882 7918 240118
rect 8002 239882 8238 240118
rect 8322 239882 8558 240118
rect 8642 239882 8878 240118
rect 226838 247842 227074 248078
rect 227158 247842 227394 248078
rect 227478 247842 227714 248078
rect 227798 247842 228034 248078
rect 228118 247842 228354 248078
rect 228438 247842 228674 248078
rect 228758 247842 228994 248078
rect 229078 247842 229314 248078
rect 229398 247842 229634 248078
rect 229718 247842 229954 248078
rect 230038 247842 230274 248078
rect 230358 247842 230594 248078
rect 226838 247522 227074 247758
rect 227158 247522 227394 247758
rect 227478 247522 227714 247758
rect 227798 247522 228034 247758
rect 228118 247522 228354 247758
rect 228438 247522 228674 247758
rect 228758 247522 228994 247758
rect 229078 247522 229314 247758
rect 229398 247522 229634 247758
rect 229718 247522 229954 247758
rect 230038 247522 230274 247758
rect 230358 247522 230594 247758
rect 226838 247202 227074 247438
rect 227158 247202 227394 247438
rect 227478 247202 227714 247438
rect 227798 247202 228034 247438
rect 228118 247202 228354 247438
rect 228438 247202 228674 247438
rect 228758 247202 228994 247438
rect 229078 247202 229314 247438
rect 229398 247202 229634 247438
rect 229718 247202 229954 247438
rect 230038 247202 230274 247438
rect 230358 247202 230594 247438
rect 226838 246882 227074 247118
rect 227158 246882 227394 247118
rect 227478 246882 227714 247118
rect 227798 246882 228034 247118
rect 228118 246882 228354 247118
rect 228438 246882 228674 247118
rect 228758 246882 228994 247118
rect 229078 246882 229314 247118
rect 229398 246882 229634 247118
rect 229718 246882 229954 247118
rect 230038 246882 230274 247118
rect 230358 246882 230594 247118
rect 226838 246562 227074 246798
rect 227158 246562 227394 246798
rect 227478 246562 227714 246798
rect 227798 246562 228034 246798
rect 228118 246562 228354 246798
rect 228438 246562 228674 246798
rect 228758 246562 228994 246798
rect 229078 246562 229314 246798
rect 229398 246562 229634 246798
rect 229718 246562 229954 246798
rect 230038 246562 230274 246798
rect 230358 246562 230594 246798
rect 226838 246242 227074 246478
rect 227158 246242 227394 246478
rect 227478 246242 227714 246478
rect 227798 246242 228034 246478
rect 228118 246242 228354 246478
rect 228438 246242 228674 246478
rect 228758 246242 228994 246478
rect 229078 246242 229314 246478
rect 229398 246242 229634 246478
rect 229718 246242 229954 246478
rect 230038 246242 230274 246478
rect 230358 246242 230594 246478
rect 226838 245922 227074 246158
rect 227158 245922 227394 246158
rect 227478 245922 227714 246158
rect 227798 245922 228034 246158
rect 228118 245922 228354 246158
rect 228438 245922 228674 246158
rect 228758 245922 228994 246158
rect 229078 245922 229314 246158
rect 229398 245922 229634 246158
rect 229718 245922 229954 246158
rect 230038 245922 230274 246158
rect 230358 245922 230594 246158
rect 226838 245602 227074 245838
rect 227158 245602 227394 245838
rect 227478 245602 227714 245838
rect 227798 245602 228034 245838
rect 228118 245602 228354 245838
rect 228438 245602 228674 245838
rect 228758 245602 228994 245838
rect 229078 245602 229314 245838
rect 229398 245602 229634 245838
rect 229718 245602 229954 245838
rect 230038 245602 230274 245838
rect 230358 245602 230594 245838
rect 226838 245282 227074 245518
rect 227158 245282 227394 245518
rect 227478 245282 227714 245518
rect 227798 245282 228034 245518
rect 228118 245282 228354 245518
rect 228438 245282 228674 245518
rect 228758 245282 228994 245518
rect 229078 245282 229314 245518
rect 229398 245282 229634 245518
rect 229718 245282 229954 245518
rect 230038 245282 230274 245518
rect 230358 245282 230594 245518
rect 226838 244962 227074 245198
rect 227158 244962 227394 245198
rect 227478 244962 227714 245198
rect 227798 244962 228034 245198
rect 228118 244962 228354 245198
rect 228438 244962 228674 245198
rect 228758 244962 228994 245198
rect 229078 244962 229314 245198
rect 229398 244962 229634 245198
rect 229718 244962 229954 245198
rect 230038 244962 230274 245198
rect 230358 244962 230594 245198
rect 226838 244642 227074 244878
rect 227158 244642 227394 244878
rect 227478 244642 227714 244878
rect 227798 244642 228034 244878
rect 228118 244642 228354 244878
rect 228438 244642 228674 244878
rect 228758 244642 228994 244878
rect 229078 244642 229314 244878
rect 229398 244642 229634 244878
rect 229718 244642 229954 244878
rect 230038 244642 230274 244878
rect 230358 244642 230594 244878
rect 226838 244322 227074 244558
rect 227158 244322 227394 244558
rect 227478 244322 227714 244558
rect 227798 244322 228034 244558
rect 228118 244322 228354 244558
rect 228438 244322 228674 244558
rect 228758 244322 228994 244558
rect 229078 244322 229314 244558
rect 229398 244322 229634 244558
rect 229718 244322 229954 244558
rect 230038 244322 230274 244558
rect 230358 244322 230594 244558
rect 226838 239882 227074 240118
rect 227158 239882 227394 240118
rect 227478 239882 227714 240118
rect 227798 239882 228034 240118
rect 228118 239882 228354 240118
rect 228438 239882 228674 240118
rect 228758 239882 228994 240118
rect 229078 239882 229314 240118
rect 229398 239882 229634 240118
rect 229718 239882 229954 240118
rect 230038 239882 230274 240118
rect 230358 239882 230594 240118
rect 30215 228682 30451 228918
rect 71882 228682 72118 228918
rect 5122 217482 5358 217718
rect 5442 217482 5678 217718
rect 5762 217482 5998 217718
rect 6082 217482 6318 217718
rect 6402 217482 6638 217718
rect 6722 217482 6958 217718
rect 7042 217482 7278 217718
rect 7362 217482 7598 217718
rect 7682 217482 7918 217718
rect 8002 217482 8238 217718
rect 8322 217482 8558 217718
rect 8642 217482 8878 217718
rect 25549 217482 25785 217718
rect 66882 217482 67118 217718
rect 114215 228682 114451 228918
rect 155882 228682 156118 228918
rect 109549 217482 109785 217718
rect 150882 217482 151118 217718
rect 198215 228682 198451 228918
rect 193549 217482 193785 217718
rect 226838 217482 227074 217718
rect 227158 217482 227394 217718
rect 227478 217482 227714 217718
rect 227798 217482 228034 217718
rect 228118 217482 228354 217718
rect 228438 217482 228674 217718
rect 228758 217482 228994 217718
rect 229078 217482 229314 217718
rect 229398 217482 229634 217718
rect 229718 217482 229954 217718
rect 230038 217482 230274 217718
rect 230358 217482 230594 217718
rect 5122 195082 5358 195318
rect 5442 195082 5678 195318
rect 5762 195082 5998 195318
rect 6082 195082 6318 195318
rect 6402 195082 6638 195318
rect 6722 195082 6958 195318
rect 7042 195082 7278 195318
rect 7362 195082 7598 195318
rect 7682 195082 7918 195318
rect 8002 195082 8238 195318
rect 8322 195082 8558 195318
rect 8642 195082 8878 195318
rect 32215 183882 32451 184118
rect 75506 183882 75742 184118
rect 116215 183882 116451 184118
rect 5122 172682 5358 172918
rect 5442 172682 5678 172918
rect 5762 172682 5998 172918
rect 6082 172682 6318 172918
rect 6402 172682 6638 172918
rect 6722 172682 6958 172918
rect 7042 172682 7278 172918
rect 7362 172682 7598 172918
rect 7682 172682 7918 172918
rect 8002 172682 8238 172918
rect 8322 172682 8558 172918
rect 8642 172682 8878 172918
rect 29549 172682 29785 172918
rect 60146 172682 60382 172918
rect 113549 172682 113785 172918
rect 32215 161482 32451 161718
rect 75506 161482 75742 161718
rect 116215 161482 116451 161718
rect 137934 156756 138170 156842
rect 137934 156692 138020 156756
rect 138020 156692 138084 156756
rect 138084 156692 138170 156756
rect 137934 156606 138170 156692
rect 5122 150282 5358 150518
rect 5442 150282 5678 150518
rect 5762 150282 5998 150518
rect 6082 150282 6318 150518
rect 6402 150282 6638 150518
rect 6722 150282 6958 150518
rect 7042 150282 7278 150518
rect 7362 150282 7598 150518
rect 7682 150282 7918 150518
rect 8002 150282 8238 150518
rect 8322 150282 8558 150518
rect 8642 150282 8878 150518
rect 5122 127882 5358 128118
rect 5442 127882 5678 128118
rect 5762 127882 5998 128118
rect 6082 127882 6318 128118
rect 6402 127882 6638 128118
rect 6722 127882 6958 128118
rect 7042 127882 7278 128118
rect 7362 127882 7598 128118
rect 7682 127882 7918 128118
rect 8002 127882 8238 128118
rect 8322 127882 8558 128118
rect 8642 127882 8878 128118
rect 25549 127882 25785 128118
rect 66882 127882 67118 128118
rect 109549 127882 109785 128118
rect 30215 116682 30451 116918
rect 114215 116682 114451 116918
rect 5122 105482 5358 105718
rect 5442 105482 5678 105718
rect 5762 105482 5998 105718
rect 6082 105482 6318 105718
rect 6402 105482 6638 105718
rect 6722 105482 6958 105718
rect 7042 105482 7278 105718
rect 7362 105482 7598 105718
rect 7682 105482 7918 105718
rect 8002 105482 8238 105718
rect 8322 105482 8558 105718
rect 8642 105482 8878 105718
rect 32215 94282 32451 94518
rect 75506 94282 75742 94518
rect 116215 94282 116451 94518
rect 5122 83082 5358 83318
rect 5442 83082 5678 83318
rect 5762 83082 5998 83318
rect 6082 83082 6318 83318
rect 6402 83082 6638 83318
rect 6722 83082 6958 83318
rect 7042 83082 7278 83318
rect 7362 83082 7598 83318
rect 7682 83082 7918 83318
rect 8002 83082 8238 83318
rect 8322 83082 8558 83318
rect 8642 83082 8878 83318
rect 29549 83082 29785 83318
rect 60146 83082 60382 83318
rect 113549 83082 113785 83318
rect 32215 71882 32451 72118
rect 75506 71882 75742 72118
rect 116215 71882 116451 72118
rect 13182 66846 13418 67082
rect 55870 66846 56106 67082
rect 5122 60682 5358 60918
rect 5442 60682 5678 60918
rect 5762 60682 5998 60918
rect 6082 60682 6318 60918
rect 6402 60682 6638 60918
rect 6722 60682 6958 60918
rect 7042 60682 7278 60918
rect 7362 60682 7598 60918
rect 7682 60682 7918 60918
rect 8002 60682 8238 60918
rect 8322 60682 8558 60918
rect 8642 60682 8878 60918
rect 226838 195082 227074 195318
rect 227158 195082 227394 195318
rect 227478 195082 227714 195318
rect 227798 195082 228034 195318
rect 228118 195082 228354 195318
rect 228438 195082 228674 195318
rect 228758 195082 228994 195318
rect 229078 195082 229314 195318
rect 229398 195082 229634 195318
rect 229718 195082 229954 195318
rect 230038 195082 230274 195318
rect 230358 195082 230594 195318
rect 193870 190620 194106 190842
rect 193870 190606 193956 190620
rect 193956 190606 194020 190620
rect 194020 190606 194106 190620
rect 209878 190756 210114 190842
rect 209878 190692 209964 190756
rect 209964 190692 210028 190756
rect 210028 190692 210114 190756
rect 209878 190606 210114 190692
rect 159506 183882 159742 184118
rect 200215 183882 200451 184118
rect 144146 172682 144382 172918
rect 197549 172682 197785 172918
rect 226838 172682 227074 172918
rect 227158 172682 227394 172918
rect 227478 172682 227714 172918
rect 227798 172682 228034 172918
rect 228118 172682 228354 172918
rect 228438 172682 228674 172918
rect 228758 172682 228994 172918
rect 229078 172682 229314 172918
rect 229398 172682 229634 172918
rect 229718 172682 229954 172918
rect 230038 172682 230274 172918
rect 230358 172682 230594 172918
rect 159506 161482 159742 161718
rect 200215 161482 200451 161718
rect 209694 156756 209930 156842
rect 209694 156692 209780 156756
rect 209780 156692 209844 156756
rect 209844 156692 209930 156756
rect 209694 156606 209930 156692
rect 226838 150282 227074 150518
rect 227158 150282 227394 150518
rect 227478 150282 227714 150518
rect 227798 150282 228034 150518
rect 228118 150282 228354 150518
rect 228438 150282 228674 150518
rect 228758 150282 228994 150518
rect 229078 150282 229314 150518
rect 229398 150282 229634 150518
rect 229718 150282 229954 150518
rect 230038 150282 230274 150518
rect 230358 150282 230594 150518
rect 150882 127882 151118 128118
rect 193549 127882 193785 128118
rect 226838 127882 227074 128118
rect 227158 127882 227394 128118
rect 227478 127882 227714 128118
rect 227798 127882 228034 128118
rect 228118 127882 228354 128118
rect 228438 127882 228674 128118
rect 228758 127882 228994 128118
rect 229078 127882 229314 128118
rect 229398 127882 229634 128118
rect 229718 127882 229954 128118
rect 230038 127882 230274 128118
rect 230358 127882 230594 128118
rect 198215 116682 198451 116918
rect 226838 105482 227074 105718
rect 227158 105482 227394 105718
rect 227478 105482 227714 105718
rect 227798 105482 228034 105718
rect 228118 105482 228354 105718
rect 228438 105482 228674 105718
rect 228758 105482 228994 105718
rect 229078 105482 229314 105718
rect 229398 105482 229634 105718
rect 229718 105482 229954 105718
rect 230038 105482 230274 105718
rect 230358 105482 230594 105718
rect 193686 96916 193922 97002
rect 193686 96852 193772 96916
rect 193772 96852 193836 96916
rect 193836 96852 193922 96916
rect 193686 96766 193922 96852
rect 209694 96780 209930 97002
rect 209694 96766 209780 96780
rect 209780 96766 209844 96780
rect 209844 96766 209930 96780
rect 159506 94282 159742 94518
rect 200215 94282 200451 94518
rect 144146 83082 144382 83318
rect 197549 83082 197785 83318
rect 226838 83082 227074 83318
rect 227158 83082 227394 83318
rect 227478 83082 227714 83318
rect 227798 83082 228034 83318
rect 228118 83082 228354 83318
rect 228438 83082 228674 83318
rect 228758 83082 228994 83318
rect 229078 83082 229314 83318
rect 229398 83082 229634 83318
rect 229718 83082 229954 83318
rect 230038 83082 230274 83318
rect 230358 83082 230594 83318
rect 159506 71882 159742 72118
rect 200215 71882 200451 72118
rect 226838 60682 227074 60918
rect 227158 60682 227394 60918
rect 227478 60682 227714 60918
rect 227798 60682 228034 60918
rect 228118 60682 228354 60918
rect 228438 60682 228674 60918
rect 228758 60682 228994 60918
rect 229078 60682 229314 60918
rect 229398 60682 229634 60918
rect 229718 60682 229954 60918
rect 230038 60682 230274 60918
rect 230358 60682 230594 60918
rect 5122 38282 5358 38518
rect 5442 38282 5678 38518
rect 5762 38282 5998 38518
rect 6082 38282 6318 38518
rect 6402 38282 6638 38518
rect 6722 38282 6958 38518
rect 7042 38282 7278 38518
rect 7362 38282 7598 38518
rect 7682 38282 7918 38518
rect 8002 38282 8238 38518
rect 8322 38282 8558 38518
rect 8642 38282 8878 38518
rect 25549 38282 25785 38518
rect 30215 27082 30451 27318
rect 66882 38282 67118 38518
rect 71882 27082 72118 27318
rect 88990 20606 89226 20842
rect 109549 38282 109785 38518
rect 114215 27082 114451 27318
rect 101502 20756 101738 20842
rect 101502 20692 101588 20756
rect 101588 20692 101652 20756
rect 101652 20692 101738 20756
rect 101502 20606 101738 20692
rect 89726 19926 89962 20162
rect 101502 20076 101738 20162
rect 101502 20012 101588 20076
rect 101588 20012 101652 20076
rect 101652 20012 101738 20076
rect 101502 19926 101738 20012
rect 154862 43046 155098 43282
rect 159462 43046 159698 43282
rect 151550 40326 151786 40562
rect 150446 39646 150682 39882
rect 150882 38282 151118 38518
rect 150446 21966 150682 22202
rect 155882 27082 156118 27318
rect 155966 21966 156202 22202
rect 173078 20606 173314 20842
rect 193549 38282 193785 38518
rect 226838 38282 227074 38518
rect 227158 38282 227394 38518
rect 227478 38282 227714 38518
rect 227798 38282 228034 38518
rect 228118 38282 228354 38518
rect 228438 38282 228674 38518
rect 228758 38282 228994 38518
rect 229078 38282 229314 38518
rect 229398 38282 229634 38518
rect 229718 38282 229954 38518
rect 230038 38282 230274 38518
rect 230358 38282 230594 38518
rect 212638 35566 212874 35802
rect 212638 34886 212874 35122
rect 198215 27082 198451 27318
rect 212638 25366 212874 25602
rect 212638 24686 212874 24922
rect 173814 21966 174050 22202
rect 185038 21980 185274 22202
rect 185038 21966 185124 21980
rect 185124 21966 185188 21980
rect 185188 21966 185274 21980
rect 212638 21286 212874 21522
rect 222206 21286 222442 21522
rect 185038 20756 185274 20842
rect 185038 20692 185124 20756
rect 185124 20692 185188 20756
rect 185188 20692 185274 20756
rect 185038 20606 185274 20692
rect 173446 19926 173682 20162
rect 185406 19926 185642 20162
rect 5122 15882 5358 16118
rect 5442 15882 5678 16118
rect 5762 15882 5998 16118
rect 6082 15882 6318 16118
rect 6402 15882 6638 16118
rect 6722 15882 6958 16118
rect 7042 15882 7278 16118
rect 7362 15882 7598 16118
rect 7682 15882 7918 16118
rect 8002 15882 8238 16118
rect 8322 15882 8558 16118
rect 8642 15882 8878 16118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 226838 15882 227074 16118
rect 227158 15882 227394 16118
rect 227478 15882 227714 16118
rect 227798 15882 228034 16118
rect 228118 15882 228354 16118
rect 228438 15882 228674 16118
rect 228758 15882 228994 16118
rect 229078 15882 229314 16118
rect 229398 15882 229634 16118
rect 229718 15882 229954 16118
rect 230038 15882 230274 16118
rect 230358 15882 230594 16118
rect 226838 8642 227074 8878
rect 227158 8642 227394 8878
rect 227478 8642 227714 8878
rect 227798 8642 228034 8878
rect 228118 8642 228354 8878
rect 228438 8642 228674 8878
rect 228758 8642 228994 8878
rect 229078 8642 229314 8878
rect 229398 8642 229634 8878
rect 229718 8642 229954 8878
rect 230038 8642 230274 8878
rect 230358 8642 230594 8878
rect 226838 8322 227074 8558
rect 227158 8322 227394 8558
rect 227478 8322 227714 8558
rect 227798 8322 228034 8558
rect 228118 8322 228354 8558
rect 228438 8322 228674 8558
rect 228758 8322 228994 8558
rect 229078 8322 229314 8558
rect 229398 8322 229634 8558
rect 229718 8322 229954 8558
rect 230038 8322 230274 8558
rect 230358 8322 230594 8558
rect 226838 8002 227074 8238
rect 227158 8002 227394 8238
rect 227478 8002 227714 8238
rect 227798 8002 228034 8238
rect 228118 8002 228354 8238
rect 228438 8002 228674 8238
rect 228758 8002 228994 8238
rect 229078 8002 229314 8238
rect 229398 8002 229634 8238
rect 229718 8002 229954 8238
rect 230038 8002 230274 8238
rect 230358 8002 230594 8238
rect 226838 7682 227074 7918
rect 227158 7682 227394 7918
rect 227478 7682 227714 7918
rect 227798 7682 228034 7918
rect 228118 7682 228354 7918
rect 228438 7682 228674 7918
rect 228758 7682 228994 7918
rect 229078 7682 229314 7918
rect 229398 7682 229634 7918
rect 229718 7682 229954 7918
rect 230038 7682 230274 7918
rect 230358 7682 230594 7918
rect 226838 7362 227074 7598
rect 227158 7362 227394 7598
rect 227478 7362 227714 7598
rect 227798 7362 228034 7598
rect 228118 7362 228354 7598
rect 228438 7362 228674 7598
rect 228758 7362 228994 7598
rect 229078 7362 229314 7598
rect 229398 7362 229634 7598
rect 229718 7362 229954 7598
rect 230038 7362 230274 7598
rect 230358 7362 230594 7598
rect 226838 7042 227074 7278
rect 227158 7042 227394 7278
rect 227478 7042 227714 7278
rect 227798 7042 228034 7278
rect 228118 7042 228354 7278
rect 228438 7042 228674 7278
rect 228758 7042 228994 7278
rect 229078 7042 229314 7278
rect 229398 7042 229634 7278
rect 229718 7042 229954 7278
rect 230038 7042 230274 7278
rect 230358 7042 230594 7278
rect 226838 6722 227074 6958
rect 227158 6722 227394 6958
rect 227478 6722 227714 6958
rect 227798 6722 228034 6958
rect 228118 6722 228354 6958
rect 228438 6722 228674 6958
rect 228758 6722 228994 6958
rect 229078 6722 229314 6958
rect 229398 6722 229634 6958
rect 229718 6722 229954 6958
rect 230038 6722 230274 6958
rect 230358 6722 230594 6958
rect 226838 6402 227074 6638
rect 227158 6402 227394 6638
rect 227478 6402 227714 6638
rect 227798 6402 228034 6638
rect 228118 6402 228354 6638
rect 228438 6402 228674 6638
rect 228758 6402 228994 6638
rect 229078 6402 229314 6638
rect 229398 6402 229634 6638
rect 229718 6402 229954 6638
rect 230038 6402 230274 6638
rect 230358 6402 230594 6638
rect 226838 6082 227074 6318
rect 227158 6082 227394 6318
rect 227478 6082 227714 6318
rect 227798 6082 228034 6318
rect 228118 6082 228354 6318
rect 228438 6082 228674 6318
rect 228758 6082 228994 6318
rect 229078 6082 229314 6318
rect 229398 6082 229634 6318
rect 229718 6082 229954 6318
rect 230038 6082 230274 6318
rect 230358 6082 230594 6318
rect 226838 5762 227074 5998
rect 227158 5762 227394 5998
rect 227478 5762 227714 5998
rect 227798 5762 228034 5998
rect 228118 5762 228354 5998
rect 228438 5762 228674 5998
rect 228758 5762 228994 5998
rect 229078 5762 229314 5998
rect 229398 5762 229634 5998
rect 229718 5762 229954 5998
rect 230038 5762 230274 5998
rect 230358 5762 230594 5998
rect 226838 5442 227074 5678
rect 227158 5442 227394 5678
rect 227478 5442 227714 5678
rect 227798 5442 228034 5678
rect 228118 5442 228354 5678
rect 228438 5442 228674 5678
rect 228758 5442 228994 5678
rect 229078 5442 229314 5678
rect 229398 5442 229634 5678
rect 229718 5442 229954 5678
rect 230038 5442 230274 5678
rect 230358 5442 230594 5678
rect 226838 5122 227074 5358
rect 227158 5122 227394 5358
rect 227478 5122 227714 5358
rect 227798 5122 228034 5358
rect 228118 5122 228354 5358
rect 228438 5122 228674 5358
rect 228758 5122 228994 5358
rect 229078 5122 229314 5358
rect 229398 5122 229634 5358
rect 229718 5122 229954 5358
rect 230038 5122 230274 5358
rect 230358 5122 230594 5358
rect 231838 228682 232074 228918
rect 232158 228682 232394 228918
rect 232478 228682 232714 228918
rect 232798 228682 233034 228918
rect 233118 228682 233354 228918
rect 233438 228682 233674 228918
rect 233758 228682 233994 228918
rect 234078 228682 234314 228918
rect 234398 228682 234634 228918
rect 234718 228682 234954 228918
rect 235038 228682 235274 228918
rect 235358 228682 235594 228918
rect 231838 206282 232074 206518
rect 232158 206282 232394 206518
rect 232478 206282 232714 206518
rect 232798 206282 233034 206518
rect 233118 206282 233354 206518
rect 233438 206282 233674 206518
rect 233758 206282 233994 206518
rect 234078 206282 234314 206518
rect 234398 206282 234634 206518
rect 234718 206282 234954 206518
rect 235038 206282 235274 206518
rect 235358 206282 235594 206518
rect 231838 183882 232074 184118
rect 232158 183882 232394 184118
rect 232478 183882 232714 184118
rect 232798 183882 233034 184118
rect 233118 183882 233354 184118
rect 233438 183882 233674 184118
rect 233758 183882 233994 184118
rect 234078 183882 234314 184118
rect 234398 183882 234634 184118
rect 234718 183882 234954 184118
rect 235038 183882 235274 184118
rect 235358 183882 235594 184118
rect 231838 161482 232074 161718
rect 232158 161482 232394 161718
rect 232478 161482 232714 161718
rect 232798 161482 233034 161718
rect 233118 161482 233354 161718
rect 233438 161482 233674 161718
rect 233758 161482 233994 161718
rect 234078 161482 234314 161718
rect 234398 161482 234634 161718
rect 234718 161482 234954 161718
rect 235038 161482 235274 161718
rect 235358 161482 235594 161718
rect 231838 139082 232074 139318
rect 232158 139082 232394 139318
rect 232478 139082 232714 139318
rect 232798 139082 233034 139318
rect 233118 139082 233354 139318
rect 233438 139082 233674 139318
rect 233758 139082 233994 139318
rect 234078 139082 234314 139318
rect 234398 139082 234634 139318
rect 234718 139082 234954 139318
rect 235038 139082 235274 139318
rect 235358 139082 235594 139318
rect 231838 116682 232074 116918
rect 232158 116682 232394 116918
rect 232478 116682 232714 116918
rect 232798 116682 233034 116918
rect 233118 116682 233354 116918
rect 233438 116682 233674 116918
rect 233758 116682 233994 116918
rect 234078 116682 234314 116918
rect 234398 116682 234634 116918
rect 234718 116682 234954 116918
rect 235038 116682 235274 116918
rect 235358 116682 235594 116918
rect 231838 94282 232074 94518
rect 232158 94282 232394 94518
rect 232478 94282 232714 94518
rect 232798 94282 233034 94518
rect 233118 94282 233354 94518
rect 233438 94282 233674 94518
rect 233758 94282 233994 94518
rect 234078 94282 234314 94518
rect 234398 94282 234634 94518
rect 234718 94282 234954 94518
rect 235038 94282 235274 94518
rect 235358 94282 235594 94518
rect 231838 71882 232074 72118
rect 232158 71882 232394 72118
rect 232478 71882 232714 72118
rect 232798 71882 233034 72118
rect 233118 71882 233354 72118
rect 233438 71882 233674 72118
rect 233758 71882 233994 72118
rect 234078 71882 234314 72118
rect 234398 71882 234634 72118
rect 234718 71882 234954 72118
rect 235038 71882 235274 72118
rect 235358 71882 235594 72118
rect 231838 49482 232074 49718
rect 232158 49482 232394 49718
rect 232478 49482 232714 49718
rect 232798 49482 233034 49718
rect 233118 49482 233354 49718
rect 233438 49482 233674 49718
rect 233758 49482 233994 49718
rect 234078 49482 234314 49718
rect 234398 49482 234634 49718
rect 234718 49482 234954 49718
rect 235038 49482 235274 49718
rect 235358 49482 235594 49718
rect 231838 27082 232074 27318
rect 232158 27082 232394 27318
rect 232478 27082 232714 27318
rect 232798 27082 233034 27318
rect 233118 27082 233354 27318
rect 233438 27082 233674 27318
rect 233758 27082 233994 27318
rect 234078 27082 234314 27318
rect 234398 27082 234634 27318
rect 234718 27082 234954 27318
rect 235038 27082 235274 27318
rect 235358 27082 235594 27318
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 231838 3642 232074 3878
rect 232158 3642 232394 3878
rect 232478 3642 232714 3878
rect 232798 3642 233034 3878
rect 233118 3642 233354 3878
rect 233438 3642 233674 3878
rect 233758 3642 233994 3878
rect 234078 3642 234314 3878
rect 234398 3642 234634 3878
rect 234718 3642 234954 3878
rect 235038 3642 235274 3878
rect 235358 3642 235594 3878
rect 231838 3322 232074 3558
rect 232158 3322 232394 3558
rect 232478 3322 232714 3558
rect 232798 3322 233034 3558
rect 233118 3322 233354 3558
rect 233438 3322 233674 3558
rect 233758 3322 233994 3558
rect 234078 3322 234314 3558
rect 234398 3322 234634 3558
rect 234718 3322 234954 3558
rect 235038 3322 235274 3558
rect 235358 3322 235594 3558
rect 231838 3002 232074 3238
rect 232158 3002 232394 3238
rect 232478 3002 232714 3238
rect 232798 3002 233034 3238
rect 233118 3002 233354 3238
rect 233438 3002 233674 3238
rect 233758 3002 233994 3238
rect 234078 3002 234314 3238
rect 234398 3002 234634 3238
rect 234718 3002 234954 3238
rect 235038 3002 235274 3238
rect 235358 3002 235594 3238
rect 231838 2682 232074 2918
rect 232158 2682 232394 2918
rect 232478 2682 232714 2918
rect 232798 2682 233034 2918
rect 233118 2682 233354 2918
rect 233438 2682 233674 2918
rect 233758 2682 233994 2918
rect 234078 2682 234314 2918
rect 234398 2682 234634 2918
rect 234718 2682 234954 2918
rect 235038 2682 235274 2918
rect 235358 2682 235594 2918
rect 231838 2362 232074 2598
rect 232158 2362 232394 2598
rect 232478 2362 232714 2598
rect 232798 2362 233034 2598
rect 233118 2362 233354 2598
rect 233438 2362 233674 2598
rect 233758 2362 233994 2598
rect 234078 2362 234314 2598
rect 234398 2362 234634 2598
rect 234718 2362 234954 2598
rect 235038 2362 235274 2598
rect 235358 2362 235594 2598
rect 231838 2042 232074 2278
rect 232158 2042 232394 2278
rect 232478 2042 232714 2278
rect 232798 2042 233034 2278
rect 233118 2042 233354 2278
rect 233438 2042 233674 2278
rect 233758 2042 233994 2278
rect 234078 2042 234314 2278
rect 234398 2042 234634 2278
rect 234718 2042 234954 2278
rect 235038 2042 235274 2278
rect 235358 2042 235594 2278
rect 231838 1722 232074 1958
rect 232158 1722 232394 1958
rect 232478 1722 232714 1958
rect 232798 1722 233034 1958
rect 233118 1722 233354 1958
rect 233438 1722 233674 1958
rect 233758 1722 233994 1958
rect 234078 1722 234314 1958
rect 234398 1722 234634 1958
rect 234718 1722 234954 1958
rect 235038 1722 235274 1958
rect 235358 1722 235594 1958
rect 231838 1402 232074 1638
rect 232158 1402 232394 1638
rect 232478 1402 232714 1638
rect 232798 1402 233034 1638
rect 233118 1402 233354 1638
rect 233438 1402 233674 1638
rect 233758 1402 233994 1638
rect 234078 1402 234314 1638
rect 234398 1402 234634 1638
rect 234718 1402 234954 1638
rect 235038 1402 235274 1638
rect 235358 1402 235594 1638
rect 231838 1082 232074 1318
rect 232158 1082 232394 1318
rect 232478 1082 232714 1318
rect 232798 1082 233034 1318
rect 233118 1082 233354 1318
rect 233438 1082 233674 1318
rect 233758 1082 233994 1318
rect 234078 1082 234314 1318
rect 234398 1082 234634 1318
rect 234718 1082 234954 1318
rect 235038 1082 235274 1318
rect 235358 1082 235594 1318
rect 231838 762 232074 998
rect 232158 762 232394 998
rect 232478 762 232714 998
rect 232798 762 233034 998
rect 233118 762 233354 998
rect 233438 762 233674 998
rect 233758 762 233994 998
rect 234078 762 234314 998
rect 234398 762 234634 998
rect 234718 762 234954 998
rect 235038 762 235274 998
rect 235358 762 235594 998
rect 231838 442 232074 678
rect 232158 442 232394 678
rect 232478 442 232714 678
rect 232798 442 233034 678
rect 233118 442 233354 678
rect 233438 442 233674 678
rect 233758 442 233994 678
rect 234078 442 234314 678
rect 234398 442 234634 678
rect 234718 442 234954 678
rect 235038 442 235274 678
rect 235358 442 235594 678
rect 231838 122 232074 358
rect 232158 122 232394 358
rect 232478 122 232714 358
rect 232798 122 233034 358
rect 233118 122 233354 358
rect 233438 122 233674 358
rect 233758 122 233994 358
rect 234078 122 234314 358
rect 234398 122 234634 358
rect 234718 122 234954 358
rect 235038 122 235274 358
rect 235358 122 235594 358
<< metal5 >>
rect 0 253078 235716 253200
rect 0 252842 122 253078
rect 358 252842 442 253078
rect 678 252842 762 253078
rect 998 252842 1082 253078
rect 1318 252842 1402 253078
rect 1638 252842 1722 253078
rect 1958 252842 2042 253078
rect 2278 252842 2362 253078
rect 2598 252842 2682 253078
rect 2918 252842 3002 253078
rect 3238 252842 3322 253078
rect 3558 252842 3642 253078
rect 3878 252842 231838 253078
rect 232074 252842 232158 253078
rect 232394 252842 232478 253078
rect 232714 252842 232798 253078
rect 233034 252842 233118 253078
rect 233354 252842 233438 253078
rect 233674 252842 233758 253078
rect 233994 252842 234078 253078
rect 234314 252842 234398 253078
rect 234634 252842 234718 253078
rect 234954 252842 235038 253078
rect 235274 252842 235358 253078
rect 235594 252842 235716 253078
rect 0 252758 235716 252842
rect 0 252522 122 252758
rect 358 252522 442 252758
rect 678 252522 762 252758
rect 998 252522 1082 252758
rect 1318 252522 1402 252758
rect 1638 252522 1722 252758
rect 1958 252522 2042 252758
rect 2278 252522 2362 252758
rect 2598 252522 2682 252758
rect 2918 252522 3002 252758
rect 3238 252522 3322 252758
rect 3558 252522 3642 252758
rect 3878 252522 231838 252758
rect 232074 252522 232158 252758
rect 232394 252522 232478 252758
rect 232714 252522 232798 252758
rect 233034 252522 233118 252758
rect 233354 252522 233438 252758
rect 233674 252522 233758 252758
rect 233994 252522 234078 252758
rect 234314 252522 234398 252758
rect 234634 252522 234718 252758
rect 234954 252522 235038 252758
rect 235274 252522 235358 252758
rect 235594 252522 235716 252758
rect 0 252438 235716 252522
rect 0 252202 122 252438
rect 358 252202 442 252438
rect 678 252202 762 252438
rect 998 252202 1082 252438
rect 1318 252202 1402 252438
rect 1638 252202 1722 252438
rect 1958 252202 2042 252438
rect 2278 252202 2362 252438
rect 2598 252202 2682 252438
rect 2918 252202 3002 252438
rect 3238 252202 3322 252438
rect 3558 252202 3642 252438
rect 3878 252202 231838 252438
rect 232074 252202 232158 252438
rect 232394 252202 232478 252438
rect 232714 252202 232798 252438
rect 233034 252202 233118 252438
rect 233354 252202 233438 252438
rect 233674 252202 233758 252438
rect 233994 252202 234078 252438
rect 234314 252202 234398 252438
rect 234634 252202 234718 252438
rect 234954 252202 235038 252438
rect 235274 252202 235358 252438
rect 235594 252202 235716 252438
rect 0 252118 235716 252202
rect 0 251882 122 252118
rect 358 251882 442 252118
rect 678 251882 762 252118
rect 998 251882 1082 252118
rect 1318 251882 1402 252118
rect 1638 251882 1722 252118
rect 1958 251882 2042 252118
rect 2278 251882 2362 252118
rect 2598 251882 2682 252118
rect 2918 251882 3002 252118
rect 3238 251882 3322 252118
rect 3558 251882 3642 252118
rect 3878 251882 231838 252118
rect 232074 251882 232158 252118
rect 232394 251882 232478 252118
rect 232714 251882 232798 252118
rect 233034 251882 233118 252118
rect 233354 251882 233438 252118
rect 233674 251882 233758 252118
rect 233994 251882 234078 252118
rect 234314 251882 234398 252118
rect 234634 251882 234718 252118
rect 234954 251882 235038 252118
rect 235274 251882 235358 252118
rect 235594 251882 235716 252118
rect 0 251798 235716 251882
rect 0 251562 122 251798
rect 358 251562 442 251798
rect 678 251562 762 251798
rect 998 251562 1082 251798
rect 1318 251562 1402 251798
rect 1638 251562 1722 251798
rect 1958 251562 2042 251798
rect 2278 251562 2362 251798
rect 2598 251562 2682 251798
rect 2918 251562 3002 251798
rect 3238 251562 3322 251798
rect 3558 251562 3642 251798
rect 3878 251562 231838 251798
rect 232074 251562 232158 251798
rect 232394 251562 232478 251798
rect 232714 251562 232798 251798
rect 233034 251562 233118 251798
rect 233354 251562 233438 251798
rect 233674 251562 233758 251798
rect 233994 251562 234078 251798
rect 234314 251562 234398 251798
rect 234634 251562 234718 251798
rect 234954 251562 235038 251798
rect 235274 251562 235358 251798
rect 235594 251562 235716 251798
rect 0 251478 235716 251562
rect 0 251242 122 251478
rect 358 251242 442 251478
rect 678 251242 762 251478
rect 998 251242 1082 251478
rect 1318 251242 1402 251478
rect 1638 251242 1722 251478
rect 1958 251242 2042 251478
rect 2278 251242 2362 251478
rect 2598 251242 2682 251478
rect 2918 251242 3002 251478
rect 3238 251242 3322 251478
rect 3558 251242 3642 251478
rect 3878 251242 231838 251478
rect 232074 251242 232158 251478
rect 232394 251242 232478 251478
rect 232714 251242 232798 251478
rect 233034 251242 233118 251478
rect 233354 251242 233438 251478
rect 233674 251242 233758 251478
rect 233994 251242 234078 251478
rect 234314 251242 234398 251478
rect 234634 251242 234718 251478
rect 234954 251242 235038 251478
rect 235274 251242 235358 251478
rect 235594 251242 235716 251478
rect 0 251158 235716 251242
rect 0 250922 122 251158
rect 358 250922 442 251158
rect 678 250922 762 251158
rect 998 250922 1082 251158
rect 1318 250922 1402 251158
rect 1638 250922 1722 251158
rect 1958 250922 2042 251158
rect 2278 250922 2362 251158
rect 2598 250922 2682 251158
rect 2918 250922 3002 251158
rect 3238 250922 3322 251158
rect 3558 250922 3642 251158
rect 3878 250922 231838 251158
rect 232074 250922 232158 251158
rect 232394 250922 232478 251158
rect 232714 250922 232798 251158
rect 233034 250922 233118 251158
rect 233354 250922 233438 251158
rect 233674 250922 233758 251158
rect 233994 250922 234078 251158
rect 234314 250922 234398 251158
rect 234634 250922 234718 251158
rect 234954 250922 235038 251158
rect 235274 250922 235358 251158
rect 235594 250922 235716 251158
rect 0 250838 235716 250922
rect 0 250602 122 250838
rect 358 250602 442 250838
rect 678 250602 762 250838
rect 998 250602 1082 250838
rect 1318 250602 1402 250838
rect 1638 250602 1722 250838
rect 1958 250602 2042 250838
rect 2278 250602 2362 250838
rect 2598 250602 2682 250838
rect 2918 250602 3002 250838
rect 3238 250602 3322 250838
rect 3558 250602 3642 250838
rect 3878 250602 231838 250838
rect 232074 250602 232158 250838
rect 232394 250602 232478 250838
rect 232714 250602 232798 250838
rect 233034 250602 233118 250838
rect 233354 250602 233438 250838
rect 233674 250602 233758 250838
rect 233994 250602 234078 250838
rect 234314 250602 234398 250838
rect 234634 250602 234718 250838
rect 234954 250602 235038 250838
rect 235274 250602 235358 250838
rect 235594 250602 235716 250838
rect 0 250518 235716 250602
rect 0 250282 122 250518
rect 358 250282 442 250518
rect 678 250282 762 250518
rect 998 250282 1082 250518
rect 1318 250282 1402 250518
rect 1638 250282 1722 250518
rect 1958 250282 2042 250518
rect 2278 250282 2362 250518
rect 2598 250282 2682 250518
rect 2918 250282 3002 250518
rect 3238 250282 3322 250518
rect 3558 250282 3642 250518
rect 3878 250282 231838 250518
rect 232074 250282 232158 250518
rect 232394 250282 232478 250518
rect 232714 250282 232798 250518
rect 233034 250282 233118 250518
rect 233354 250282 233438 250518
rect 233674 250282 233758 250518
rect 233994 250282 234078 250518
rect 234314 250282 234398 250518
rect 234634 250282 234718 250518
rect 234954 250282 235038 250518
rect 235274 250282 235358 250518
rect 235594 250282 235716 250518
rect 0 250198 235716 250282
rect 0 249962 122 250198
rect 358 249962 442 250198
rect 678 249962 762 250198
rect 998 249962 1082 250198
rect 1318 249962 1402 250198
rect 1638 249962 1722 250198
rect 1958 249962 2042 250198
rect 2278 249962 2362 250198
rect 2598 249962 2682 250198
rect 2918 249962 3002 250198
rect 3238 249962 3322 250198
rect 3558 249962 3642 250198
rect 3878 249962 231838 250198
rect 232074 249962 232158 250198
rect 232394 249962 232478 250198
rect 232714 249962 232798 250198
rect 233034 249962 233118 250198
rect 233354 249962 233438 250198
rect 233674 249962 233758 250198
rect 233994 249962 234078 250198
rect 234314 249962 234398 250198
rect 234634 249962 234718 250198
rect 234954 249962 235038 250198
rect 235274 249962 235358 250198
rect 235594 249962 235716 250198
rect 0 249878 235716 249962
rect 0 249642 122 249878
rect 358 249642 442 249878
rect 678 249642 762 249878
rect 998 249642 1082 249878
rect 1318 249642 1402 249878
rect 1638 249642 1722 249878
rect 1958 249642 2042 249878
rect 2278 249642 2362 249878
rect 2598 249642 2682 249878
rect 2918 249642 3002 249878
rect 3238 249642 3322 249878
rect 3558 249642 3642 249878
rect 3878 249642 231838 249878
rect 232074 249642 232158 249878
rect 232394 249642 232478 249878
rect 232714 249642 232798 249878
rect 233034 249642 233118 249878
rect 233354 249642 233438 249878
rect 233674 249642 233758 249878
rect 233994 249642 234078 249878
rect 234314 249642 234398 249878
rect 234634 249642 234718 249878
rect 234954 249642 235038 249878
rect 235274 249642 235358 249878
rect 235594 249642 235716 249878
rect 0 249558 235716 249642
rect 0 249322 122 249558
rect 358 249322 442 249558
rect 678 249322 762 249558
rect 998 249322 1082 249558
rect 1318 249322 1402 249558
rect 1638 249322 1722 249558
rect 1958 249322 2042 249558
rect 2278 249322 2362 249558
rect 2598 249322 2682 249558
rect 2918 249322 3002 249558
rect 3238 249322 3322 249558
rect 3558 249322 3642 249558
rect 3878 249322 231838 249558
rect 232074 249322 232158 249558
rect 232394 249322 232478 249558
rect 232714 249322 232798 249558
rect 233034 249322 233118 249558
rect 233354 249322 233438 249558
rect 233674 249322 233758 249558
rect 233994 249322 234078 249558
rect 234314 249322 234398 249558
rect 234634 249322 234718 249558
rect 234954 249322 235038 249558
rect 235274 249322 235358 249558
rect 235594 249322 235716 249558
rect 0 249200 235716 249322
rect 5000 248078 230716 248200
rect 5000 247842 5122 248078
rect 5358 247842 5442 248078
rect 5678 247842 5762 248078
rect 5998 247842 6082 248078
rect 6318 247842 6402 248078
rect 6638 247842 6722 248078
rect 6958 247842 7042 248078
rect 7278 247842 7362 248078
rect 7598 247842 7682 248078
rect 7918 247842 8002 248078
rect 8238 247842 8322 248078
rect 8558 247842 8642 248078
rect 8878 247842 226838 248078
rect 227074 247842 227158 248078
rect 227394 247842 227478 248078
rect 227714 247842 227798 248078
rect 228034 247842 228118 248078
rect 228354 247842 228438 248078
rect 228674 247842 228758 248078
rect 228994 247842 229078 248078
rect 229314 247842 229398 248078
rect 229634 247842 229718 248078
rect 229954 247842 230038 248078
rect 230274 247842 230358 248078
rect 230594 247842 230716 248078
rect 5000 247758 230716 247842
rect 5000 247522 5122 247758
rect 5358 247522 5442 247758
rect 5678 247522 5762 247758
rect 5998 247522 6082 247758
rect 6318 247522 6402 247758
rect 6638 247522 6722 247758
rect 6958 247522 7042 247758
rect 7278 247522 7362 247758
rect 7598 247522 7682 247758
rect 7918 247522 8002 247758
rect 8238 247522 8322 247758
rect 8558 247522 8642 247758
rect 8878 247522 226838 247758
rect 227074 247522 227158 247758
rect 227394 247522 227478 247758
rect 227714 247522 227798 247758
rect 228034 247522 228118 247758
rect 228354 247522 228438 247758
rect 228674 247522 228758 247758
rect 228994 247522 229078 247758
rect 229314 247522 229398 247758
rect 229634 247522 229718 247758
rect 229954 247522 230038 247758
rect 230274 247522 230358 247758
rect 230594 247522 230716 247758
rect 5000 247438 230716 247522
rect 5000 247202 5122 247438
rect 5358 247202 5442 247438
rect 5678 247202 5762 247438
rect 5998 247202 6082 247438
rect 6318 247202 6402 247438
rect 6638 247202 6722 247438
rect 6958 247202 7042 247438
rect 7278 247202 7362 247438
rect 7598 247202 7682 247438
rect 7918 247202 8002 247438
rect 8238 247202 8322 247438
rect 8558 247202 8642 247438
rect 8878 247202 226838 247438
rect 227074 247202 227158 247438
rect 227394 247202 227478 247438
rect 227714 247202 227798 247438
rect 228034 247202 228118 247438
rect 228354 247202 228438 247438
rect 228674 247202 228758 247438
rect 228994 247202 229078 247438
rect 229314 247202 229398 247438
rect 229634 247202 229718 247438
rect 229954 247202 230038 247438
rect 230274 247202 230358 247438
rect 230594 247202 230716 247438
rect 5000 247118 230716 247202
rect 5000 246882 5122 247118
rect 5358 246882 5442 247118
rect 5678 246882 5762 247118
rect 5998 246882 6082 247118
rect 6318 246882 6402 247118
rect 6638 246882 6722 247118
rect 6958 246882 7042 247118
rect 7278 246882 7362 247118
rect 7598 246882 7682 247118
rect 7918 246882 8002 247118
rect 8238 246882 8322 247118
rect 8558 246882 8642 247118
rect 8878 246882 226838 247118
rect 227074 246882 227158 247118
rect 227394 246882 227478 247118
rect 227714 246882 227798 247118
rect 228034 246882 228118 247118
rect 228354 246882 228438 247118
rect 228674 246882 228758 247118
rect 228994 246882 229078 247118
rect 229314 246882 229398 247118
rect 229634 246882 229718 247118
rect 229954 246882 230038 247118
rect 230274 246882 230358 247118
rect 230594 246882 230716 247118
rect 5000 246798 230716 246882
rect 5000 246562 5122 246798
rect 5358 246562 5442 246798
rect 5678 246562 5762 246798
rect 5998 246562 6082 246798
rect 6318 246562 6402 246798
rect 6638 246562 6722 246798
rect 6958 246562 7042 246798
rect 7278 246562 7362 246798
rect 7598 246562 7682 246798
rect 7918 246562 8002 246798
rect 8238 246562 8322 246798
rect 8558 246562 8642 246798
rect 8878 246562 226838 246798
rect 227074 246562 227158 246798
rect 227394 246562 227478 246798
rect 227714 246562 227798 246798
rect 228034 246562 228118 246798
rect 228354 246562 228438 246798
rect 228674 246562 228758 246798
rect 228994 246562 229078 246798
rect 229314 246562 229398 246798
rect 229634 246562 229718 246798
rect 229954 246562 230038 246798
rect 230274 246562 230358 246798
rect 230594 246562 230716 246798
rect 5000 246478 230716 246562
rect 5000 246242 5122 246478
rect 5358 246242 5442 246478
rect 5678 246242 5762 246478
rect 5998 246242 6082 246478
rect 6318 246242 6402 246478
rect 6638 246242 6722 246478
rect 6958 246242 7042 246478
rect 7278 246242 7362 246478
rect 7598 246242 7682 246478
rect 7918 246242 8002 246478
rect 8238 246242 8322 246478
rect 8558 246242 8642 246478
rect 8878 246242 226838 246478
rect 227074 246242 227158 246478
rect 227394 246242 227478 246478
rect 227714 246242 227798 246478
rect 228034 246242 228118 246478
rect 228354 246242 228438 246478
rect 228674 246242 228758 246478
rect 228994 246242 229078 246478
rect 229314 246242 229398 246478
rect 229634 246242 229718 246478
rect 229954 246242 230038 246478
rect 230274 246242 230358 246478
rect 230594 246242 230716 246478
rect 5000 246158 230716 246242
rect 5000 245922 5122 246158
rect 5358 245922 5442 246158
rect 5678 245922 5762 246158
rect 5998 245922 6082 246158
rect 6318 245922 6402 246158
rect 6638 245922 6722 246158
rect 6958 245922 7042 246158
rect 7278 245922 7362 246158
rect 7598 245922 7682 246158
rect 7918 245922 8002 246158
rect 8238 245922 8322 246158
rect 8558 245922 8642 246158
rect 8878 245922 226838 246158
rect 227074 245922 227158 246158
rect 227394 245922 227478 246158
rect 227714 245922 227798 246158
rect 228034 245922 228118 246158
rect 228354 245922 228438 246158
rect 228674 245922 228758 246158
rect 228994 245922 229078 246158
rect 229314 245922 229398 246158
rect 229634 245922 229718 246158
rect 229954 245922 230038 246158
rect 230274 245922 230358 246158
rect 230594 245922 230716 246158
rect 5000 245838 230716 245922
rect 5000 245602 5122 245838
rect 5358 245602 5442 245838
rect 5678 245602 5762 245838
rect 5998 245602 6082 245838
rect 6318 245602 6402 245838
rect 6638 245602 6722 245838
rect 6958 245602 7042 245838
rect 7278 245602 7362 245838
rect 7598 245602 7682 245838
rect 7918 245602 8002 245838
rect 8238 245602 8322 245838
rect 8558 245602 8642 245838
rect 8878 245602 226838 245838
rect 227074 245602 227158 245838
rect 227394 245602 227478 245838
rect 227714 245602 227798 245838
rect 228034 245602 228118 245838
rect 228354 245602 228438 245838
rect 228674 245602 228758 245838
rect 228994 245602 229078 245838
rect 229314 245602 229398 245838
rect 229634 245602 229718 245838
rect 229954 245602 230038 245838
rect 230274 245602 230358 245838
rect 230594 245602 230716 245838
rect 5000 245518 230716 245602
rect 5000 245282 5122 245518
rect 5358 245282 5442 245518
rect 5678 245282 5762 245518
rect 5998 245282 6082 245518
rect 6318 245282 6402 245518
rect 6638 245282 6722 245518
rect 6958 245282 7042 245518
rect 7278 245282 7362 245518
rect 7598 245282 7682 245518
rect 7918 245282 8002 245518
rect 8238 245282 8322 245518
rect 8558 245282 8642 245518
rect 8878 245282 226838 245518
rect 227074 245282 227158 245518
rect 227394 245282 227478 245518
rect 227714 245282 227798 245518
rect 228034 245282 228118 245518
rect 228354 245282 228438 245518
rect 228674 245282 228758 245518
rect 228994 245282 229078 245518
rect 229314 245282 229398 245518
rect 229634 245282 229718 245518
rect 229954 245282 230038 245518
rect 230274 245282 230358 245518
rect 230594 245282 230716 245518
rect 5000 245198 230716 245282
rect 5000 244962 5122 245198
rect 5358 244962 5442 245198
rect 5678 244962 5762 245198
rect 5998 244962 6082 245198
rect 6318 244962 6402 245198
rect 6638 244962 6722 245198
rect 6958 244962 7042 245198
rect 7278 244962 7362 245198
rect 7598 244962 7682 245198
rect 7918 244962 8002 245198
rect 8238 244962 8322 245198
rect 8558 244962 8642 245198
rect 8878 244962 226838 245198
rect 227074 244962 227158 245198
rect 227394 244962 227478 245198
rect 227714 244962 227798 245198
rect 228034 244962 228118 245198
rect 228354 244962 228438 245198
rect 228674 244962 228758 245198
rect 228994 244962 229078 245198
rect 229314 244962 229398 245198
rect 229634 244962 229718 245198
rect 229954 244962 230038 245198
rect 230274 244962 230358 245198
rect 230594 244962 230716 245198
rect 5000 244878 230716 244962
rect 5000 244642 5122 244878
rect 5358 244642 5442 244878
rect 5678 244642 5762 244878
rect 5998 244642 6082 244878
rect 6318 244642 6402 244878
rect 6638 244642 6722 244878
rect 6958 244642 7042 244878
rect 7278 244642 7362 244878
rect 7598 244642 7682 244878
rect 7918 244642 8002 244878
rect 8238 244642 8322 244878
rect 8558 244642 8642 244878
rect 8878 244642 226838 244878
rect 227074 244642 227158 244878
rect 227394 244642 227478 244878
rect 227714 244642 227798 244878
rect 228034 244642 228118 244878
rect 228354 244642 228438 244878
rect 228674 244642 228758 244878
rect 228994 244642 229078 244878
rect 229314 244642 229398 244878
rect 229634 244642 229718 244878
rect 229954 244642 230038 244878
rect 230274 244642 230358 244878
rect 230594 244642 230716 244878
rect 5000 244558 230716 244642
rect 5000 244322 5122 244558
rect 5358 244322 5442 244558
rect 5678 244322 5762 244558
rect 5998 244322 6082 244558
rect 6318 244322 6402 244558
rect 6638 244322 6722 244558
rect 6958 244322 7042 244558
rect 7278 244322 7362 244558
rect 7598 244322 7682 244558
rect 7918 244322 8002 244558
rect 8238 244322 8322 244558
rect 8558 244322 8642 244558
rect 8878 244322 226838 244558
rect 227074 244322 227158 244558
rect 227394 244322 227478 244558
rect 227714 244322 227798 244558
rect 228034 244322 228118 244558
rect 228354 244322 228438 244558
rect 228674 244322 228758 244558
rect 228994 244322 229078 244558
rect 229314 244322 229398 244558
rect 229634 244322 229718 244558
rect 229954 244322 230038 244558
rect 230274 244322 230358 244558
rect 230594 244322 230716 244558
rect 5000 244200 230716 244322
rect 0 240118 235716 240160
rect 0 239882 5122 240118
rect 5358 239882 5442 240118
rect 5678 239882 5762 240118
rect 5998 239882 6082 240118
rect 6318 239882 6402 240118
rect 6638 239882 6722 240118
rect 6958 239882 7042 240118
rect 7278 239882 7362 240118
rect 7598 239882 7682 240118
rect 7918 239882 8002 240118
rect 8238 239882 8322 240118
rect 8558 239882 8642 240118
rect 8878 239882 226838 240118
rect 227074 239882 227158 240118
rect 227394 239882 227478 240118
rect 227714 239882 227798 240118
rect 228034 239882 228118 240118
rect 228354 239882 228438 240118
rect 228674 239882 228758 240118
rect 228994 239882 229078 240118
rect 229314 239882 229398 240118
rect 229634 239882 229718 240118
rect 229954 239882 230038 240118
rect 230274 239882 230358 240118
rect 230594 239882 235716 240118
rect 0 239840 235716 239882
rect 0 228918 235716 228960
rect 0 228682 122 228918
rect 358 228682 442 228918
rect 678 228682 762 228918
rect 998 228682 1082 228918
rect 1318 228682 1402 228918
rect 1638 228682 1722 228918
rect 1958 228682 2042 228918
rect 2278 228682 2362 228918
rect 2598 228682 2682 228918
rect 2918 228682 3002 228918
rect 3238 228682 3322 228918
rect 3558 228682 3642 228918
rect 3878 228682 30215 228918
rect 30451 228682 71882 228918
rect 72118 228682 114215 228918
rect 114451 228682 155882 228918
rect 156118 228682 198215 228918
rect 198451 228682 231838 228918
rect 232074 228682 232158 228918
rect 232394 228682 232478 228918
rect 232714 228682 232798 228918
rect 233034 228682 233118 228918
rect 233354 228682 233438 228918
rect 233674 228682 233758 228918
rect 233994 228682 234078 228918
rect 234314 228682 234398 228918
rect 234634 228682 234718 228918
rect 234954 228682 235038 228918
rect 235274 228682 235358 228918
rect 235594 228682 235716 228918
rect 0 228640 235716 228682
rect 0 217718 235716 217760
rect 0 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 25549 217718
rect 25785 217482 66882 217718
rect 67118 217482 109549 217718
rect 109785 217482 150882 217718
rect 151118 217482 193549 217718
rect 193785 217482 226838 217718
rect 227074 217482 227158 217718
rect 227394 217482 227478 217718
rect 227714 217482 227798 217718
rect 228034 217482 228118 217718
rect 228354 217482 228438 217718
rect 228674 217482 228758 217718
rect 228994 217482 229078 217718
rect 229314 217482 229398 217718
rect 229634 217482 229718 217718
rect 229954 217482 230038 217718
rect 230274 217482 230358 217718
rect 230594 217482 235716 217718
rect 0 217440 235716 217482
rect 0 206518 235716 206560
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 231838 206518
rect 232074 206282 232158 206518
rect 232394 206282 232478 206518
rect 232714 206282 232798 206518
rect 233034 206282 233118 206518
rect 233354 206282 233438 206518
rect 233674 206282 233758 206518
rect 233994 206282 234078 206518
rect 234314 206282 234398 206518
rect 234634 206282 234718 206518
rect 234954 206282 235038 206518
rect 235274 206282 235358 206518
rect 235594 206282 235716 206518
rect 0 206240 235716 206282
rect 0 195318 235716 195360
rect 0 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 226838 195318
rect 227074 195082 227158 195318
rect 227394 195082 227478 195318
rect 227714 195082 227798 195318
rect 228034 195082 228118 195318
rect 228354 195082 228438 195318
rect 228674 195082 228758 195318
rect 228994 195082 229078 195318
rect 229314 195082 229398 195318
rect 229634 195082 229718 195318
rect 229954 195082 230038 195318
rect 230274 195082 230358 195318
rect 230594 195082 235716 195318
rect 0 195040 235716 195082
rect 193828 190842 210156 190884
rect 193828 190606 193870 190842
rect 194106 190606 209878 190842
rect 210114 190606 210156 190842
rect 193828 190564 210156 190606
rect 0 184118 235716 184160
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 32215 184118
rect 32451 183882 75506 184118
rect 75742 183882 116215 184118
rect 116451 183882 159506 184118
rect 159742 183882 200215 184118
rect 200451 183882 231838 184118
rect 232074 183882 232158 184118
rect 232394 183882 232478 184118
rect 232714 183882 232798 184118
rect 233034 183882 233118 184118
rect 233354 183882 233438 184118
rect 233674 183882 233758 184118
rect 233994 183882 234078 184118
rect 234314 183882 234398 184118
rect 234634 183882 234718 184118
rect 234954 183882 235038 184118
rect 235274 183882 235358 184118
rect 235594 183882 235716 184118
rect 0 183840 235716 183882
rect 0 172918 235716 172960
rect 0 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 29549 172918
rect 29785 172682 60146 172918
rect 60382 172682 113549 172918
rect 113785 172682 144146 172918
rect 144382 172682 197549 172918
rect 197785 172682 226838 172918
rect 227074 172682 227158 172918
rect 227394 172682 227478 172918
rect 227714 172682 227798 172918
rect 228034 172682 228118 172918
rect 228354 172682 228438 172918
rect 228674 172682 228758 172918
rect 228994 172682 229078 172918
rect 229314 172682 229398 172918
rect 229634 172682 229718 172918
rect 229954 172682 230038 172918
rect 230274 172682 230358 172918
rect 230594 172682 235716 172918
rect 0 172640 235716 172682
rect 0 161718 235716 161760
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 32215 161718
rect 32451 161482 75506 161718
rect 75742 161482 116215 161718
rect 116451 161482 159506 161718
rect 159742 161482 200215 161718
rect 200451 161482 231838 161718
rect 232074 161482 232158 161718
rect 232394 161482 232478 161718
rect 232714 161482 232798 161718
rect 233034 161482 233118 161718
rect 233354 161482 233438 161718
rect 233674 161482 233758 161718
rect 233994 161482 234078 161718
rect 234314 161482 234398 161718
rect 234634 161482 234718 161718
rect 234954 161482 235038 161718
rect 235274 161482 235358 161718
rect 235594 161482 235716 161718
rect 0 161440 235716 161482
rect 137892 156842 209972 156884
rect 137892 156606 137934 156842
rect 138170 156606 209694 156842
rect 209930 156606 209972 156842
rect 137892 156564 209972 156606
rect 0 150518 235716 150560
rect 0 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 226838 150518
rect 227074 150282 227158 150518
rect 227394 150282 227478 150518
rect 227714 150282 227798 150518
rect 228034 150282 228118 150518
rect 228354 150282 228438 150518
rect 228674 150282 228758 150518
rect 228994 150282 229078 150518
rect 229314 150282 229398 150518
rect 229634 150282 229718 150518
rect 229954 150282 230038 150518
rect 230274 150282 230358 150518
rect 230594 150282 235716 150518
rect 0 150240 235716 150282
rect 0 139318 235716 139360
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 231838 139318
rect 232074 139082 232158 139318
rect 232394 139082 232478 139318
rect 232714 139082 232798 139318
rect 233034 139082 233118 139318
rect 233354 139082 233438 139318
rect 233674 139082 233758 139318
rect 233994 139082 234078 139318
rect 234314 139082 234398 139318
rect 234634 139082 234718 139318
rect 234954 139082 235038 139318
rect 235274 139082 235358 139318
rect 235594 139082 235716 139318
rect 0 139040 235716 139082
rect 0 128118 235716 128160
rect 0 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 25549 128118
rect 25785 127882 66882 128118
rect 67118 127882 109549 128118
rect 109785 127882 150882 128118
rect 151118 127882 193549 128118
rect 193785 127882 226838 128118
rect 227074 127882 227158 128118
rect 227394 127882 227478 128118
rect 227714 127882 227798 128118
rect 228034 127882 228118 128118
rect 228354 127882 228438 128118
rect 228674 127882 228758 128118
rect 228994 127882 229078 128118
rect 229314 127882 229398 128118
rect 229634 127882 229718 128118
rect 229954 127882 230038 128118
rect 230274 127882 230358 128118
rect 230594 127882 235716 128118
rect 0 127840 235716 127882
rect 0 116918 235716 116960
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 30215 116918
rect 30451 116682 114215 116918
rect 114451 116682 198215 116918
rect 198451 116682 231838 116918
rect 232074 116682 232158 116918
rect 232394 116682 232478 116918
rect 232714 116682 232798 116918
rect 233034 116682 233118 116918
rect 233354 116682 233438 116918
rect 233674 116682 233758 116918
rect 233994 116682 234078 116918
rect 234314 116682 234398 116918
rect 234634 116682 234718 116918
rect 234954 116682 235038 116918
rect 235274 116682 235358 116918
rect 235594 116682 235716 116918
rect 0 116640 235716 116682
rect 0 105718 235716 105760
rect 0 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 226838 105718
rect 227074 105482 227158 105718
rect 227394 105482 227478 105718
rect 227714 105482 227798 105718
rect 228034 105482 228118 105718
rect 228354 105482 228438 105718
rect 228674 105482 228758 105718
rect 228994 105482 229078 105718
rect 229314 105482 229398 105718
rect 229634 105482 229718 105718
rect 229954 105482 230038 105718
rect 230274 105482 230358 105718
rect 230594 105482 235716 105718
rect 0 105440 235716 105482
rect 193644 97002 209972 97044
rect 193644 96766 193686 97002
rect 193922 96766 209694 97002
rect 209930 96766 209972 97002
rect 193644 96724 209972 96766
rect 0 94518 235716 94560
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 32215 94518
rect 32451 94282 75506 94518
rect 75742 94282 116215 94518
rect 116451 94282 159506 94518
rect 159742 94282 200215 94518
rect 200451 94282 231838 94518
rect 232074 94282 232158 94518
rect 232394 94282 232478 94518
rect 232714 94282 232798 94518
rect 233034 94282 233118 94518
rect 233354 94282 233438 94518
rect 233674 94282 233758 94518
rect 233994 94282 234078 94518
rect 234314 94282 234398 94518
rect 234634 94282 234718 94518
rect 234954 94282 235038 94518
rect 235274 94282 235358 94518
rect 235594 94282 235716 94518
rect 0 94240 235716 94282
rect 0 83318 235716 83360
rect 0 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 29549 83318
rect 29785 83082 60146 83318
rect 60382 83082 113549 83318
rect 113785 83082 144146 83318
rect 144382 83082 197549 83318
rect 197785 83082 226838 83318
rect 227074 83082 227158 83318
rect 227394 83082 227478 83318
rect 227714 83082 227798 83318
rect 228034 83082 228118 83318
rect 228354 83082 228438 83318
rect 228674 83082 228758 83318
rect 228994 83082 229078 83318
rect 229314 83082 229398 83318
rect 229634 83082 229718 83318
rect 229954 83082 230038 83318
rect 230274 83082 230358 83318
rect 230594 83082 235716 83318
rect 0 83040 235716 83082
rect 0 72118 235716 72160
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 32215 72118
rect 32451 71882 75506 72118
rect 75742 71882 116215 72118
rect 116451 71882 159506 72118
rect 159742 71882 200215 72118
rect 200451 71882 231838 72118
rect 232074 71882 232158 72118
rect 232394 71882 232478 72118
rect 232714 71882 232798 72118
rect 233034 71882 233118 72118
rect 233354 71882 233438 72118
rect 233674 71882 233758 72118
rect 233994 71882 234078 72118
rect 234314 71882 234398 72118
rect 234634 71882 234718 72118
rect 234954 71882 235038 72118
rect 235274 71882 235358 72118
rect 235594 71882 235716 72118
rect 0 71840 235716 71882
rect 13140 67082 56148 67124
rect 13140 66846 13182 67082
rect 13418 66846 55870 67082
rect 56106 66846 56148 67082
rect 13140 66804 56148 66846
rect 0 60918 235716 60960
rect 0 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 226838 60918
rect 227074 60682 227158 60918
rect 227394 60682 227478 60918
rect 227714 60682 227798 60918
rect 228034 60682 228118 60918
rect 228354 60682 228438 60918
rect 228674 60682 228758 60918
rect 228994 60682 229078 60918
rect 229314 60682 229398 60918
rect 229634 60682 229718 60918
rect 229954 60682 230038 60918
rect 230274 60682 230358 60918
rect 230594 60682 235716 60918
rect 0 60640 235716 60682
rect 0 49718 235716 49760
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 231838 49718
rect 232074 49482 232158 49718
rect 232394 49482 232478 49718
rect 232714 49482 232798 49718
rect 233034 49482 233118 49718
rect 233354 49482 233438 49718
rect 233674 49482 233758 49718
rect 233994 49482 234078 49718
rect 234314 49482 234398 49718
rect 234634 49482 234718 49718
rect 234954 49482 235038 49718
rect 235274 49482 235358 49718
rect 235594 49482 235716 49718
rect 0 49440 235716 49482
rect 151876 43282 155140 43324
rect 151876 43046 154862 43282
rect 155098 43046 155140 43282
rect 151876 43004 155140 43046
rect 159420 43282 159740 43324
rect 159420 43046 159462 43282
rect 159698 43046 159740 43282
rect 151876 40604 152196 43004
rect 159420 40604 159740 43046
rect 151508 40562 152196 40604
rect 151508 40326 151550 40562
rect 151786 40326 152196 40562
rect 151508 40284 152196 40326
rect 152612 40284 159740 40604
rect 152612 39924 152932 40284
rect 150404 39882 152932 39924
rect 150404 39646 150446 39882
rect 150682 39646 152932 39882
rect 150404 39604 152932 39646
rect 0 38518 235716 38560
rect 0 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 25549 38518
rect 25785 38282 66882 38518
rect 67118 38282 109549 38518
rect 109785 38282 150882 38518
rect 151118 38282 193549 38518
rect 193785 38282 226838 38518
rect 227074 38282 227158 38518
rect 227394 38282 227478 38518
rect 227714 38282 227798 38518
rect 228034 38282 228118 38518
rect 228354 38282 228438 38518
rect 228674 38282 228758 38518
rect 228994 38282 229078 38518
rect 229314 38282 229398 38518
rect 229634 38282 229718 38518
rect 229954 38282 230038 38518
rect 230274 38282 230358 38518
rect 230594 38282 235716 38518
rect 0 38240 235716 38282
rect 211860 35802 212916 35844
rect 211860 35566 212638 35802
rect 212874 35566 212916 35802
rect 211860 35524 212916 35566
rect 211860 35164 212180 35524
rect 211860 35122 212916 35164
rect 211860 34886 212638 35122
rect 212874 34886 212916 35122
rect 211860 34844 212916 34886
rect 0 27318 235716 27360
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 30215 27318
rect 30451 27082 71882 27318
rect 72118 27082 114215 27318
rect 114451 27082 155882 27318
rect 156118 27082 198215 27318
rect 198451 27082 231838 27318
rect 232074 27082 232158 27318
rect 232394 27082 232478 27318
rect 232714 27082 232798 27318
rect 233034 27082 233118 27318
rect 233354 27082 233438 27318
rect 233674 27082 233758 27318
rect 233994 27082 234078 27318
rect 234314 27082 234398 27318
rect 234634 27082 234718 27318
rect 234954 27082 235038 27318
rect 235274 27082 235358 27318
rect 235594 27082 235716 27318
rect 0 27040 235716 27082
rect 212412 25602 212916 25644
rect 212412 25366 212638 25602
rect 212874 25366 212916 25602
rect 212412 25324 212916 25366
rect 212412 24964 212732 25324
rect 212412 24922 212916 24964
rect 212412 24686 212638 24922
rect 212874 24686 212916 24922
rect 212412 24644 212916 24686
rect 150404 22202 156244 22244
rect 150404 21966 150446 22202
rect 150682 21966 155966 22202
rect 156202 21966 156244 22202
rect 150404 21924 156244 21966
rect 173772 22202 185316 22244
rect 173772 21966 173814 22202
rect 174050 21966 185038 22202
rect 185274 21966 185316 22202
rect 173772 21924 185316 21966
rect 212596 21522 222484 21564
rect 212596 21286 212638 21522
rect 212874 21286 222206 21522
rect 222442 21286 222484 21522
rect 212596 21244 222484 21286
rect 88948 20842 101780 20884
rect 88948 20606 88990 20842
rect 89226 20606 101502 20842
rect 101738 20606 101780 20842
rect 88948 20564 101780 20606
rect 173036 20842 185316 20884
rect 173036 20606 173078 20842
rect 173314 20606 185038 20842
rect 185274 20606 185316 20842
rect 173036 20564 185316 20606
rect 89684 20162 101780 20204
rect 89684 19926 89726 20162
rect 89962 19926 101502 20162
rect 101738 19926 101780 20162
rect 89684 19884 101780 19926
rect 173404 20162 185684 20204
rect 173404 19926 173446 20162
rect 173682 19926 185406 20162
rect 185642 19926 185684 20162
rect 173404 19884 185684 19926
rect 0 16118 235716 16160
rect 0 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 226838 16118
rect 227074 15882 227158 16118
rect 227394 15882 227478 16118
rect 227714 15882 227798 16118
rect 228034 15882 228118 16118
rect 228354 15882 228438 16118
rect 228674 15882 228758 16118
rect 228994 15882 229078 16118
rect 229314 15882 229398 16118
rect 229634 15882 229718 16118
rect 229954 15882 230038 16118
rect 230274 15882 230358 16118
rect 230594 15882 235716 16118
rect 0 15840 235716 15882
rect 5000 8878 230716 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 226838 8878
rect 227074 8642 227158 8878
rect 227394 8642 227478 8878
rect 227714 8642 227798 8878
rect 228034 8642 228118 8878
rect 228354 8642 228438 8878
rect 228674 8642 228758 8878
rect 228994 8642 229078 8878
rect 229314 8642 229398 8878
rect 229634 8642 229718 8878
rect 229954 8642 230038 8878
rect 230274 8642 230358 8878
rect 230594 8642 230716 8878
rect 5000 8558 230716 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 226838 8558
rect 227074 8322 227158 8558
rect 227394 8322 227478 8558
rect 227714 8322 227798 8558
rect 228034 8322 228118 8558
rect 228354 8322 228438 8558
rect 228674 8322 228758 8558
rect 228994 8322 229078 8558
rect 229314 8322 229398 8558
rect 229634 8322 229718 8558
rect 229954 8322 230038 8558
rect 230274 8322 230358 8558
rect 230594 8322 230716 8558
rect 5000 8238 230716 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 226838 8238
rect 227074 8002 227158 8238
rect 227394 8002 227478 8238
rect 227714 8002 227798 8238
rect 228034 8002 228118 8238
rect 228354 8002 228438 8238
rect 228674 8002 228758 8238
rect 228994 8002 229078 8238
rect 229314 8002 229398 8238
rect 229634 8002 229718 8238
rect 229954 8002 230038 8238
rect 230274 8002 230358 8238
rect 230594 8002 230716 8238
rect 5000 7918 230716 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 226838 7918
rect 227074 7682 227158 7918
rect 227394 7682 227478 7918
rect 227714 7682 227798 7918
rect 228034 7682 228118 7918
rect 228354 7682 228438 7918
rect 228674 7682 228758 7918
rect 228994 7682 229078 7918
rect 229314 7682 229398 7918
rect 229634 7682 229718 7918
rect 229954 7682 230038 7918
rect 230274 7682 230358 7918
rect 230594 7682 230716 7918
rect 5000 7598 230716 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 226838 7598
rect 227074 7362 227158 7598
rect 227394 7362 227478 7598
rect 227714 7362 227798 7598
rect 228034 7362 228118 7598
rect 228354 7362 228438 7598
rect 228674 7362 228758 7598
rect 228994 7362 229078 7598
rect 229314 7362 229398 7598
rect 229634 7362 229718 7598
rect 229954 7362 230038 7598
rect 230274 7362 230358 7598
rect 230594 7362 230716 7598
rect 5000 7278 230716 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 226838 7278
rect 227074 7042 227158 7278
rect 227394 7042 227478 7278
rect 227714 7042 227798 7278
rect 228034 7042 228118 7278
rect 228354 7042 228438 7278
rect 228674 7042 228758 7278
rect 228994 7042 229078 7278
rect 229314 7042 229398 7278
rect 229634 7042 229718 7278
rect 229954 7042 230038 7278
rect 230274 7042 230358 7278
rect 230594 7042 230716 7278
rect 5000 6958 230716 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 226838 6958
rect 227074 6722 227158 6958
rect 227394 6722 227478 6958
rect 227714 6722 227798 6958
rect 228034 6722 228118 6958
rect 228354 6722 228438 6958
rect 228674 6722 228758 6958
rect 228994 6722 229078 6958
rect 229314 6722 229398 6958
rect 229634 6722 229718 6958
rect 229954 6722 230038 6958
rect 230274 6722 230358 6958
rect 230594 6722 230716 6958
rect 5000 6638 230716 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 226838 6638
rect 227074 6402 227158 6638
rect 227394 6402 227478 6638
rect 227714 6402 227798 6638
rect 228034 6402 228118 6638
rect 228354 6402 228438 6638
rect 228674 6402 228758 6638
rect 228994 6402 229078 6638
rect 229314 6402 229398 6638
rect 229634 6402 229718 6638
rect 229954 6402 230038 6638
rect 230274 6402 230358 6638
rect 230594 6402 230716 6638
rect 5000 6318 230716 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 226838 6318
rect 227074 6082 227158 6318
rect 227394 6082 227478 6318
rect 227714 6082 227798 6318
rect 228034 6082 228118 6318
rect 228354 6082 228438 6318
rect 228674 6082 228758 6318
rect 228994 6082 229078 6318
rect 229314 6082 229398 6318
rect 229634 6082 229718 6318
rect 229954 6082 230038 6318
rect 230274 6082 230358 6318
rect 230594 6082 230716 6318
rect 5000 5998 230716 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 226838 5998
rect 227074 5762 227158 5998
rect 227394 5762 227478 5998
rect 227714 5762 227798 5998
rect 228034 5762 228118 5998
rect 228354 5762 228438 5998
rect 228674 5762 228758 5998
rect 228994 5762 229078 5998
rect 229314 5762 229398 5998
rect 229634 5762 229718 5998
rect 229954 5762 230038 5998
rect 230274 5762 230358 5998
rect 230594 5762 230716 5998
rect 5000 5678 230716 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 226838 5678
rect 227074 5442 227158 5678
rect 227394 5442 227478 5678
rect 227714 5442 227798 5678
rect 228034 5442 228118 5678
rect 228354 5442 228438 5678
rect 228674 5442 228758 5678
rect 228994 5442 229078 5678
rect 229314 5442 229398 5678
rect 229634 5442 229718 5678
rect 229954 5442 230038 5678
rect 230274 5442 230358 5678
rect 230594 5442 230716 5678
rect 5000 5358 230716 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 226838 5358
rect 227074 5122 227158 5358
rect 227394 5122 227478 5358
rect 227714 5122 227798 5358
rect 228034 5122 228118 5358
rect 228354 5122 228438 5358
rect 228674 5122 228758 5358
rect 228994 5122 229078 5358
rect 229314 5122 229398 5358
rect 229634 5122 229718 5358
rect 229954 5122 230038 5358
rect 230274 5122 230358 5358
rect 230594 5122 230716 5358
rect 5000 5000 230716 5122
rect 0 3878 235716 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 231838 3878
rect 232074 3642 232158 3878
rect 232394 3642 232478 3878
rect 232714 3642 232798 3878
rect 233034 3642 233118 3878
rect 233354 3642 233438 3878
rect 233674 3642 233758 3878
rect 233994 3642 234078 3878
rect 234314 3642 234398 3878
rect 234634 3642 234718 3878
rect 234954 3642 235038 3878
rect 235274 3642 235358 3878
rect 235594 3642 235716 3878
rect 0 3558 235716 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 231838 3558
rect 232074 3322 232158 3558
rect 232394 3322 232478 3558
rect 232714 3322 232798 3558
rect 233034 3322 233118 3558
rect 233354 3322 233438 3558
rect 233674 3322 233758 3558
rect 233994 3322 234078 3558
rect 234314 3322 234398 3558
rect 234634 3322 234718 3558
rect 234954 3322 235038 3558
rect 235274 3322 235358 3558
rect 235594 3322 235716 3558
rect 0 3238 235716 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 231838 3238
rect 232074 3002 232158 3238
rect 232394 3002 232478 3238
rect 232714 3002 232798 3238
rect 233034 3002 233118 3238
rect 233354 3002 233438 3238
rect 233674 3002 233758 3238
rect 233994 3002 234078 3238
rect 234314 3002 234398 3238
rect 234634 3002 234718 3238
rect 234954 3002 235038 3238
rect 235274 3002 235358 3238
rect 235594 3002 235716 3238
rect 0 2918 235716 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 231838 2918
rect 232074 2682 232158 2918
rect 232394 2682 232478 2918
rect 232714 2682 232798 2918
rect 233034 2682 233118 2918
rect 233354 2682 233438 2918
rect 233674 2682 233758 2918
rect 233994 2682 234078 2918
rect 234314 2682 234398 2918
rect 234634 2682 234718 2918
rect 234954 2682 235038 2918
rect 235274 2682 235358 2918
rect 235594 2682 235716 2918
rect 0 2598 235716 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 231838 2598
rect 232074 2362 232158 2598
rect 232394 2362 232478 2598
rect 232714 2362 232798 2598
rect 233034 2362 233118 2598
rect 233354 2362 233438 2598
rect 233674 2362 233758 2598
rect 233994 2362 234078 2598
rect 234314 2362 234398 2598
rect 234634 2362 234718 2598
rect 234954 2362 235038 2598
rect 235274 2362 235358 2598
rect 235594 2362 235716 2598
rect 0 2278 235716 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 231838 2278
rect 232074 2042 232158 2278
rect 232394 2042 232478 2278
rect 232714 2042 232798 2278
rect 233034 2042 233118 2278
rect 233354 2042 233438 2278
rect 233674 2042 233758 2278
rect 233994 2042 234078 2278
rect 234314 2042 234398 2278
rect 234634 2042 234718 2278
rect 234954 2042 235038 2278
rect 235274 2042 235358 2278
rect 235594 2042 235716 2278
rect 0 1958 235716 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 231838 1958
rect 232074 1722 232158 1958
rect 232394 1722 232478 1958
rect 232714 1722 232798 1958
rect 233034 1722 233118 1958
rect 233354 1722 233438 1958
rect 233674 1722 233758 1958
rect 233994 1722 234078 1958
rect 234314 1722 234398 1958
rect 234634 1722 234718 1958
rect 234954 1722 235038 1958
rect 235274 1722 235358 1958
rect 235594 1722 235716 1958
rect 0 1638 235716 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 231838 1638
rect 232074 1402 232158 1638
rect 232394 1402 232478 1638
rect 232714 1402 232798 1638
rect 233034 1402 233118 1638
rect 233354 1402 233438 1638
rect 233674 1402 233758 1638
rect 233994 1402 234078 1638
rect 234314 1402 234398 1638
rect 234634 1402 234718 1638
rect 234954 1402 235038 1638
rect 235274 1402 235358 1638
rect 235594 1402 235716 1638
rect 0 1318 235716 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 231838 1318
rect 232074 1082 232158 1318
rect 232394 1082 232478 1318
rect 232714 1082 232798 1318
rect 233034 1082 233118 1318
rect 233354 1082 233438 1318
rect 233674 1082 233758 1318
rect 233994 1082 234078 1318
rect 234314 1082 234398 1318
rect 234634 1082 234718 1318
rect 234954 1082 235038 1318
rect 235274 1082 235358 1318
rect 235594 1082 235716 1318
rect 0 998 235716 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 231838 998
rect 232074 762 232158 998
rect 232394 762 232478 998
rect 232714 762 232798 998
rect 233034 762 233118 998
rect 233354 762 233438 998
rect 233674 762 233758 998
rect 233994 762 234078 998
rect 234314 762 234398 998
rect 234634 762 234718 998
rect 234954 762 235038 998
rect 235274 762 235358 998
rect 235594 762 235716 998
rect 0 678 235716 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 231838 678
rect 232074 442 232158 678
rect 232394 442 232478 678
rect 232714 442 232798 678
rect 233034 442 233118 678
rect 233354 442 233438 678
rect 233674 442 233758 678
rect 233994 442 234078 678
rect 234314 442 234398 678
rect 234634 442 234718 678
rect 234954 442 235038 678
rect 235274 442 235358 678
rect 235594 442 235716 678
rect 0 358 235716 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 231838 358
rect 232074 122 232158 358
rect 232394 122 232478 358
rect 232714 122 232798 358
rect 233034 122 233118 358
rect 233354 122 233438 358
rect 233674 122 233758 358
rect 233994 122 234078 358
rect 234314 122 234398 358
rect 234634 122 234718 358
rect 234954 122 235038 358
rect 235274 122 235358 358
rect 235594 122 235716 358
rect 0 0 235716 122
use grid_clb  grid_clb_1__1_
timestamp 1605114789
transform 1 0 55896 0 1 59824
box 0 0 40000 40000
use sb_0__0_  sb_0__0_
timestamp 1605114789
transform 1 0 19896 0 1 18824
box 0 0 28000 27720
use cby_0__1_  cby_0__1_
timestamp 1605114789
transform 1 0 25896 0 1 59824
box 0 0 16000 40000
use cbx_1__0_  cbx_1__0_
timestamp 1605114789
transform 1 0 60896 0 1 20824
box 0 0 30000 24000
use grid_clb  grid_clb_2__1_
timestamp 1605114789
transform 1 0 139896 0 1 59824
box 0 0 40000 40000
use sb_1__0_  sb_1__0_
timestamp 1605114789
transform 1 0 103896 0 1 18824
box 0 0 28000 28000
use cby_1__1_  cby_1__1_
timestamp 1605114789
transform 1 0 109896 0 1 59824
box 0 0 16000 40000
use cbx_1__0_  cbx_2__0_
timestamp 1605114789
transform 1 0 144896 0 1 20824
box 0 0 30000 24000
use sb_2__0_  sb_2__0_
timestamp 1605114789
transform 1 0 187896 0 1 18824
box 0 0 28000 28000
use cby_2__1_  cby_2__1_
timestamp 1605114789
transform 1 0 193896 0 1 59824
box 0 0 16000 40000
use sb_0__1_  sb_0__1_
timestamp 1605114789
transform 1 0 19896 0 1 112824
box 0 0 28000 28000
use cbx_1__1_  cbx_1__1_
timestamp 1605114789
transform 1 0 60896 0 1 114824
box 0 0 30000 24000
use sb_1__1_  sb_1__1_
timestamp 1605114789
transform 1 0 103896 0 1 112824
box 0 0 28000 28000
use cbx_1__1_  cbx_2__1_
timestamp 1605114789
transform 1 0 144896 0 1 114824
box 0 0 30000 24000
use sb_2__1_  sb_2__1_
timestamp 1605114789
transform 1 0 187896 0 1 112824
box 0 0 28000 28000
use grid_clb  grid_clb_1__2_
timestamp 1605114789
transform 1 0 55896 0 1 153824
box 0 0 40000 40000
use cby_0__1_  cby_0__2_
timestamp 1605114789
transform 1 0 25896 0 1 153824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1605114789
transform 1 0 139896 0 1 153824
box 0 0 40000 40000
use cby_1__1_  cby_1__2_
timestamp 1605114789
transform 1 0 109896 0 1 153824
box 0 0 16000 40000
use cby_2__1_  cby_2__2_
timestamp 1605114789
transform 1 0 193896 0 1 153824
box 0 0 16000 40000
use sb_0__2_  sb_0__2_
timestamp 1605114789
transform 1 0 19896 0 1 206824
box 0 0 28000 28000
use cbx_1__2_  cbx_1__2_
timestamp 1605114789
transform 1 0 60896 0 1 208824
box 0 0 30000 24000
use sb_1__2_  sb_1__2_
timestamp 1605114789
transform 1 0 103896 0 1 206824
box 0 0 28000 28000
use cbx_1__2_  cbx_2__2_
timestamp 1605114789
transform 1 0 144896 0 1 208824
box 0 0 30000 24000
use sb_2__2_  sb_2__2_
timestamp 1605114789
transform 1 0 187896 0 1 206824
box 0 0 28000 28000
<< labels >>
rlabel metal3 s 9896 44056 10376 44176 6 Test_en
port 0 nsew default input
rlabel metal3 s 225416 205352 225896 205472 6 ccff_head
port 1 nsew default input
rlabel metal3 s 9896 20528 10376 20648 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 67720 10376 67840 6 clk
port 3 nsew default input
rlabel metal2 s 27854 244344 27910 244824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 4 nsew default tristate
rlabel metal2 s 120866 8824 120922 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
port 5 nsew default tristate
rlabel metal2 s 126846 8824 126902 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
port 6 nsew default tristate
rlabel metal2 s 132826 8824 132882 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
port 7 nsew default tristate
rlabel metal2 s 138806 8824 138862 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
port 8 nsew default tristate
rlabel metal2 s 144786 8824 144842 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
port 9 nsew default tristate
rlabel metal2 s 150858 8824 150914 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
port 10 nsew default tristate
rlabel metal3 s 9896 91248 10376 91368 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
port 11 nsew default tristate
rlabel metal3 s 9896 162104 10376 162224 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
port 12 nsew default tristate
rlabel metal2 s 63826 244344 63882 244824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 13 nsew default tristate
rlabel metal3 s 225416 48000 225896 48120 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 14 nsew default tristate
rlabel metal3 s 225416 126744 225896 126864 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 15 nsew default tristate
rlabel metal2 s 12858 8824 12914 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 16 nsew default tristate
rlabel metal2 s 18838 8824 18894 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 17 nsew default tristate
rlabel metal2 s 24818 8824 24874 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
port 18 nsew default tristate
rlabel metal2 s 30798 8824 30854 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
port 19 nsew default tristate
rlabel metal2 s 36778 8824 36834 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
port 20 nsew default tristate
rlabel metal2 s 42850 8824 42906 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
port 21 nsew default tristate
rlabel metal2 s 99798 244344 99854 244824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 22 nsew default input
rlabel metal2 s 156838 8824 156894 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[10]
port 23 nsew default input
rlabel metal2 s 162818 8824 162874 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[11]
port 24 nsew default input
rlabel metal2 s 168798 8824 168854 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[12]
port 25 nsew default input
rlabel metal2 s 174870 8824 174926 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[13]
port 26 nsew default input
rlabel metal2 s 180850 8824 180906 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[14]
port 27 nsew default input
rlabel metal2 s 186830 8824 186886 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[15]
port 28 nsew default input
rlabel metal3 s 9896 114912 10376 115032 6 gfpga_pad_EMBEDDED_IO_SOC_IN[16]
port 29 nsew default input
rlabel metal3 s 9896 185632 10376 185752 6 gfpga_pad_EMBEDDED_IO_SOC_IN[17]
port 30 nsew default input
rlabel metal2 s 135862 244344 135918 244824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 31 nsew default input
rlabel metal3 s 225416 74248 225896 74368 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 32 nsew default input
rlabel metal3 s 225416 152856 225896 152976 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 33 nsew default input
rlabel metal2 s 48830 8824 48886 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 34 nsew default input
rlabel metal2 s 54810 8824 54866 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 35 nsew default input
rlabel metal2 s 60790 8824 60846 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[6]
port 36 nsew default input
rlabel metal2 s 66862 8824 66918 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[7]
port 37 nsew default input
rlabel metal2 s 72842 8824 72898 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[8]
port 38 nsew default input
rlabel metal2 s 78822 8824 78878 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[9]
port 39 nsew default input
rlabel metal2 s 171834 244344 171890 244824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 40 nsew default tristate
rlabel metal2 s 192810 8824 192866 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
port 41 nsew default tristate
rlabel metal2 s 198790 8824 198846 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
port 42 nsew default tristate
rlabel metal2 s 204862 8824 204918 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
port 43 nsew default tristate
rlabel metal2 s 210842 8824 210898 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
port 44 nsew default tristate
rlabel metal2 s 216822 8824 216878 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
port 45 nsew default tristate
rlabel metal2 s 222802 8824 222858 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
port 46 nsew default tristate
rlabel metal3 s 9896 138440 10376 138560 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
port 47 nsew default tristate
rlabel metal3 s 9896 209296 10376 209416 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
port 48 nsew default tristate
rlabel metal2 s 207806 244344 207862 244824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 49 nsew default tristate
rlabel metal3 s 225416 100496 225896 100616 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 50 nsew default tristate
rlabel metal3 s 225416 179104 225896 179224 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 51 nsew default tristate
rlabel metal2 s 84802 8824 84858 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 52 nsew default tristate
rlabel metal2 s 90782 8824 90838 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 53 nsew default tristate
rlabel metal2 s 96854 8824 96910 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
port 54 nsew default tristate
rlabel metal2 s 102834 8824 102890 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
port 55 nsew default tristate
rlabel metal2 s 108814 8824 108870 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
port 56 nsew default tristate
rlabel metal2 s 114794 8824 114850 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
port 57 nsew default tristate
rlabel metal3 s 225416 21888 225896 22008 6 prog_clk
port 58 nsew default input
rlabel metal3 s 9896 232824 10376 232944 6 sc_head
port 59 nsew default input
rlabel metal3 s 225416 231600 225896 231720 6 sc_tail
port 60 nsew default tristate
rlabel metal5 s 5000 5000 230716 9000 8 VPWR
port 61 nsew default input
rlabel metal5 s 0 0 235716 4000 8 VGND
port 62 nsew default input
<< properties >>
string FIXED_BBOX 0 0 235716 253200
<< end >>
