* NGSPICE file created from sb_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_1__2_ SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP bottom_left_grid_pin_42_
+ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_
+ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11] chanx_right_in[12]
+ chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16] chanx_right_in[17]
+ chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3]
+ chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7] chanx_right_in[8]
+ chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11] chanx_right_out[12]
+ chanx_right_out[13] chanx_right_out[14] chanx_right_out[15] chanx_right_out[16]
+ chanx_right_out[17] chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11]
+ chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15]
+ chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0]
+ chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12] chany_bottom_out[13]
+ chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16] chany_bottom_out[17]
+ chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] left_bottom_grid_pin_34_
+ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_
+ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_ left_bottom_grid_pin_41_ left_top_grid_pin_1_
+ prog_clk right_bottom_grid_pin_34_ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_
+ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_
+ right_bottom_grid_pin_41_ right_top_grid_pin_1_ VPWR VGND
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_3.mux_l1_in_2_/S mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A0 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A1 mux_left_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_062_ _062_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__S mux_bottom_track_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__S mux_bottom_track_7.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_3__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_114_ _114_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l1_in_0_ bottom_left_grid_pin_46_ chanx_right_in[13] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l2_in_1__A1 mux_left_track_33.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_028_ _028_/HI _028_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_19.mux_l2_in_0_/S
+ mux_bottom_track_21.mux_l1_in_1_/S mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_16.mux_l3_in_0__S mux_right_track_16.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_19.mux_l2_in_0__S mux_bottom_track_19.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _117_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A1 mux_left_track_33.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_2__A0 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[4] mux_bottom_track_3.mux_l1_in_2_/S
+ mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0__A1 chanx_right_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/S mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A mux_left_track_1.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__A0 mux_left_track_9.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_061_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l2_in_2__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_5.mux_l2_in_1_/S
+ mux_bottom_track_5.mux_l3_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l4_in_0__A0 mux_left_track_9.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_113_ _113_/A chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_4.mux_l2_in_2__S mux_right_track_4.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.mux_l2_in_3_ _042_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _066_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_1__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l2_in_1__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_23.mux_l1_in_0__S mux_bottom_track_23.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/S mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_27.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__A1 mux_left_track_9.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_060_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A0 mux_right_track_4.mux_l1_in_5_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__061__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_5.mux_l1_in_3_/S
+ mux_bottom_track_5.mux_l2_in_1_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l4_in_0__A1 mux_left_track_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_112_ _112_/A chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__056__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A0 mux_right_track_4.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l2_in_1__S mux_left_track_25.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0__S mux_bottom_track_15.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A0 mux_right_track_4.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A0 mux_bottom_track_13.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__064__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_11.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__059__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A0 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_2__A1 mux_right_track_4.mux_l1_in_4_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_3_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_111_ _111_/A chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__072__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__A1 mux_right_track_4.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_2__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 mux_bottom_track_5.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__067__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A0 mux_bottom_track_21.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_1_ chany_bottom_in[9] chany_bottom_in[2] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l4_in_0__A1 mux_right_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0__A1 mux_bottom_track_13.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__080__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__075__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_110_ _110_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_21.mux_l1_in_1__A1 chanx_left_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_11.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l2_in_0_/S mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l3_in_0_/X
+ _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__083__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_21.mux_l2_in_0__A1 mux_bottom_track_21.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_41_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_24.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__078__A _078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_6__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__S mux_bottom_track_11.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__091__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_11.mux_l3_in_0_/S
+ mux_bottom_track_13.mux_l1_in_1_/S mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 chany_bottom_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_6__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l2_in_0_/S mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l3_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l1_in_1_/X mux_bottom_track_13.mux_l1_in_0_/X
+ mux_bottom_track_13.mux_l2_in_0_/S mux_bottom_track_13.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l1_in_0_ right_bottom_grid_pin_37_ right_top_grid_pin_1_ mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__089__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chanx_right_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_13.mux_l1_in_1_ _045_/HI chanx_left_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _094_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l2_in_1_ _051_/HI chanx_left_in[18] mux_bottom_track_25.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_099_ chanx_left_in[0] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1_ _028_/HI chanx_left_in[15] mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l4_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_11.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_19.mux_l1_in_1_/S mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 mux_right_track_24.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l2_in_3__A0 _029_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__A1 chanx_left_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l2_in_3_ _032_/HI left_bottom_grid_pin_40_ mux_left_track_3.mux_l2_in_0_/S
+ mux_left_track_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.mux_l1_in_0_ bottom_left_grid_pin_44_ chanx_right_in[10] mux_bottom_track_13.mux_l1_in_1_/S
+ mux_bottom_track_13.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l3_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_0_ bottom_left_grid_pin_42_ mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_0_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_13.mux_l1_in_1__S mux_bottom_track_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_098_ _098_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A0 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l4_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_16.mux_l1_in_2__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ chanx_left_in[8] mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_0_/S mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l3_in_1_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 mux_right_track_32.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_5_ chany_bottom_in[17] chany_bottom_in[10] mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_3__A1 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l4_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A0 mux_bottom_track_19.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_38_ left_bottom_grid_pin_36_ mux_left_track_3.mux_l2_in_0_/S
+ mux_left_track_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_21.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_3_ _041_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_3_/S
+ mux_right_track_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_097_ _097_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_32.mux_l1_in_1__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l3_in_1_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ chanx_right_in[19] chanx_right_in[18] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ chany_bottom_in[3] right_bottom_grid_pin_41_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_19.mux_l1_in_1__A1 chanx_left_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[8] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _114_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_5__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l3_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_19.mux_l2_in_0__A1 mux_bottom_track_19.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l2_in_1_ left_bottom_grid_pin_34_ chany_bottom_in[14] mux_left_track_3.mux_l2_in_0_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_3__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A mux_left_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__100__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_5.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 mux_left_track_5.mux_l1_in_5_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_3_/S mux_right_track_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_096_ _096_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_0.mux_l1_in_2_/S mux_right_track_0.mux_l2_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_1__S mux_bottom_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_15.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_24.mux_l1_in_3__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_3_ _037_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l3_in_1__A0 mux_left_track_5.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_40_ right_bottom_grid_pin_39_
+ mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__S mux_bottom_track_19.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__A1 mux_bottom_track_27.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__103__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l4_in_0__A0 mux_left_track_5.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_1_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l1_in_3__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_095_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 mux_left_track_5.mux_l1_in_4_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_3_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_right_track_0.mux_l1_in_2_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l2_in_0__A0 mux_left_track_33.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] chany_bottom_in[15] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_38_ right_bottom_grid_pin_37_
+ mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_1__A1 mux_left_track_5.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_24.mux_l2_in_1_/S
+ mux_right_track_24.mux_l3_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_5.mux_l4_in_0__A1 mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_1__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A0 mux_right_track_0.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_33.mux_l2_in_1_/S ccff_tail
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l2_in_3__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l4_in_0__S mux_left_track_3.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_3_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l2_in_3__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_094_ _094_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l4_in_0__A0 mux_right_track_0.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_1__S mux_left_track_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l2_in_0__A1 mux_left_track_33.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_077_ _077_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_35_
+ mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l2_in_1_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l2_in_2__A1 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_21.mux_l2_in_0__S mux_bottom_track_21.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l1_in_6__A0 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_15.mux_l1_in_0__S mux_bottom_track_15.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l2_in_0_/S mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_1__A1 mux_right_track_0.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l2_in_1_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 mux_bottom_track_1.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l3_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_093_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_0.mux_l4_in_0__A1 mux_right_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l1_in_3_ _054_/HI chanx_left_in[7] mux_bottom_track_5.mux_l1_in_3_/S
+ mux_bottom_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_076_ _076_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ right_bottom_grid_pin_34_
+ mux_right_track_16.mux_l1_in_3_/S mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ right_bottom_grid_pin_34_ right_top_grid_pin_1_ mux_right_track_4.mux_l1_in_2_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _096_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_17.mux_l2_in_1__S mux_left_track_17.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chanx_right_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_3_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_6__A1 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_21.mux_l2_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/S mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_0_/S
+ mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_prog_clk clkbuf_2_0_0_prog_clk/X clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l2_in_1_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_092_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A mux_left_track_3.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_3__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l1_in_2_ chanx_left_in[5] bottom_left_grid_pin_48_ mux_bottom_track_5.mux_l1_in_3_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_075_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__S mux_right_track_4.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l4_in_0__S mux_right_track_2.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l3_in_1__S mux_left_track_5.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A0 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _090_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l3_in_1__S mux_right_track_8.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ _058_/A SC_OUT_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_7.mux_l2_in_1_/S
+ mux_bottom_track_7.mux_l3_in_0_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l1_in_1_/X mux_bottom_track_19.mux_l1_in_0_/X
+ mux_bottom_track_19.mux_l2_in_0_/S mux_bottom_track_19.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l1_in_1_/X mux_bottom_track_21.mux_l1_in_0_/X
+ mux_bottom_track_21.mux_l2_in_0_/S mux_bottom_track_21.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_19.mux_l1_in_1_ _048_/HI chanx_left_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A mux_left_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__S mux_bottom_track_23.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_21.mux_l1_in_1_ _049_/HI chanx_left_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0__S mux_bottom_track_11.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_091_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_32.mux_l3_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A0 mux_bottom_track_11.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A0 bottom_left_grid_pin_48_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_5.mux_l1_in_3_/S mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _074_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_057_ _057_/A SC_OUT_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l2_in_1_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_7.mux_l3_in_0__S mux_bottom_track_7.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A mux_left_track_9.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_3_ _035_/HI left_bottom_grid_pin_41_ mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_3_ _036_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l1_in_0_ bottom_left_grid_pin_47_ chanx_right_in[14] mux_bottom_track_19.mux_l1_in_1_/S
+ mux_bottom_track_19.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_1__A1 chanx_left_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__065__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.mux_l1_in_0_ bottom_left_grid_pin_48_ chanx_right_in[16] mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ _090_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__A1 mux_bottom_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_21.mux_l1_in_0__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _116_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_3_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_073_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_3__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l3_in_0_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__073__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_27.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_056_ SC_IN_BOT SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_7.mux_l1_in_3_/S mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_3__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__068__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l3_in_1__S mux_left_track_1.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A0 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l3_in_1__S mux_right_track_4.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l1_in_3_ _030_/HI left_bottom_grid_pin_38_ mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_37_ left_top_grid_pin_1_ mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l3_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] chany_bottom_in[19] mux_right_track_0.mux_l2_in_0_/S
+ mux_right_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_7.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__081__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _062_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l2_in_0__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__S mux_right_track_32.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A0 mux_bottom_track_15.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l2_in_1_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__084__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_5__A1 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l2_in_0_/S mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_34_ chany_bottom_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ _107_/A chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[9] mux_left_track_9.mux_l2_in_1_/S
+ mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__079__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_1_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__S mux_bottom_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_1__S mux_bottom_track_11.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__S mux_left_track_25.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_15.mux_l1_in_1__A1 chanx_left_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A0 mux_bottom_track_7.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[5] right_bottom_grid_pin_41_ mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A0 mux_bottom_track_23.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__087__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0__A1 mux_bottom_track_15.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A0 mux_bottom_track_7.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_19.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_3_ _039_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chanx_right_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_13.mux_l2_in_0_/S
+ mux_bottom_track_15.mux_l1_in_1_/S mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_106_ _106_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_1_ chany_bottom_in[10] chany_bottom_in[3] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A0 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[2] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_1_/S mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__095__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_2__A1 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_0_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_1__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l3_in_1__S mux_right_track_0.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_3.mux_l2_in_2__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A0 mux_left_track_1.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_1__A1 mux_bottom_track_7.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.mux_l2_in_0__A1 mux_bottom_track_23.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_0.mux_l1_in_2_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l4_in_0__A0 mux_left_track_1.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_070_ _070_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_7.mux_l3_in_0__A1 mux_bottom_track_7.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_3__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] chany_bottom_in[14] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__098__A _098_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A0 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_13.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_105_ _105_/A chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chanx_right_in[17] chanx_right_in[8] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l2_in_2__A1 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A mux_left_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l4_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _098_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_3_ _043_/HI chanx_left_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_1__A1 mux_left_track_1.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_35_ right_top_grid_pin_1_ mux_right_track_0.mux_l1_in_2_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_1_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_1.mux_l4_in_0__A1 mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A0 bottom_left_grid_pin_43_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_1_ chany_bottom_in[7] chany_bottom_in[0] mux_right_track_24.mux_l1_in_3_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_3__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l1_in_0__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l4_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ chanx_right_in[11] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_41_ left_bottom_grid_pin_40_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_2_ chanx_left_in[1] bottom_left_grid_pin_48_ mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 mux_left_track_5.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l2_in_2__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l1_in_1_/X mux_bottom_track_15.mux_l1_in_0_/X
+ mux_bottom_track_15.mux_l2_in_0_/S mux_bottom_track_15.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_27.mux_l1_in_0__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_23.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_3__A0 _032_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_39_ right_bottom_grid_pin_35_
+ mux_right_track_24.mux_l1_in_3_/S mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_16.mux_l1_in_3__A1 chanx_left_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_15.mux_l1_in_1_ _046_/HI chanx_left_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l3_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_4_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_103_ chanx_right_in[7] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_5_ left_bottom_grid_pin_39_ left_bottom_grid_pin_38_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_5.mux_l1_in_4_/S mux_left_track_5.mux_l2_in_1_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_21.mux_l1_in_0__S mux_bottom_track_21.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l1_in_1__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_6__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_1.mux_l1_in_0_/S mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_8.mux_l3_in_1_/S mux_right_track_8.mux_l4_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__101__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_3__A1 chanx_left_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l2_in_3__A1 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_3_ _034_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_1_/S
+ mux_left_track_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_7.mux_l1_in_2__S mux_bottom_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_15.mux_l1_in_0_ bottom_left_grid_pin_45_ chanx_right_in[12] mux_bottom_track_15.mux_l1_in_1_/S
+ mux_bottom_track_15.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_2.mux_l1_in_0_/S mux_right_track_2.mux_l2_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_bottom_track_27.mux_l2_in_0_ _052_/HI mux_bottom_track_27.mux_l1_in_0_/X mux_bottom_track_27.mux_l2_in_0_/S
+ mux_bottom_track_27.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0__S mux_bottom_track_13.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _118_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_102_ chanx_right_in[3] chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_5.mux_l1_in_4_ left_bottom_grid_pin_37_ left_bottom_grid_pin_36_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_16.mux_l2_in_1__S mux_right_track_16.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_19.mux_l1_in_1__S mux_bottom_track_19.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_4_/S
+ mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__104__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_0_ bottom_left_grid_pin_42_ chanx_right_in[2] mux_bottom_track_1.mux_l1_in_0_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_1_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_7.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_3__A0 _030_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_2_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ chanx_right_in[1] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_032_ _032_/HI _032_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_2_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_35_ left_bottom_grid_pin_34_ mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_46_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l1_in_5__A0 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_27.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[15] mux_bottom_track_27.mux_l1_in_0_/S
+ mux_bottom_track_27.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _070_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_3__A0 _031_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_6__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_25.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_3__A1 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_100_ chanx_right_in[0] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_031_ _031_/HI _031_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_2__S mux_bottom_track_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_left_grid_pin_44_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__118__A _118_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_15.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_1_ chany_bottom_in[15] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_3_ _031_/HI left_bottom_grid_pin_39_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_5__A1 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__S mux_bottom_track_7.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_2__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_1__S mux_bottom_track_15.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_25.mux_l1_in_3__A1 left_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l3_in_1__A0 mux_right_track_2.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l3_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_030_ _030_/HI _030_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_1_ chany_bottom_in[8] chany_bottom_in[1] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_35_ chany_bottom_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A0 mux_right_track_2.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_3_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A0 chanx_left_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_23.mux_l2_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A1 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__S mux_left_track_33.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_1_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_9.mux_l2_in_3__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l3_in_1__A1 mux_right_track_2.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_3.mux_l1_in_2_/S
+ mux_bottom_track_3.mux_l2_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 mux_bottom_track_3.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_11.mux_l3_in_0_ mux_bottom_track_11.mux_l2_in_1_/X mux_bottom_track_11.mux_l2_in_0_/X
+ mux_bottom_track_11.mux_l3_in_0_/S mux_bottom_track_11.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A mux_left_track_5.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_0_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l1_in_4_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_9.mux_l4_in_0__S mux_left_track_9.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_089_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__060__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l4_in_0__A1 mux_right_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_11.mux_l2_in_0__A1 mux_bottom_track_11.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.mux_l2_in_1_ _044_/HI chanx_left_in[19] mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_9.mux_l2_in_0_/S
+ mux_bottom_track_9.mux_l3_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chanx_right_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_1_ _040_/HI chanx_left_in[10] mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_25.mux_l2_in_0__S mux_left_track_25.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_27.mux_l2_in_0__S mux_bottom_track_27.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_2_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__063__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_3__A1 left_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_2_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 mux_bottom_track_3.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_11.mux_l2_in_0_/S
+ mux_bottom_track_11.mux_l3_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_0_ chanx_right_in[18] chanx_right_in[9] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_088_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l1_in_3_ _055_/HI chanx_left_in[11] mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_11.mux_l2_in_0_ chanx_left_in[9] mux_bottom_track_11.mux_l1_in_0_/X
+ mux_bottom_track_11.mux_l2_in_0_/S mux_bottom_track_11.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__071__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l2_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l3_in_0__S mux_left_track_17.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A0 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__066__A _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 right_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ mux_bottom_track_7.mux_l3_in_0_/S mux_bottom_track_7.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l1_in_3_/X mux_bottom_track_7.mux_l1_in_2_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_4__A1 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l2_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__069__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A0 bottom_left_grid_pin_47_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A0 bottom_left_grid_pin_49_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _086_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_11.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_2_ chanx_left_in[6] bottom_left_grid_pin_49_ mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l4_in_0__S mux_left_track_5.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_3__A1 mux_right_track_4.mux_l1_in_6_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_7.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l4_in_0__S mux_right_track_8.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0__A1 chanx_right_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A0 mux_bottom_track_7.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_3_ _029_/HI left_bottom_grid_pin_41_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_11.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[9] mux_bottom_track_11.mux_l1_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l1_in_1_/X mux_bottom_track_23.mux_l1_in_0_/X
+ mux_bottom_track_23.mux_l2_in_0_/S mux_bottom_track_23.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_9.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l2_in_1__S mux_left_track_33.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_0_ right_bottom_grid_pin_40_ right_bottom_grid_pin_36_
+ mux_right_track_32.mux_l1_in_0_/S mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_23.mux_l2_in_0__S mux_bottom_track_23.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_23.mux_l1_in_1_ _050_/HI chanx_left_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S mux_bottom_track_7.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_086_ _086_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_11.mux_l1_in_0_/S mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__085__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_7.mux_l1_in_1__A1 bottom_left_grid_pin_45_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_23.mux_l1_in_0__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_7.mux_l1_in_1_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_7.mux_l1_in_3_/S mux_bottom_track_7.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l2_in_0_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0__A1 mux_bottom_track_7.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_39_ left_bottom_grid_pin_37_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_3_ _038_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__088__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.mux_l1_in_0_ bottom_left_grid_pin_49_ chanx_right_in[17] mux_bottom_track_23.mux_l1_in_0_/S
+ mux_bottom_track_23.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A0 mux_right_track_8.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 left_top_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l4_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_7.mux_l1_in_0_ bottom_left_grid_pin_43_ chanx_right_in[6] mux_bottom_track_7.mux_l1_in_3_/S
+ mux_bottom_track_7.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X _115_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l4_in_0__A0 mux_right_track_8.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_15.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l1_in_0_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_left_track_1.mux_l2_in_1_ left_bottom_grid_pin_35_ left_top_grid_pin_1_ mux_left_track_1.mux_l2_in_0_/S
+ mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l2_in_3__S mux_left_track_3.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l4_in_0__S mux_left_track_1.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_4.mux_l4_in_0__S mux_right_track_4.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] chany_bottom_in[18] mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l3_in_1__A1 mux_right_track_8.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_084_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_left_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 _028_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 mux_right_track_16.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0__S mux_bottom_track_13.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_067_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l4_in_0__A1 mux_right_track_8.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A0 mux_right_track_16.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_1_ chany_bottom_in[13] chany_bottom_in[6] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l2_in_2__A0 left_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l2_in_1_ chany_bottom_in[11] chany_bottom_in[4] mux_right_track_2.mux_l2_in_0_/S
+ mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_11.mux_l3_in_0__S mux_bottom_track_11.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2__A1 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 mux_right_track_24.mux_l1_in_3_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_3.mux_l3_in_1__A0 mux_left_track_3.mux_l2_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_083_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 chanx_left_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_1__A1 mux_right_track_16.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_066_ _066_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A0 mux_left_track_3.mux_l3_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l3_in_0__A1 mux_right_track_16.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_ mux_right_track_4.mux_l3_in_1_/S mux_right_track_4.mux_l4_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_118_ _118_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l1_in_2__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l2_in_1__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[2] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l2_in_2__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_3__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__S mux_left_track_5.mux_l1_in_4_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l4_in_0__S mux_right_track_0.mux_l4_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l3_in_1__S mux_left_track_3.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l2_in_1_ _033_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_1_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 mux_right_track_24.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l2_in_2__S mux_left_track_9.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l3_in_0__A0 mux_right_track_32.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l3_in_1__A1 mux_left_track_3.mux_l2_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _082_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_2.mux_l1_in_0_/S mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_40_ left_bottom_grid_pin_36_
+ mux_left_track_33.mux_l1_in_0_/S mux_left_track_33.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_left_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_27.mux_l2_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_3.mux_l4_in_0__A1 mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_left_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_21.mux_l1_in_1__S mux_bottom_track_21.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0__S mux_bottom_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_13.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_117_ _117_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_4.mux_l2_in_3_/S mux_right_track_4.mux_l3_in_1_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l1_in_2__S mux_right_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2__A0 left_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_32.mux_l2_in_1__A1 chanx_left_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D mux_left_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 mux_left_track_17.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_3_ _053_/HI chanx_left_in[4] mux_bottom_track_3.mux_l1_in_2_/S
+ mux_bottom_track_3.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l3_in_0__A1 mux_right_track_32.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _097_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D mux_right_track_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_7.mux_l1_in_3__S mux_bottom_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_081_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_0_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_2.mux_l1_in_0_/S mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 bottom_left_grid_pin_42_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_1_ chany_bottom_in[19] chany_bottom_in[12] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_4__A0 left_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_left_track_17.mux_l1_in_2__S mux_left_track_17.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A0 mux_left_track_17.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_064_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_4.mux_l1_in_2_/S mux_right_track_4.mux_l2_in_3_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_left_track_5.mux_l2_in_3__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_116_ _116_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 left_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l2_in_1__A0 mux_left_track_25.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l2_in_1__A1 mux_left_track_17.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_2_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_3.mux_l1_in_2_/S
+ mux_bottom_track_3.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l3_in_0__A0 mux_left_track_25.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_4.mux_l1_in_4__S mux_right_track_4.mux_l1_in_2_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_0_ chany_bottom_in[5] chanx_right_in[10] mux_left_track_33.mux_l1_in_0_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l3_in_1__S mux_right_track_2.mux_l3_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__108__A _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_23.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_4__A1 left_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_2__S mux_left_track_5.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_17.mux_l3_in_0__A1 mux_left_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_2__S mux_right_track_8.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_2__A0 left_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_2_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 mux_left_track_5.mux_l1_in_6_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_115_ _115_/A chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l2_in_1__A0 _033_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l1_in_1_ _047_/HI chanx_left_in[13] mux_bottom_track_17.mux_l1_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_029_ _029_/HI _029_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_21.mux_l1_in_1_/S
+ mux_bottom_track_21.mux_l2_in_0_/S mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_left_track_25.mux_l2_in_1__A1 mux_left_track_25.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l3_in_0__A0 mux_left_track_33.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_27.mux_l1_in_0__S mux_bottom_track_27.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

