magic
tech sky130A
magscale 1 2
timestamp 1606236195
<< locali >>
rect 9229 5151 9263 5253
rect 9321 5083 9355 5253
rect 7389 4471 7423 4641
<< viali >>
rect 1593 6409 1627 6443
rect 11713 6409 11747 6443
rect 2881 6273 2915 6307
rect 4169 6273 4203 6307
rect 7021 6273 7055 6307
rect 7389 6273 7423 6307
rect 8401 6273 8435 6307
rect 9045 6273 9079 6307
rect 10517 6273 10551 6307
rect 12725 6273 12759 6307
rect 14105 6273 14139 6307
rect 1409 6205 1443 6239
rect 1961 6205 1995 6239
rect 5457 6205 5491 6239
rect 5825 6205 5859 6239
rect 11529 6205 11563 6239
rect 2605 6137 2639 6171
rect 2697 6137 2731 6171
rect 4261 6137 4295 6171
rect 5181 6137 5215 6171
rect 6193 6137 6227 6171
rect 7113 6137 7147 6171
rect 8493 6137 8527 6171
rect 10241 6137 10275 6171
rect 10333 6137 10367 6171
rect 12817 6137 12851 6171
rect 13737 6137 13771 6171
rect 14197 6137 14231 6171
rect 15117 6137 15151 6171
rect 2145 6069 2179 6103
rect 9229 5865 9263 5899
rect 9873 5865 9907 5899
rect 10425 5865 10459 5899
rect 12403 5865 12437 5899
rect 14289 5865 14323 5899
rect 14841 5865 14875 5899
rect 1869 5797 1903 5831
rect 1961 5797 1995 5831
rect 4215 5797 4249 5831
rect 4629 5797 4663 5831
rect 4721 5797 4755 5831
rect 6377 5797 6411 5831
rect 6469 5797 6503 5831
rect 7757 5797 7791 5831
rect 7849 5797 7883 5831
rect 10885 5797 10919 5831
rect 10977 5797 11011 5831
rect 12909 5797 12943 5831
rect 3157 5729 3191 5763
rect 4123 5729 4157 5763
rect 9045 5729 9079 5763
rect 9689 5729 9723 5763
rect 10241 5729 10275 5763
rect 12332 5729 12366 5763
rect 14105 5729 14139 5763
rect 14657 5729 14691 5763
rect 2145 5661 2179 5695
rect 5457 5661 5491 5695
rect 7389 5661 7423 5695
rect 8769 5661 8803 5695
rect 11897 5661 11931 5695
rect 12817 5661 12851 5695
rect 13829 5661 13863 5695
rect 3341 5525 3375 5559
rect 1961 5321 1995 5355
rect 10379 5321 10413 5355
rect 13185 5321 13219 5355
rect 14105 5321 14139 5355
rect 2329 5253 2363 5287
rect 3709 5253 3743 5287
rect 9229 5253 9263 5287
rect 7849 5185 7883 5219
rect 8585 5185 8619 5219
rect 1777 5117 1811 5151
rect 2697 5117 2731 5151
rect 4077 5117 4111 5151
rect 5089 5117 5123 5151
rect 5356 5117 5390 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 7573 5117 7607 5151
rect 8217 5117 8251 5151
rect 8861 5117 8895 5151
rect 9229 5117 9263 5151
rect 9321 5253 9355 5287
rect 9597 5253 9631 5287
rect 14657 5253 14691 5287
rect 9413 5117 9447 5151
rect 10308 5117 10342 5151
rect 13001 5117 13035 5151
rect 13921 5117 13955 5151
rect 14473 5117 14507 5151
rect 3065 5049 3099 5083
rect 4445 5049 4479 5083
rect 9321 5049 9355 5083
rect 6469 4981 6503 5015
rect 9045 4981 9079 5015
rect 5457 4777 5491 4811
rect 9275 4777 9309 4811
rect 4322 4709 4356 4743
rect 6092 4709 6126 4743
rect 7726 4709 7760 4743
rect 1593 4641 1627 4675
rect 2412 4641 2446 4675
rect 7389 4641 7423 4675
rect 9172 4641 9206 4675
rect 10828 4641 10862 4675
rect 14013 4641 14047 4675
rect 2145 4573 2179 4607
rect 4077 4573 4111 4607
rect 5825 4573 5859 4607
rect 1777 4505 1811 4539
rect 7481 4573 7515 4607
rect 3525 4437 3559 4471
rect 7205 4437 7239 4471
rect 7389 4437 7423 4471
rect 8861 4437 8895 4471
rect 10931 4437 10965 4471
rect 14197 4437 14231 4471
rect 4261 4233 4295 4267
rect 2881 4097 2915 4131
rect 4629 4097 4663 4131
rect 6929 4097 6963 4131
rect 7941 4097 7975 4131
rect 10977 4097 11011 4131
rect 1869 4029 1903 4063
rect 2237 4029 2271 4063
rect 2605 4029 2639 4063
rect 3148 4029 3182 4063
rect 5917 4029 5951 4063
rect 8217 4029 8251 4063
rect 4721 3961 4755 3995
rect 5641 3961 5675 3995
rect 7021 3961 7055 3995
rect 11069 3961 11103 3995
rect 11989 3961 12023 3995
rect 6101 3893 6135 3927
rect 8401 3893 8435 3927
rect 3249 3689 3283 3723
rect 7573 3689 7607 3723
rect 8079 3689 8113 3723
rect 2136 3621 2170 3655
rect 3663 3621 3697 3655
rect 4261 3621 4295 3655
rect 3560 3553 3594 3587
rect 5733 3553 5767 3587
rect 6000 3553 6034 3587
rect 7389 3553 7423 3587
rect 7976 3553 8010 3587
rect 1869 3485 1903 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 7113 3349 7147 3383
rect 3249 3145 3283 3179
rect 7389 3077 7423 3111
rect 4859 3009 4893 3043
rect 5273 3009 5307 3043
rect 2513 2941 2547 2975
rect 3065 2941 3099 2975
rect 3709 2941 3743 2975
rect 4077 2941 4111 2975
rect 4756 2941 4790 2975
rect 6837 2941 6871 2975
rect 7205 2941 7239 2975
rect 9781 2941 9815 2975
rect 4445 2873 4479 2907
rect 5365 2873 5399 2907
rect 6285 2873 6319 2907
rect 2697 2805 2731 2839
rect 9965 2805 9999 2839
rect 3065 2601 3099 2635
rect 3617 2601 3651 2635
rect 4261 2601 4295 2635
rect 5411 2601 5445 2635
rect 1941 2465 1975 2499
rect 3433 2465 3467 2499
rect 4077 2465 4111 2499
rect 5308 2465 5342 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 7297 2465 7331 2499
rect 7941 2465 7975 2499
rect 1685 2397 1719 2431
rect 7665 2397 7699 2431
rect 6469 2261 6503 2295
rect 8125 2261 8159 2295
<< metal1 >>
rect 3418 7080 3424 7132
rect 3476 7120 3482 7132
rect 8938 7120 8944 7132
rect 3476 7092 8944 7120
rect 3476 7080 3482 7092
rect 8938 7080 8944 7092
rect 8996 7080 9002 7132
rect 3050 6876 3056 6928
rect 3108 6916 3114 6928
rect 7742 6916 7748 6928
rect 3108 6888 7748 6916
rect 3108 6876 3114 6888
rect 7742 6876 7748 6888
rect 7800 6876 7806 6928
rect 13078 6672 13084 6724
rect 13136 6712 13142 6724
rect 13538 6712 13544 6724
rect 13136 6684 13544 6712
rect 13136 6672 13142 6684
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 198 6400 204 6452
rect 256 6440 262 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 256 6412 1593 6440
rect 256 6400 262 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 11698 6440 11704 6452
rect 1581 6403 1639 6409
rect 7024 6412 11560 6440
rect 11659 6412 11704 6440
rect 1118 6332 1124 6384
rect 1176 6372 1182 6384
rect 2590 6372 2596 6384
rect 1176 6344 2596 6372
rect 1176 6332 1182 6344
rect 1412 6245 1440 6344
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 1964 6276 2881 6304
rect 1964 6245 1992 6276
rect 2869 6273 2881 6276
rect 2915 6273 2927 6307
rect 4154 6304 4160 6316
rect 4115 6276 4160 6304
rect 2869 6267 2927 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 7024 6313 7052 6412
rect 9122 6372 9128 6384
rect 8404 6344 9128 6372
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7374 6304 7380 6316
rect 7335 6276 7380 6304
rect 7009 6267 7067 6273
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 8404 6313 8432 6344
rect 9122 6332 9128 6344
rect 9180 6332 9186 6384
rect 11532 6372 11560 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 15194 6372 15200 6384
rect 11532 6344 15200 6372
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 8389 6267 8447 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10226 6304 10232 6316
rect 9732 6276 10232 6304
rect 9732 6264 9738 6276
rect 10226 6264 10232 6276
rect 10284 6304 10290 6316
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10284 6276 10517 6304
rect 10284 6264 10290 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12216 6276 12725 6304
rect 12216 6264 12222 6276
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6304 14151 6307
rect 16206 6304 16212 6316
rect 14139 6276 16212 6304
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1949 6239 2007 6245
rect 1949 6205 1961 6239
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5132 6208 5457 6236
rect 5132 6196 5138 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5810 6236 5816 6248
rect 5771 6208 5816 6236
rect 5445 6199 5503 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 11204 6208 11529 6236
rect 11204 6196 11210 6208
rect 11517 6205 11529 6208
rect 11563 6236 11575 6239
rect 11974 6236 11980 6248
rect 11563 6208 11980 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 2593 6171 2651 6177
rect 2593 6168 2605 6171
rect 1728 6140 2605 6168
rect 1728 6128 1734 6140
rect 2593 6137 2605 6140
rect 2639 6137 2651 6171
rect 2593 6131 2651 6137
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6137 2743 6171
rect 2685 6131 2743 6137
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 4522 6168 4528 6180
rect 4295 6140 4528 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 2498 6100 2504 6112
rect 2179 6072 2504 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 2700 6100 2728 6131
rect 4522 6128 4528 6140
rect 4580 6128 4586 6180
rect 5166 6168 5172 6180
rect 5079 6140 5172 6168
rect 5166 6128 5172 6140
rect 5224 6168 5230 6180
rect 5350 6168 5356 6180
rect 5224 6140 5356 6168
rect 5224 6128 5230 6140
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 6181 6171 6239 6177
rect 6181 6137 6193 6171
rect 6227 6137 6239 6171
rect 6181 6131 6239 6137
rect 7101 6171 7159 6177
rect 7101 6137 7113 6171
rect 7147 6168 7159 6171
rect 8481 6171 8539 6177
rect 7147 6140 8248 6168
rect 7147 6137 7159 6140
rect 7101 6131 7159 6137
rect 3326 6100 3332 6112
rect 2700 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 6196 6100 6224 6131
rect 6914 6100 6920 6112
rect 6196 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 7374 6100 7380 6112
rect 7064 6072 7380 6100
rect 7064 6060 7070 6072
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8220 6100 8248 6140
rect 8481 6137 8493 6171
rect 8527 6168 8539 6171
rect 8754 6168 8760 6180
rect 8527 6140 8760 6168
rect 8527 6137 8539 6140
rect 8481 6131 8539 6137
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 9214 6100 9220 6112
rect 8220 6072 9220 6100
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 10244 6100 10272 6131
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 10376 6140 10421 6168
rect 10376 6128 10382 6140
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 12342 6168 12348 6180
rect 10560 6140 12348 6168
rect 10560 6128 10566 6140
rect 12342 6128 12348 6140
rect 12400 6168 12406 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12400 6140 12817 6168
rect 12400 6128 12406 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 13725 6171 13783 6177
rect 13725 6137 13737 6171
rect 13771 6168 13783 6171
rect 13906 6168 13912 6180
rect 13771 6140 13912 6168
rect 13771 6137 13783 6140
rect 13725 6131 13783 6137
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 14090 6128 14096 6180
rect 14148 6168 14154 6180
rect 14185 6171 14243 6177
rect 14185 6168 14197 6171
rect 14148 6140 14197 6168
rect 14148 6128 14154 6140
rect 14185 6137 14197 6140
rect 14231 6137 14243 6171
rect 15102 6168 15108 6180
rect 15063 6140 15108 6168
rect 14185 6131 14243 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 15654 6100 15660 6112
rect 10244 6072 15660 6100
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6328 5868 6408 5896
rect 6328 5856 6334 5868
rect 1854 5828 1860 5840
rect 1815 5800 1860 5828
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 1949 5831 2007 5837
rect 1949 5797 1961 5831
rect 1995 5828 2007 5831
rect 4203 5831 4261 5837
rect 4203 5828 4215 5831
rect 1995 5800 4215 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 4203 5797 4215 5800
rect 4249 5797 4261 5831
rect 4614 5828 4620 5840
rect 4575 5800 4620 5828
rect 4203 5791 4261 5797
rect 4614 5788 4620 5800
rect 4672 5788 4678 5840
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 6380 5837 6408 5868
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 8996 5868 9229 5896
rect 8996 5856 9002 5868
rect 9217 5865 9229 5868
rect 9263 5865 9275 5899
rect 9217 5859 9275 5865
rect 9861 5899 9919 5905
rect 9861 5865 9873 5899
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 6365 5831 6423 5837
rect 4764 5800 4809 5828
rect 4764 5788 4770 5800
rect 6365 5797 6377 5831
rect 6411 5797 6423 5831
rect 6365 5791 6423 5797
rect 6457 5831 6515 5837
rect 6457 5797 6469 5831
rect 6503 5828 6515 5831
rect 6914 5828 6920 5840
rect 6503 5800 6920 5828
rect 6503 5797 6515 5800
rect 6457 5791 6515 5797
rect 6914 5788 6920 5800
rect 6972 5828 6978 5840
rect 7742 5828 7748 5840
rect 6972 5800 7236 5828
rect 7703 5800 7748 5828
rect 6972 5788 6978 5800
rect 3145 5763 3203 5769
rect 3145 5729 3157 5763
rect 3191 5729 3203 5763
rect 3145 5723 3203 5729
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 3160 5624 3188 5723
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 4111 5763 4169 5769
rect 4111 5760 4123 5763
rect 3384 5732 4123 5760
rect 3384 5720 3390 5732
rect 4111 5729 4123 5732
rect 4157 5729 4169 5763
rect 4111 5723 4169 5729
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 7208 5624 7236 5800
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 7892 5800 7937 5828
rect 7892 5788 7898 5800
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 9876 5828 9904 5859
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10413 5899 10471 5905
rect 10413 5896 10425 5899
rect 10192 5868 10425 5896
rect 10192 5856 10198 5868
rect 10413 5865 10425 5868
rect 10459 5865 10471 5899
rect 10413 5859 10471 5865
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 12391 5899 12449 5905
rect 10652 5868 11008 5896
rect 10652 5856 10658 5868
rect 8720 5800 9904 5828
rect 8720 5788 8726 5800
rect 10686 5788 10692 5840
rect 10744 5828 10750 5840
rect 10980 5837 11008 5868
rect 12391 5865 12403 5899
rect 12437 5896 12449 5899
rect 14090 5896 14096 5908
rect 12437 5868 14096 5896
rect 12437 5865 12449 5868
rect 12391 5859 12449 5865
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 14240 5868 14289 5896
rect 14240 5856 14246 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14700 5868 14841 5896
rect 14700 5856 14706 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 10873 5831 10931 5837
rect 10873 5828 10885 5831
rect 10744 5800 10885 5828
rect 10744 5788 10750 5800
rect 10873 5797 10885 5800
rect 10919 5797 10931 5831
rect 10873 5791 10931 5797
rect 10965 5831 11023 5837
rect 10965 5797 10977 5831
rect 11011 5797 11023 5831
rect 12897 5831 12955 5837
rect 12897 5828 12909 5831
rect 10965 5791 11023 5797
rect 11716 5800 12909 5828
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 10226 5760 10232 5772
rect 10187 5732 10232 5760
rect 9677 5723 9735 5729
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 8662 5692 8668 5704
rect 7423 5664 8668 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 9692 5692 9720 5723
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 8803 5664 9720 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 7558 5624 7564 5636
rect 3160 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 8772 5624 8800 5655
rect 11716 5624 11744 5800
rect 12897 5797 12909 5800
rect 12943 5828 12955 5831
rect 12943 5800 14136 5828
rect 12943 5797 12955 5800
rect 12897 5791 12955 5797
rect 12342 5769 12348 5772
rect 12320 5763 12348 5769
rect 12320 5729 12332 5763
rect 12320 5723 12348 5729
rect 12342 5720 12348 5723
rect 12400 5720 12406 5772
rect 14108 5769 14136 5800
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5661 11943 5695
rect 12802 5692 12808 5704
rect 12763 5664 12808 5692
rect 11885 5655 11943 5661
rect 8352 5596 8800 5624
rect 8864 5596 11744 5624
rect 11900 5624 11928 5655
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13817 5695 13875 5701
rect 13817 5661 13829 5695
rect 13863 5692 13875 5695
rect 13998 5692 14004 5704
rect 13863 5664 14004 5692
rect 13863 5661 13875 5664
rect 13817 5655 13875 5661
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14458 5624 14464 5636
rect 11900 5596 14464 5624
rect 8352 5584 8358 5596
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3329 5559 3387 5565
rect 3329 5556 3341 5559
rect 2832 5528 3341 5556
rect 2832 5516 2838 5528
rect 3329 5525 3341 5528
rect 3375 5525 3387 5559
rect 3329 5519 3387 5525
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 8864 5556 8892 5596
rect 14458 5584 14464 5596
rect 14516 5584 14522 5636
rect 7800 5528 8892 5556
rect 7800 5516 7806 5528
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 14660 5556 14688 5723
rect 10468 5528 14688 5556
rect 10468 5516 10474 5528
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 2682 5352 2688 5364
rect 1995 5324 2688 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5408 5324 6040 5352
rect 5408 5312 5414 5324
rect 1854 5244 1860 5296
rect 1912 5284 1918 5296
rect 2317 5287 2375 5293
rect 2317 5284 2329 5287
rect 1912 5256 2329 5284
rect 1912 5244 1918 5256
rect 2317 5253 2329 5256
rect 2363 5284 2375 5287
rect 3697 5287 3755 5293
rect 3697 5284 3709 5287
rect 2363 5256 3709 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 3697 5253 3709 5256
rect 3743 5284 3755 5287
rect 5074 5284 5080 5296
rect 3743 5256 5080 5284
rect 3743 5253 3755 5256
rect 3697 5247 3755 5253
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 6012 5284 6040 5324
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 7708 5324 10272 5352
rect 7708 5312 7714 5324
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 6012 5256 9229 5284
rect 9217 5253 9229 5256
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 9309 5287 9367 5293
rect 9309 5253 9321 5287
rect 9355 5284 9367 5287
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 9355 5256 9597 5284
rect 9355 5253 9367 5256
rect 9309 5247 9367 5253
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 10244 5284 10272 5324
rect 10318 5312 10324 5364
rect 10376 5361 10382 5364
rect 10376 5355 10425 5361
rect 10376 5321 10379 5355
rect 10413 5321 10425 5355
rect 13170 5352 13176 5364
rect 13131 5324 13176 5352
rect 10376 5315 10425 5321
rect 10376 5312 10382 5315
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 13688 5324 14105 5352
rect 13688 5312 13694 5324
rect 14093 5321 14105 5324
rect 14139 5321 14151 5355
rect 14093 5315 14151 5321
rect 12802 5284 12808 5296
rect 10244 5256 12808 5284
rect 9585 5247 9643 5253
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 14645 5287 14703 5293
rect 14645 5284 14657 5287
rect 13780 5256 14657 5284
rect 13780 5244 13786 5256
rect 14645 5253 14657 5256
rect 14691 5253 14703 5287
rect 14645 5247 14703 5253
rect 658 5176 664 5228
rect 716 5216 722 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 716 5188 4752 5216
rect 716 5176 722 5188
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5148 1823 5151
rect 2130 5148 2136 5160
rect 1811 5120 2136 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 2774 5148 2780 5160
rect 2731 5120 2780 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4246 5148 4252 5160
rect 4111 5120 4252 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4246 5108 4252 5120
rect 4304 5108 4310 5160
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3326 5080 3332 5092
rect 3099 5052 3332 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 4433 5083 4491 5089
rect 4433 5049 4445 5083
rect 4479 5080 4491 5083
rect 4614 5080 4620 5092
rect 4479 5052 4620 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 4724 5080 4752 5188
rect 6840 5188 7849 5216
rect 6840 5160 6868 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 8754 5216 8760 5228
rect 8619 5188 8760 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8754 5176 8760 5188
rect 8812 5216 8818 5228
rect 15102 5216 15108 5228
rect 8812 5188 9536 5216
rect 8812 5176 8818 5188
rect 5074 5148 5080 5160
rect 5035 5120 5080 5148
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5344 5151 5402 5157
rect 5344 5117 5356 5151
rect 5390 5148 5402 5151
rect 5810 5148 5816 5160
rect 5390 5120 5816 5148
rect 5390 5117 5402 5120
rect 5344 5111 5402 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7190 5148 7196 5160
rect 7151 5120 7196 5148
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 7742 5148 7748 5160
rect 7607 5120 7748 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 8202 5148 8208 5160
rect 8163 5120 8208 5148
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8720 5120 8861 5148
rect 8720 5108 8726 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 9263 5120 9413 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9508 5148 9536 5188
rect 13004 5188 15108 5216
rect 10296 5151 10354 5157
rect 10296 5148 10308 5151
rect 9508 5120 10308 5148
rect 9401 5111 9459 5117
rect 10296 5117 10308 5120
rect 10342 5148 10354 5151
rect 10410 5148 10416 5160
rect 10342 5120 10416 5148
rect 10342 5117 10354 5120
rect 10296 5111 10354 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13004 5157 13032 5188
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12768 5120 13001 5148
rect 12768 5108 12774 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 13906 5148 13912 5160
rect 13867 5120 13912 5148
rect 12989 5111 13047 5117
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 14458 5148 14464 5160
rect 14419 5120 14464 5148
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 6914 5080 6920 5092
rect 4724 5052 6920 5080
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 7064 5052 9321 5080
rect 7064 5040 7070 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9309 5043 9367 5049
rect 6457 5015 6515 5021
rect 6457 4981 6469 5015
rect 6503 5012 6515 5015
rect 7190 5012 7196 5024
rect 6503 4984 7196 5012
rect 6503 4981 6515 4984
rect 6457 4975 6515 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 5012 9091 5015
rect 12434 5012 12440 5024
rect 9079 4984 12440 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 4706 4808 4712 4820
rect 2556 4780 4712 4808
rect 2556 4768 2562 4780
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5810 4808 5816 4820
rect 5491 4780 5816 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 9214 4768 9220 4820
rect 9272 4817 9278 4820
rect 9272 4811 9321 4817
rect 9272 4777 9275 4811
rect 9309 4777 9321 4811
rect 9272 4771 9321 4777
rect 9272 4768 9278 4771
rect 1596 4712 3372 4740
rect 1596 4681 1624 4712
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 2400 4675 2458 4681
rect 2400 4641 2412 4675
rect 2446 4672 2458 4675
rect 2774 4672 2780 4684
rect 2446 4644 2780 4672
rect 2446 4641 2458 4644
rect 2400 4635 2458 4641
rect 2774 4632 2780 4644
rect 2832 4672 2838 4684
rect 3234 4672 3240 4684
rect 2832 4644 3240 4672
rect 2832 4632 2838 4644
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3344 4672 3372 4712
rect 4246 4700 4252 4752
rect 4304 4749 4310 4752
rect 4304 4743 4368 4749
rect 4304 4709 4322 4743
rect 4356 4709 4368 4743
rect 4304 4703 4368 4709
rect 6080 4743 6138 4749
rect 6080 4709 6092 4743
rect 6126 4740 6138 4743
rect 6126 4712 7144 4740
rect 6126 4709 6138 4712
rect 6080 4703 6138 4709
rect 4304 4700 4310 4703
rect 4614 4672 4620 4684
rect 3344 4644 4620 4672
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 7116 4672 7144 4712
rect 7190 4700 7196 4752
rect 7248 4740 7254 4752
rect 7714 4743 7772 4749
rect 7714 4740 7726 4743
rect 7248 4712 7726 4740
rect 7248 4700 7254 4712
rect 7714 4709 7726 4712
rect 7760 4709 7772 4743
rect 7714 4703 7772 4709
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 5828 4644 6868 4672
rect 7116 4644 7389 4672
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 5828 4613 5856 4644
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1728 4576 2145 4604
rect 1728 4564 1734 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 6840 4604 6868 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 9160 4675 9218 4681
rect 9160 4672 9172 4675
rect 7616 4644 9172 4672
rect 7616 4632 7622 4644
rect 9160 4641 9172 4644
rect 9206 4641 9218 4675
rect 9160 4635 9218 4641
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 10816 4675 10874 4681
rect 10816 4672 10828 4675
rect 10652 4644 10828 4672
rect 10652 4632 10658 4644
rect 10816 4641 10828 4644
rect 10862 4641 10874 4675
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 10816 4635 10874 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 6840 4576 7481 4604
rect 5813 4567 5871 4573
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 1762 4536 1768 4548
rect 1723 4508 1768 4536
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 2148 4468 2176 4567
rect 4080 4536 4108 4567
rect 5718 4536 5724 4548
rect 3068 4508 4108 4536
rect 3068 4468 3096 4508
rect 2148 4440 3096 4468
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3513 4471 3571 4477
rect 3513 4468 3525 4471
rect 3200 4440 3525 4468
rect 3200 4428 3206 4440
rect 3513 4437 3525 4440
rect 3559 4437 3571 4471
rect 4080 4468 4108 4508
rect 5552 4508 5724 4536
rect 5074 4468 5080 4480
rect 4080 4440 5080 4468
rect 3513 4431 3571 4437
rect 5074 4428 5080 4440
rect 5132 4468 5138 4480
rect 5552 4468 5580 4508
rect 5718 4496 5724 4508
rect 5776 4536 5782 4548
rect 5828 4536 5856 4567
rect 5776 4508 5856 4536
rect 5776 4496 5782 4508
rect 5132 4440 5580 4468
rect 5132 4428 5138 4440
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 7006 4468 7012 4480
rect 5684 4440 7012 4468
rect 5684 4428 5690 4440
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7190 4468 7196 4480
rect 7151 4440 7196 4468
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4468 7435 4471
rect 8202 4468 8208 4480
rect 7423 4440 8208 4468
rect 7423 4437 7435 4440
rect 7377 4431 7435 4437
rect 8202 4428 8208 4440
rect 8260 4468 8266 4480
rect 8849 4471 8907 4477
rect 8849 4468 8861 4471
rect 8260 4440 8861 4468
rect 8260 4428 8266 4440
rect 8849 4437 8861 4440
rect 8895 4437 8907 4471
rect 8849 4431 8907 4437
rect 10919 4471 10977 4477
rect 10919 4437 10931 4471
rect 10965 4468 10977 4471
rect 11054 4468 11060 4480
rect 10965 4440 11060 4468
rect 10965 4437 10977 4440
rect 10919 4431 10977 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 14826 4468 14832 4480
rect 14231 4440 14832 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 4246 4264 4252 4276
rect 3108 4236 4108 4264
rect 4207 4236 4252 4264
rect 3108 4224 3114 4236
rect 4080 4196 4108 4236
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 6822 4264 6828 4276
rect 5224 4236 6828 4264
rect 5224 4224 5230 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 4080 4168 4660 4196
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 4632 4137 4660 4168
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 16666 4196 16672 4208
rect 4764 4168 16672 4196
rect 4764 4156 4770 4168
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 1728 4100 2881 4128
rect 1728 4088 1734 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5500 4100 5948 4128
rect 5500 4088 5506 4100
rect 1854 4060 1860 4072
rect 1815 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2225 4023 2283 4029
rect 2240 3992 2268 4023
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 3142 4069 3148 4072
rect 3136 4060 3148 4069
rect 2976 4032 3148 4060
rect 2976 3992 3004 4032
rect 3136 4023 3148 4032
rect 3142 4020 3148 4023
rect 3200 4020 3206 4072
rect 5920 4069 5948 4100
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7929 4131 7987 4137
rect 6972 4100 7017 4128
rect 6972 4088 6978 4100
rect 7929 4097 7941 4131
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 12434 4128 12440 4140
rect 11011 4100 12440 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4029 5963 4063
rect 7944 4060 7972 4091
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7944 4032 8217 4060
rect 5905 4023 5963 4029
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 2240 3964 3004 3992
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3961 4767 3995
rect 5626 3992 5632 4004
rect 5587 3964 5632 3992
rect 4709 3955 4767 3961
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 4724 3924 4752 3955
rect 5626 3952 5632 3964
rect 5684 3952 5690 4004
rect 7006 3992 7012 4004
rect 6967 3964 7012 3992
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11974 3992 11980 4004
rect 11112 3964 11157 3992
rect 11935 3964 11980 3992
rect 11112 3952 11118 3964
rect 11974 3952 11980 3964
rect 12032 3952 12038 4004
rect 2648 3896 4752 3924
rect 6089 3927 6147 3933
rect 2648 3884 2654 3896
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 8294 3924 8300 3936
rect 6135 3896 8300 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 13722 3924 13728 3936
rect 8435 3896 13728 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 3234 3720 3240 3732
rect 3195 3692 3240 3720
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7156 3692 7573 3720
rect 7156 3680 7162 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 8067 3723 8125 3729
rect 8067 3720 8079 3723
rect 7892 3692 8079 3720
rect 7892 3680 7898 3692
rect 8067 3689 8079 3692
rect 8113 3689 8125 3723
rect 8067 3683 8125 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 12526 3720 12532 3732
rect 8352 3692 12532 3720
rect 8352 3680 8358 3692
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 2124 3655 2182 3661
rect 2124 3621 2136 3655
rect 2170 3652 2182 3655
rect 3050 3652 3056 3664
rect 2170 3624 3056 3652
rect 2170 3621 2182 3624
rect 2124 3615 2182 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3651 3655 3709 3661
rect 3651 3621 3663 3655
rect 3697 3652 3709 3655
rect 4249 3655 4307 3661
rect 4249 3652 4261 3655
rect 3697 3624 4261 3652
rect 3697 3621 3709 3624
rect 3651 3615 3709 3621
rect 4249 3621 4261 3624
rect 4295 3621 4307 3655
rect 4249 3615 4307 3621
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 9766 3652 9772 3664
rect 5684 3624 9772 3652
rect 5684 3612 5690 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 2590 3544 2596 3596
rect 2648 3584 2654 3596
rect 3548 3587 3606 3593
rect 3548 3584 3560 3587
rect 2648 3556 3560 3584
rect 2648 3544 2654 3556
rect 3548 3553 3560 3556
rect 3594 3553 3606 3587
rect 5718 3584 5724 3596
rect 5679 3556 5724 3584
rect 3548 3547 3606 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 5988 3587 6046 3593
rect 5988 3553 6000 3587
rect 6034 3584 6046 3587
rect 7190 3584 7196 3596
rect 6034 3556 7196 3584
rect 6034 3553 6046 3556
rect 5988 3547 6046 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7374 3584 7380 3596
rect 7335 3556 7380 3584
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7742 3544 7748 3596
rect 7800 3584 7806 3596
rect 7964 3587 8022 3593
rect 7964 3584 7976 3587
rect 7800 3556 7976 3584
rect 7800 3544 7806 3556
rect 7964 3553 7976 3556
rect 8010 3553 8022 3587
rect 7964 3547 8022 3553
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1728 3488 1869 3516
rect 1728 3476 1734 3488
rect 1857 3485 1869 3488
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4154 3516 4160 3528
rect 4115 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 3804 3448 3832 3476
rect 4062 3448 4068 3460
rect 3804 3420 4068 3448
rect 4062 3408 4068 3420
rect 4120 3448 4126 3460
rect 4448 3448 4476 3479
rect 4120 3420 4476 3448
rect 4120 3408 4126 3420
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 3200 3148 3249 3176
rect 3200 3136 3206 3148
rect 3237 3145 3249 3148
rect 3283 3145 3295 3179
rect 3237 3139 3295 3145
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 12434 3176 12440 3188
rect 4212 3148 12440 3176
rect 4212 3136 4218 3148
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 7377 3111 7435 3117
rect 7377 3108 7389 3111
rect 2516 3080 7389 3108
rect 2516 2981 2544 3080
rect 7377 3077 7389 3080
rect 7423 3108 7435 3111
rect 10594 3108 10600 3120
rect 7423 3080 10600 3108
rect 7423 3077 7435 3080
rect 7377 3071 7435 3077
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 2740 3012 4200 3040
rect 2740 3000 2746 3012
rect 2501 2975 2559 2981
rect 2501 2941 2513 2975
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2648 2944 3065 2972
rect 2648 2932 2654 2944
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 3694 2972 3700 2984
rect 3655 2944 3700 2972
rect 3053 2935 3111 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 4080 2904 4108 2935
rect 3068 2876 4108 2904
rect 3068 2848 3096 2876
rect 2130 2796 2136 2848
rect 2188 2836 2194 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2188 2808 2697 2836
rect 2188 2796 2194 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 2685 2799 2743 2805
rect 3050 2796 3056 2848
rect 3108 2796 3114 2848
rect 4172 2836 4200 3012
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 4847 3043 4905 3049
rect 4847 3040 4859 3043
rect 4580 3012 4859 3040
rect 4580 3000 4586 3012
rect 4847 3009 4859 3012
rect 4893 3009 4905 3043
rect 4847 3003 4905 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 12526 3040 12532 3052
rect 5307 3012 12532 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4744 2975 4802 2981
rect 4744 2972 4756 2975
rect 4672 2944 4756 2972
rect 4672 2932 4678 2944
rect 4744 2941 4756 2944
rect 4790 2941 4802 2975
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 4744 2935 4802 2941
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 9766 2972 9772 2984
rect 9727 2944 9772 2972
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 4430 2904 4436 2916
rect 4391 2876 4436 2904
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 5350 2864 5356 2916
rect 5408 2904 5414 2916
rect 6273 2907 6331 2913
rect 5408 2876 5453 2904
rect 5408 2864 5414 2876
rect 6273 2873 6285 2907
rect 6319 2873 6331 2907
rect 6273 2867 6331 2873
rect 6288 2836 6316 2867
rect 4172 2808 6316 2836
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2836 10011 2839
rect 10594 2836 10600 2848
rect 9999 2808 10600 2836
rect 9999 2805 10011 2808
rect 9953 2799 10011 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2601 3663 2635
rect 3605 2595 3663 2601
rect 4249 2635 4307 2641
rect 4249 2601 4261 2635
rect 4295 2632 4307 2635
rect 4338 2632 4344 2644
rect 4295 2604 4344 2632
rect 4295 2601 4307 2604
rect 4249 2595 4307 2601
rect 3620 2564 3648 2595
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 5350 2592 5356 2644
rect 5408 2641 5414 2644
rect 5408 2635 5457 2641
rect 5408 2601 5411 2635
rect 5445 2601 5457 2635
rect 13078 2632 13084 2644
rect 5408 2595 5457 2601
rect 6932 2604 13084 2632
rect 5408 2592 5414 2595
rect 6932 2564 6960 2604
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 3620 2536 6960 2564
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7064 2536 7972 2564
rect 7064 2524 7070 2536
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 1929 2499 1987 2505
rect 1929 2496 1941 2499
rect 1452 2468 1941 2496
rect 1452 2456 1458 2468
rect 1929 2465 1941 2468
rect 1975 2465 1987 2499
rect 1929 2459 1987 2465
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 3421 2499 3479 2505
rect 3421 2496 3433 2499
rect 3384 2468 3433 2496
rect 3384 2456 3390 2468
rect 3421 2465 3433 2468
rect 3467 2465 3479 2499
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 3421 2459 3479 2465
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4430 2456 4436 2508
rect 4488 2496 4494 2508
rect 5296 2499 5354 2505
rect 5296 2496 5308 2499
rect 4488 2468 5308 2496
rect 4488 2456 4494 2468
rect 5296 2465 5308 2468
rect 5342 2496 5354 2499
rect 6273 2499 6331 2505
rect 5342 2468 6224 2496
rect 5342 2465 5354 2468
rect 5296 2459 5354 2465
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 6196 2360 6224 2468
rect 6273 2465 6285 2499
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6288 2428 6316 2459
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6880 2468 6929 2496
rect 6880 2456 6886 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7944 2505 7972 2536
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 7156 2468 7297 2496
rect 7156 2456 7162 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 6288 2400 7665 2428
rect 7653 2397 7665 2400
rect 7699 2428 7711 2431
rect 10502 2428 10508 2440
rect 7699 2400 10508 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 6196 2332 6592 2360
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6420 2264 6469 2292
rect 6420 2252 6426 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6564 2292 6592 2332
rect 7006 2292 7012 2304
rect 6564 2264 7012 2292
rect 6457 2255 6515 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 8113 2295 8171 2301
rect 8113 2261 8125 2295
rect 8159 2292 8171 2295
rect 10962 2292 10968 2304
rect 8159 2264 10968 2292
rect 8159 2261 8171 2264
rect 8113 2255 8171 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 7098 2088 7104 2100
rect 3292 2060 7104 2088
rect 3292 2048 3298 2060
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 10962 1300 10968 1352
rect 11020 1340 11026 1352
rect 12710 1340 12716 1352
rect 11020 1312 12716 1340
rect 11020 1300 11026 1312
rect 12710 1300 12716 1312
rect 12768 1300 12774 1352
<< via1 >>
rect 3424 7080 3476 7132
rect 8944 7080 8996 7132
rect 3056 6876 3108 6928
rect 7748 6876 7800 6928
rect 13084 6672 13136 6724
rect 13544 6672 13596 6724
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 204 6400 256 6452
rect 11704 6443 11756 6452
rect 1124 6332 1176 6384
rect 2596 6332 2648 6384
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 9128 6332 9180 6384
rect 11704 6409 11713 6443
rect 11713 6409 11747 6443
rect 11747 6409 11756 6443
rect 11704 6400 11756 6409
rect 15200 6332 15252 6384
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9680 6264 9732 6316
rect 10232 6264 10284 6316
rect 12164 6264 12216 6316
rect 16212 6264 16264 6316
rect 5080 6196 5132 6248
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 11152 6196 11204 6248
rect 11980 6196 12032 6248
rect 1676 6128 1728 6180
rect 2504 6060 2556 6112
rect 4528 6128 4580 6180
rect 5172 6171 5224 6180
rect 5172 6137 5181 6171
rect 5181 6137 5215 6171
rect 5215 6137 5224 6171
rect 5172 6128 5224 6137
rect 5356 6128 5408 6180
rect 3332 6060 3384 6112
rect 6920 6060 6972 6112
rect 7012 6060 7064 6112
rect 7380 6060 7432 6112
rect 8760 6128 8812 6180
rect 9220 6060 9272 6112
rect 10324 6171 10376 6180
rect 10324 6137 10333 6171
rect 10333 6137 10367 6171
rect 10367 6137 10376 6171
rect 10324 6128 10376 6137
rect 10508 6128 10560 6180
rect 12348 6128 12400 6180
rect 13912 6128 13964 6180
rect 14096 6128 14148 6180
rect 15108 6171 15160 6180
rect 15108 6137 15117 6171
rect 15117 6137 15151 6171
rect 15151 6137 15160 6171
rect 15108 6128 15160 6137
rect 15660 6060 15712 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 6276 5856 6328 5908
rect 1860 5831 1912 5840
rect 1860 5797 1869 5831
rect 1869 5797 1903 5831
rect 1903 5797 1912 5831
rect 1860 5788 1912 5797
rect 4620 5831 4672 5840
rect 4620 5797 4629 5831
rect 4629 5797 4663 5831
rect 4663 5797 4672 5831
rect 4620 5788 4672 5797
rect 4712 5831 4764 5840
rect 4712 5797 4721 5831
rect 4721 5797 4755 5831
rect 4755 5797 4764 5831
rect 8944 5856 8996 5908
rect 4712 5788 4764 5797
rect 6920 5788 6972 5840
rect 7748 5831 7800 5840
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 3332 5720 3384 5772
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 7748 5797 7757 5831
rect 7757 5797 7791 5831
rect 7791 5797 7800 5831
rect 7748 5788 7800 5797
rect 7840 5831 7892 5840
rect 7840 5797 7849 5831
rect 7849 5797 7883 5831
rect 7883 5797 7892 5831
rect 7840 5788 7892 5797
rect 8668 5788 8720 5840
rect 10140 5856 10192 5908
rect 10600 5856 10652 5908
rect 10692 5788 10744 5840
rect 14096 5856 14148 5908
rect 14188 5856 14240 5908
rect 14648 5856 14700 5908
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 10232 5763 10284 5772
rect 8668 5652 8720 5704
rect 10232 5729 10241 5763
rect 10241 5729 10275 5763
rect 10275 5729 10284 5763
rect 10232 5720 10284 5729
rect 7564 5584 7616 5636
rect 8300 5584 8352 5636
rect 12348 5763 12400 5772
rect 12348 5729 12366 5763
rect 12366 5729 12400 5763
rect 12348 5720 12400 5729
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 14004 5652 14056 5704
rect 2780 5516 2832 5568
rect 7748 5516 7800 5568
rect 14464 5584 14516 5636
rect 10416 5516 10468 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 2688 5312 2740 5364
rect 5356 5312 5408 5364
rect 1860 5244 1912 5296
rect 5080 5244 5132 5296
rect 7656 5312 7708 5364
rect 10324 5312 10376 5364
rect 13176 5355 13228 5364
rect 13176 5321 13185 5355
rect 13185 5321 13219 5355
rect 13219 5321 13228 5355
rect 13176 5312 13228 5321
rect 13636 5312 13688 5364
rect 12808 5244 12860 5296
rect 13728 5244 13780 5296
rect 664 5176 716 5228
rect 2136 5108 2188 5160
rect 2780 5108 2832 5160
rect 4252 5108 4304 5160
rect 3332 5040 3384 5092
rect 4620 5040 4672 5092
rect 8760 5176 8812 5228
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 5816 5108 5868 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 7748 5108 7800 5160
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 8668 5108 8720 5160
rect 10416 5108 10468 5160
rect 12716 5108 12768 5160
rect 15108 5176 15160 5228
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 6920 5040 6972 5092
rect 7012 5040 7064 5092
rect 7196 4972 7248 5024
rect 12440 4972 12492 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 2504 4768 2556 4820
rect 4712 4768 4764 4820
rect 5816 4768 5868 4820
rect 9220 4768 9272 4820
rect 2780 4632 2832 4684
rect 3240 4632 3292 4684
rect 4252 4700 4304 4752
rect 4620 4632 4672 4684
rect 7196 4700 7248 4752
rect 1676 4564 1728 4616
rect 7564 4632 7616 4684
rect 10600 4632 10652 4684
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 1768 4539 1820 4548
rect 1768 4505 1777 4539
rect 1777 4505 1811 4539
rect 1811 4505 1820 4539
rect 1768 4496 1820 4505
rect 3148 4428 3200 4480
rect 5080 4428 5132 4480
rect 5724 4496 5776 4548
rect 5632 4428 5684 4480
rect 7012 4428 7064 4480
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 8208 4428 8260 4480
rect 11060 4428 11112 4480
rect 14832 4428 14884 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 3056 4224 3108 4276
rect 4252 4267 4304 4276
rect 4252 4233 4261 4267
rect 4261 4233 4295 4267
rect 4295 4233 4304 4267
rect 4252 4224 4304 4233
rect 5172 4224 5224 4276
rect 6828 4224 6880 4276
rect 1676 4088 1728 4140
rect 4712 4156 4764 4208
rect 16672 4156 16724 4208
rect 5448 4088 5500 4140
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 1860 4020 1912 4029
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 3148 4063 3200 4072
rect 3148 4029 3182 4063
rect 3182 4029 3200 4063
rect 3148 4020 3200 4029
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 12440 4088 12492 4140
rect 5632 3995 5684 4004
rect 2596 3884 2648 3936
rect 5632 3961 5641 3995
rect 5641 3961 5675 3995
rect 5675 3961 5684 3995
rect 5632 3952 5684 3961
rect 7012 3995 7064 4004
rect 7012 3961 7021 3995
rect 7021 3961 7055 3995
rect 7055 3961 7064 3995
rect 7012 3952 7064 3961
rect 11060 3995 11112 4004
rect 11060 3961 11069 3995
rect 11069 3961 11103 3995
rect 11103 3961 11112 3995
rect 11980 3995 12032 4004
rect 11060 3952 11112 3961
rect 11980 3961 11989 3995
rect 11989 3961 12023 3995
rect 12023 3961 12032 3995
rect 11980 3952 12032 3961
rect 8300 3884 8352 3936
rect 13728 3884 13780 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 7104 3680 7156 3732
rect 7840 3680 7892 3732
rect 8300 3680 8352 3732
rect 12532 3680 12584 3732
rect 3056 3612 3108 3664
rect 5632 3612 5684 3664
rect 9772 3612 9824 3664
rect 2596 3544 2648 3596
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 7196 3544 7248 3596
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 7748 3544 7800 3596
rect 1676 3476 1728 3528
rect 3792 3476 3844 3528
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4068 3408 4120 3460
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 3148 3136 3200 3188
rect 4160 3136 4212 3188
rect 12440 3136 12492 3188
rect 10600 3068 10652 3120
rect 2688 3000 2740 3052
rect 2596 2932 2648 2984
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 2136 2796 2188 2848
rect 3056 2796 3108 2848
rect 4528 3000 4580 3052
rect 12532 3000 12584 3052
rect 4620 2932 4672 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 4436 2907 4488 2916
rect 4436 2873 4445 2907
rect 4445 2873 4479 2907
rect 4479 2873 4488 2907
rect 4436 2864 4488 2873
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 10600 2796 10652 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 4344 2592 4396 2644
rect 5356 2592 5408 2644
rect 13084 2592 13136 2644
rect 7012 2524 7064 2576
rect 1400 2456 1452 2508
rect 3332 2456 3384 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 4436 2456 4488 2508
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 6828 2456 6880 2508
rect 7104 2456 7156 2508
rect 10508 2388 10560 2440
rect 6368 2252 6420 2304
rect 7012 2252 7064 2304
rect 10968 2252 11020 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 3240 2048 3292 2100
rect 7104 2048 7156 2100
rect 10968 1300 11020 1352
rect 12716 1300 12768 1352
<< metal2 >>
rect 202 8520 258 9000
rect 662 8520 718 9000
rect 1122 8520 1178 9000
rect 1674 8520 1730 9000
rect 2134 8520 2190 9000
rect 2686 8520 2742 9000
rect 3146 8520 3202 9000
rect 3422 8664 3478 8673
rect 3422 8599 3478 8608
rect 216 6458 244 8520
rect 204 6452 256 6458
rect 204 6394 256 6400
rect 676 5234 704 8520
rect 1136 6390 1164 8520
rect 1124 6384 1176 6390
rect 1124 6326 1176 6332
rect 1688 6186 1716 8520
rect 1858 6216 1914 6225
rect 1676 6180 1728 6186
rect 1858 6151 1914 6160
rect 1676 6122 1728 6128
rect 1872 5846 1900 6151
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 2148 5710 2176 8520
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 664 5228 716 5234
rect 664 5170 716 5176
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1766 4584 1822 4593
rect 1688 4146 1716 4558
rect 1766 4519 1768 4528
rect 1820 4519 1822 4528
rect 1768 4490 1820 4496
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3534 1716 4082
rect 1872 4078 1900 5238
rect 2148 5166 2176 5646
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2516 4826 2544 6054
rect 2608 5250 2636 6326
rect 2700 5370 2728 8520
rect 3054 7848 3110 7857
rect 3054 7783 3110 7792
rect 3068 6934 3096 7783
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5409 2820 5510
rect 2778 5400 2834 5409
rect 2688 5364 2740 5370
rect 2778 5335 2834 5344
rect 2688 5306 2740 5312
rect 2608 5222 2728 5250
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1412 1329 1440 2450
rect 1688 2446 1716 3470
rect 1872 2961 1900 4014
rect 2608 3942 2636 4014
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2608 3602 2636 3878
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2608 2990 2636 3538
rect 2700 3058 2728 5222
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4690 2820 5102
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3160 4570 3188 8520
rect 3436 7138 3464 8599
rect 3698 8520 3754 9000
rect 4158 8520 4214 9000
rect 4618 8520 4674 9000
rect 5170 8520 5226 9000
rect 5630 8520 5686 9000
rect 6182 8520 6238 9000
rect 6642 8520 6698 9000
rect 7194 8520 7250 9000
rect 7654 8520 7710 9000
rect 8206 8520 8262 9000
rect 8666 8520 8722 9000
rect 9126 8520 9182 9000
rect 9678 8520 9734 9000
rect 10138 8520 10194 9000
rect 10690 8520 10746 9000
rect 11150 8520 11206 9000
rect 11702 8520 11758 9000
rect 12162 8520 12218 9000
rect 12714 8520 12770 9000
rect 13174 8520 13230 9000
rect 13634 8520 13690 9000
rect 14186 8520 14242 9000
rect 14646 8520 14702 9000
rect 15198 8520 15254 9000
rect 15658 8520 15714 9000
rect 16210 8520 16266 9000
rect 16670 8520 16726 9000
rect 3424 7132 3476 7138
rect 3424 7074 3476 7080
rect 3712 6746 3740 8520
rect 4172 7834 4200 8520
rect 4172 7806 4384 7834
rect 4158 7032 4214 7041
rect 4158 6967 4214 6976
rect 3712 6718 3832 6746
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5778 3372 6054
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3344 5098 3372 5714
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3068 4542 3188 4570
rect 3068 4282 3096 4542
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 3160 4078 3188 4422
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3146 3768 3202 3777
rect 3252 3738 3280 4626
rect 3146 3703 3202 3712
rect 3240 3732 3292 3738
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2596 2984 2648 2990
rect 1858 2952 1914 2961
rect 2596 2926 2648 2932
rect 1858 2887 1914 2896
rect 3068 2854 3096 3606
rect 3160 3194 3188 3703
rect 3240 3674 3292 3680
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1398 1320 1454 1329
rect 1398 1255 1454 1264
rect 1688 513 1716 2382
rect 1674 504 1730 513
rect 2148 480 2176 2790
rect 3068 2650 3096 2790
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3344 2514 3372 5034
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3804 3534 3832 6718
rect 4172 6322 4200 6967
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4252 5160 4304 5166
rect 4252 5102 4304 5108
rect 4264 4758 4292 5102
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4264 4282 4292 4694
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3700 2984 3752 2990
rect 3698 2952 3700 2961
rect 3752 2952 3754 2961
rect 3698 2887 3754 2896
rect 4080 2514 4108 3402
rect 4172 3194 4200 3470
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4356 2650 4384 7806
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4540 3058 4568 6122
rect 4632 5846 4660 8520
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4620 5092 4672 5098
rect 4724 5080 4752 5782
rect 5092 5302 5120 6190
rect 5184 6186 5212 8520
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 5368 5370 5396 6122
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5080 5296 5132 5302
rect 5132 5244 5212 5250
rect 5080 5238 5212 5244
rect 5092 5222 5212 5238
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4672 5052 4752 5080
rect 4620 5034 4672 5040
rect 4632 4690 4660 5034
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4632 2990 4660 4626
rect 4724 4214 4752 4762
rect 5092 4486 5120 5102
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5184 4282 5212 5222
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 5460 4146 5488 5646
rect 5644 4486 5672 8520
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 5166 5856 6190
rect 6196 6100 6224 8520
rect 6656 6338 6684 8520
rect 7208 7834 7236 8520
rect 7116 7806 7236 7834
rect 6656 6310 7052 6338
rect 7024 6118 7052 6310
rect 6920 6112 6972 6118
rect 6196 6072 6316 6100
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 6288 5914 6316 6072
rect 6920 6054 6972 6060
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6932 5846 6960 6054
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 5828 4826 5856 5102
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5644 3670 5672 3946
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5736 3602 5764 4490
rect 6840 4282 6868 5102
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6840 2990 6868 4218
rect 6932 4146 6960 5034
rect 7024 4486 7052 5034
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4448 2514 4476 2858
rect 5368 2650 5396 2858
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 6840 2514 6868 2926
rect 7024 2582 7052 3946
rect 7116 3738 7144 7806
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 6118 7420 6258
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 5030 7236 5102
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4758 7236 4966
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7208 3602 7236 4422
rect 7392 3602 7420 6054
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 4690 7604 5578
rect 7668 5370 7696 8520
rect 7748 6928 7800 6934
rect 7748 6870 7800 6876
rect 7760 5846 7788 6870
rect 8220 6066 8248 8520
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8220 6038 8340 6066
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7760 5166 7788 5510
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7760 3602 7788 5102
rect 7852 3738 7880 5782
rect 8312 5642 8340 6038
rect 8680 5846 8708 8520
rect 8944 7132 8996 7138
rect 8944 7074 8996 7080
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8680 5166 8708 5646
rect 8772 5234 8800 6122
rect 8956 5914 8984 7074
rect 9140 6390 9168 8520
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 9692 6322 9720 8520
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9048 5778 9076 6258
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8220 4486 8248 5102
rect 9232 4826 9260 6054
rect 10152 5914 10180 8520
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10244 5778 10272 6258
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10336 5370 10364 6122
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10428 5166 10456 5510
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8312 3738 8340 3878
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7024 2310 7052 2518
rect 7116 2514 7144 3334
rect 7208 2990 7236 3538
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 9784 2990 9812 3606
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3238 2136 3294 2145
rect 3421 2128 3717 2148
rect 3238 2071 3240 2080
rect 3292 2071 3294 2080
rect 3240 2042 3292 2048
rect 6380 480 6408 2246
rect 7116 2106 7144 2450
rect 10520 2446 10548 6122
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10612 4690 10640 5850
rect 10704 5846 10732 8520
rect 11164 6254 11192 8520
rect 11716 6458 11744 8520
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 12176 6322 12204 8520
rect 12438 6352 12494 6361
rect 12164 6316 12216 6322
rect 12438 6287 12494 6296
rect 12164 6258 12216 6264
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 3126 10640 4626
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4010 11100 4422
rect 11992 4010 12020 6190
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12360 5778 12388 6122
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12452 5030 12480 6287
rect 12530 5264 12586 5273
rect 12530 5199 12586 5208
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 12452 3505 12480 4082
rect 12544 3738 12572 5199
rect 12728 5166 12756 8520
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12820 5302 12848 5646
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12438 3496 12494 3505
rect 12438 3431 12494 3440
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 10612 480 10640 2790
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 12452 2417 12480 3130
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12438 2408 12494 2417
rect 12438 2343 12494 2352
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1358 11008 2246
rect 12544 1465 12572 2994
rect 13096 2650 13124 6666
rect 13188 5370 13216 8520
rect 13648 7834 13676 8520
rect 13726 8392 13782 8401
rect 13726 8327 13782 8336
rect 13556 7806 13676 7834
rect 13556 6730 13584 7806
rect 13740 7698 13768 8327
rect 13648 7670 13768 7698
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13648 5370 13676 7670
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13740 5302 13768 7375
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13924 5166 13952 6122
rect 14108 5914 14136 6122
rect 14200 5914 14228 8520
rect 14660 5914 14688 8520
rect 15212 6390 15240 8520
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 14016 4690 14044 5646
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14476 5166 14504 5578
rect 15120 5234 15148 6122
rect 15672 6118 15700 8520
rect 16224 6322 16252 8520
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14832 4480 14884 4486
rect 13726 4448 13782 4457
rect 13282 4380 13578 4400
rect 14832 4422 14884 4428
rect 13726 4383 13782 4392
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13740 3942 13768 4383
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 12530 1456 12586 1465
rect 12530 1391 12586 1400
rect 10968 1352 11020 1358
rect 10968 1294 11020 1300
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 12728 513 12756 1294
rect 12714 504 12770 513
rect 1674 439 1730 448
rect 2134 0 2190 480
rect 6366 0 6422 480
rect 10598 0 10654 480
rect 14844 480 14872 4422
rect 16684 4214 16712 8520
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 12714 439 12770 448
rect 14830 0 14886 480
<< via2 >>
rect 3422 8608 3478 8664
rect 1858 6160 1914 6216
rect 1766 4548 1822 4584
rect 1766 4528 1768 4548
rect 1768 4528 1820 4548
rect 1820 4528 1822 4548
rect 3054 7792 3110 7848
rect 2778 5344 2834 5400
rect 4158 6976 4214 7032
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3146 3712 3202 3768
rect 1858 2896 1914 2952
rect 1398 1264 1454 1320
rect 1674 448 1730 504
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3698 2932 3700 2952
rect 3700 2932 3752 2952
rect 3752 2932 3754 2952
rect 3698 2896 3754 2932
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3238 2100 3294 2136
rect 3238 2080 3240 2100
rect 3240 2080 3292 2100
rect 3292 2080 3294 2100
rect 12438 6296 12494 6352
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 12530 5208 12586 5264
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 12438 3440 12494 3496
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 12438 2352 12494 2408
rect 13726 8336 13782 8392
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13726 7384 13782 7440
rect 13726 4392 13782 4448
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 12530 1400 12586 1456
rect 12714 448 12770 504
<< metal3 >>
rect 0 8666 480 8696
rect 3417 8666 3483 8669
rect 0 8664 3483 8666
rect 0 8608 3422 8664
rect 3478 8608 3483 8664
rect 0 8606 3483 8608
rect 0 8576 480 8606
rect 3417 8603 3483 8606
rect 13721 8394 13787 8397
rect 16520 8394 17000 8424
rect 13721 8392 17000 8394
rect 13721 8336 13726 8392
rect 13782 8336 17000 8392
rect 13721 8334 17000 8336
rect 13721 8331 13787 8334
rect 16520 8304 17000 8334
rect 0 7850 480 7880
rect 3049 7850 3115 7853
rect 0 7848 3115 7850
rect 0 7792 3054 7848
rect 3110 7792 3115 7848
rect 0 7790 3115 7792
rect 0 7760 480 7790
rect 3049 7787 3115 7790
rect 13721 7442 13787 7445
rect 16520 7442 17000 7472
rect 13721 7440 17000 7442
rect 13721 7384 13726 7440
rect 13782 7384 17000 7440
rect 13721 7382 17000 7384
rect 13721 7379 13787 7382
rect 16520 7352 17000 7382
rect 0 7034 480 7064
rect 4153 7034 4219 7037
rect 0 7032 4219 7034
rect 0 6976 4158 7032
rect 4214 6976 4219 7032
rect 0 6974 4219 6976
rect 0 6944 480 6974
rect 4153 6971 4219 6974
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 16520 6490 17000 6520
rect 13678 6430 17000 6490
rect 12433 6354 12499 6357
rect 13678 6354 13738 6430
rect 16520 6400 17000 6430
rect 12433 6352 13738 6354
rect 12433 6296 12438 6352
rect 12494 6296 13738 6352
rect 12433 6294 13738 6296
rect 12433 6291 12499 6294
rect 0 6218 480 6248
rect 1853 6218 1919 6221
rect 0 6216 1919 6218
rect 0 6160 1858 6216
rect 1914 6160 1919 6216
rect 0 6158 1919 6160
rect 0 6128 480 6158
rect 1853 6155 1919 6158
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 3409 5472 3729 5473
rect 0 5402 480 5432
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 2773 5402 2839 5405
rect 16520 5402 17000 5432
rect 0 5400 2839 5402
rect 0 5344 2778 5400
rect 2834 5344 2839 5400
rect 0 5342 2839 5344
rect 0 5312 480 5342
rect 2773 5339 2839 5342
rect 13678 5342 17000 5402
rect 12525 5266 12591 5269
rect 13678 5266 13738 5342
rect 16520 5312 17000 5342
rect 12525 5264 13738 5266
rect 12525 5208 12530 5264
rect 12586 5208 13738 5264
rect 12525 5206 13738 5208
rect 12525 5203 12591 5206
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 0 4586 480 4616
rect 1761 4586 1827 4589
rect 0 4584 1827 4586
rect 0 4528 1766 4584
rect 1822 4528 1827 4584
rect 0 4526 1827 4528
rect 0 4496 480 4526
rect 1761 4523 1827 4526
rect 13721 4450 13787 4453
rect 16520 4450 17000 4480
rect 13721 4448 17000 4450
rect 13721 4392 13726 4448
rect 13782 4392 17000 4448
rect 13721 4390 17000 4392
rect 13721 4387 13787 4390
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 16520 4360 17000 4390
rect 13270 4319 13590 4320
rect 5874 3840 6194 3841
rect 0 3770 480 3800
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3141 3770 3207 3773
rect 0 3768 3207 3770
rect 0 3712 3146 3768
rect 3202 3712 3207 3768
rect 0 3710 3207 3712
rect 0 3680 480 3710
rect 3141 3707 3207 3710
rect 12433 3498 12499 3501
rect 16520 3498 17000 3528
rect 12433 3496 17000 3498
rect 12433 3440 12438 3496
rect 12494 3440 17000 3496
rect 12433 3438 17000 3440
rect 12433 3435 12499 3438
rect 16520 3408 17000 3438
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 0 2954 480 2984
rect 1853 2954 1919 2957
rect 3693 2954 3759 2957
rect 0 2952 3759 2954
rect 0 2896 1858 2952
rect 1914 2896 3698 2952
rect 3754 2896 3759 2952
rect 0 2894 3759 2896
rect 0 2864 480 2894
rect 1853 2891 1919 2894
rect 3693 2891 3759 2894
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 12433 2410 12499 2413
rect 16520 2410 17000 2440
rect 12433 2408 17000 2410
rect 12433 2352 12438 2408
rect 12494 2352 17000 2408
rect 12433 2350 17000 2352
rect 12433 2347 12499 2350
rect 16520 2320 17000 2350
rect 3409 2208 3729 2209
rect 0 2138 480 2168
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 3233 2138 3299 2141
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 2048 480 2078
rect 3233 2075 3299 2078
rect 12525 1458 12591 1461
rect 16520 1458 17000 1488
rect 12525 1456 17000 1458
rect 12525 1400 12530 1456
rect 12586 1400 17000 1456
rect 12525 1398 17000 1400
rect 12525 1395 12591 1398
rect 16520 1368 17000 1398
rect 0 1322 480 1352
rect 1393 1322 1459 1325
rect 0 1320 1459 1322
rect 0 1264 1398 1320
rect 1454 1264 1459 1320
rect 0 1262 1459 1264
rect 0 1232 480 1262
rect 1393 1259 1459 1262
rect 0 506 480 536
rect 1669 506 1735 509
rect 0 504 1735 506
rect 0 448 1674 504
rect 1730 448 1735 504
rect 0 446 1735 448
rect 0 416 480 446
rect 1669 443 1735 446
rect 12709 506 12775 509
rect 16520 506 17000 536
rect 12709 504 17000 506
rect 12709 448 12714 504
rect 12770 448 17000 504
rect 12709 446 17000 448
rect 12709 443 12775 446
rect 16520 416 17000 446
<< via3 >>
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 6560 3729 6576
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 6016 6195 6576
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 6560 8660 6576
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 6016 11125 6576
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 13270 6560 13590 6576
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__buf_2  _02_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1656 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1605641404
transform 1 0 3036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1605641404
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22
timestamp 1605641404
transform 1 0 3128 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1605641404
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_25
timestamp 1605641404
transform 1 0 3404 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5152 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4416 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1605641404
transform 1 0 5520 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1605641404
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1605641404
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _01_
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1605641404
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1605641404
transform 1 0 7912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1605641404
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_78
timestamp 1605641404
transform 1 0 8280 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_71
timestamp 1605641404
transform 1 0 7636 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_83
timestamp 1605641404
transform 1 0 8740 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1605641404
transform 1 0 9752 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1605641404
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_91
timestamp 1605641404
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1605641404
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1605641404
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1605641404
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1605641404
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1840 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1605641404
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_23
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1605641404
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1605641404
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1605641404
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1605641404
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1605641404
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _00_
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 7912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1605641404
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_24
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1605641404
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1605641404
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1605641404
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1605641404
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1605641404
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_25
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1605641404
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2852 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1605641404
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 4508 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1605641404
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1605641404
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1605641404
transform 1 0 5888 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_26
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_56
timestamp 1605641404
transform 1 0 6256 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1605641404
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1605641404
transform 1 0 8188 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1605641404
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1605641404
transform 1 0 8556 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1605641404
transform 1 0 9660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 10856 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_3_105
timestamp 1605641404
transform 1 0 10764 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_27
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1605641404
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1605641404
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1605641404
transform 1 0 14628 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1605641404
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1605641404
transform 1 0 1564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2116 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1605641404
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5796 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1605641404
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7452 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1605641404
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 10764 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_108
timestamp 1605641404
transform 1 0 11040 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_120
timestamp 1605641404
transform 1 0 12144 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1605641404
transform 1 0 13248 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1605641404
transform 1 0 13984 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_144
timestamp 1605641404
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1605641404
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1605641404
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 2300 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1605641404
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_22
timestamp 1605641404
transform 1 0 3128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_37
timestamp 1605641404
transform 1 0 4508 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1605641404
transform 1 0 8832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1605641404
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1605641404
transform 1 0 9384 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 10212 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1605641404
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1605641404
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_102
timestamp 1605641404
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1605641404
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1605641404
transform 1 0 12972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_133
timestamp 1605641404
transform 1 0 13340 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1605641404
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1605641404
transform 1 0 14444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_143
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1605641404
transform 1 0 14812 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1605641404
transform 1 0 1932 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 1748 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1605641404
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1605641404
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1605641404
transform 1 0 3128 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 4048 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1605641404
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_20
timestamp 1605641404
transform 1 0 2944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_26
timestamp 1605641404
transform 1 0 3496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1605641404
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 1605641404
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 4508 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1605641404
transform 1 0 5428 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_35
timestamp 1605641404
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_50
timestamp 1605641404
transform 1 0 5704 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1605641404
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 6900 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_56
timestamp 1605641404
transform 1 0 6256 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 7636 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 8280 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1605641404
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1605641404
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1605641404
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1605641404
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1605641404
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1605641404
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1605641404
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1605641404
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1605641404
transform 1 0 9660 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1605641404
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1605641404
transform 1 0 11500 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 10764 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_6_103
timestamp 1605641404
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_111
timestamp 1605641404
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_117
timestamp 1605641404
transform 1 0 11868 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 12696 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1605641404
transform 1 0 12236 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 12604 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1605641404
transform 1 0 12512 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_118
timestamp 1605641404
transform 1 0 11960 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1605641404
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1605641404
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1605641404
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 13984 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_6_139
timestamp 1605641404
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1605641404
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1605641404
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1605641404
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1605641404
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_156
timestamp 1605641404
transform 1 0 15456 0 1 5984
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 2864 480 2984 6 IO_ISOL_N
port 0 nsew default input
rlabel metal3 s 0 1232 480 1352 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 2048 480 2168 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 16520 416 17000 536 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 3 nsew default tristate
rlabel metal2 s 13634 8520 13690 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 4 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 5 nsew default tristate
rlabel metal3 s 0 4496 480 4616 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 6 nsew default tristate
rlabel metal3 s 0 5312 480 5432 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 7 nsew default tristate
rlabel metal2 s 14186 8520 14242 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 8 nsew default tristate
rlabel metal2 s 14646 8520 14702 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 9 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 10 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 11 nsew default tristate
rlabel metal3 s 16520 1368 17000 1488 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 12 nsew default input
rlabel metal3 s 0 6128 480 6248 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 13 nsew default input
rlabel metal3 s 16520 2320 17000 2440 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 14 nsew default input
rlabel metal3 s 0 6944 480 7064 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 15 nsew default input
rlabel metal2 s 15198 8520 15254 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 16 nsew default input
rlabel metal3 s 0 7760 480 7880 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 17 nsew default input
rlabel metal2 s 15658 8520 15714 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 18 nsew default input
rlabel metal3 s 16520 3408 17000 3528 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 19 nsew default input
rlabel metal2 s 16210 8520 16266 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 20 nsew default input
rlabel metal3 s 16520 4360 17000 4480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 21 nsew default tristate
rlabel metal2 s 16670 8520 16726 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 22 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 23 nsew default tristate
rlabel metal3 s 16520 5312 17000 5432 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 24 nsew default tristate
rlabel metal3 s 16520 6400 17000 6520 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 25 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 26 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 27 nsew default tristate
rlabel metal3 s 16520 7352 17000 7472 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 28 nsew default tristate
rlabel metal3 s 16520 8304 17000 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 29 nsew default tristate
rlabel metal3 s 0 416 480 536 6 prog_clk
port 30 nsew default input
rlabel metal2 s 662 8520 718 9000 6 top_width_0_height_0__pin_0_
port 31 nsew default input
rlabel metal2 s 7654 8520 7710 9000 6 top_width_0_height_0__pin_10_
port 32 nsew default input
rlabel metal2 s 8206 8520 8262 9000 6 top_width_0_height_0__pin_11_lower
port 33 nsew default tristate
rlabel metal2 s 8666 8520 8722 9000 6 top_width_0_height_0__pin_11_upper
port 34 nsew default tristate
rlabel metal2 s 9126 8520 9182 9000 6 top_width_0_height_0__pin_12_
port 35 nsew default input
rlabel metal2 s 9678 8520 9734 9000 6 top_width_0_height_0__pin_13_lower
port 36 nsew default tristate
rlabel metal2 s 10138 8520 10194 9000 6 top_width_0_height_0__pin_13_upper
port 37 nsew default tristate
rlabel metal2 s 10690 8520 10746 9000 6 top_width_0_height_0__pin_14_
port 38 nsew default input
rlabel metal2 s 11150 8520 11206 9000 6 top_width_0_height_0__pin_15_lower
port 39 nsew default tristate
rlabel metal2 s 11702 8520 11758 9000 6 top_width_0_height_0__pin_15_upper
port 40 nsew default tristate
rlabel metal2 s 12162 8520 12218 9000 6 top_width_0_height_0__pin_16_
port 41 nsew default input
rlabel metal2 s 12714 8520 12770 9000 6 top_width_0_height_0__pin_17_lower
port 42 nsew default tristate
rlabel metal2 s 13174 8520 13230 9000 6 top_width_0_height_0__pin_17_upper
port 43 nsew default tristate
rlabel metal2 s 1122 8520 1178 9000 6 top_width_0_height_0__pin_1_lower
port 44 nsew default tristate
rlabel metal2 s 202 8520 258 9000 6 top_width_0_height_0__pin_1_upper
port 45 nsew default tristate
rlabel metal2 s 1674 8520 1730 9000 6 top_width_0_height_0__pin_2_
port 46 nsew default input
rlabel metal2 s 2134 8520 2190 9000 6 top_width_0_height_0__pin_3_lower
port 47 nsew default tristate
rlabel metal2 s 2686 8520 2742 9000 6 top_width_0_height_0__pin_3_upper
port 48 nsew default tristate
rlabel metal2 s 3146 8520 3202 9000 6 top_width_0_height_0__pin_4_
port 49 nsew default input
rlabel metal2 s 3698 8520 3754 9000 6 top_width_0_height_0__pin_5_lower
port 50 nsew default tristate
rlabel metal2 s 4158 8520 4214 9000 6 top_width_0_height_0__pin_5_upper
port 51 nsew default tristate
rlabel metal2 s 4618 8520 4674 9000 6 top_width_0_height_0__pin_6_
port 52 nsew default input
rlabel metal2 s 5170 8520 5226 9000 6 top_width_0_height_0__pin_7_lower
port 53 nsew default tristate
rlabel metal2 s 5630 8520 5686 9000 6 top_width_0_height_0__pin_7_upper
port 54 nsew default tristate
rlabel metal2 s 6182 8520 6238 9000 6 top_width_0_height_0__pin_8_
port 55 nsew default input
rlabel metal2 s 6642 8520 6698 9000 6 top_width_0_height_0__pin_9_lower
port 56 nsew default tristate
rlabel metal2 s 7194 8520 7250 9000 6 top_width_0_height_0__pin_9_upper
port 57 nsew default tristate
rlabel metal4 s 3409 2128 3729 6576 6 VPWR
port 58 nsew default input
rlabel metal4 s 5875 2128 6195 6576 6 VGND
port 59 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 9000
<< end >>
