magic
tech sky130A
magscale 1 2
timestamp 1605013573
<< viali >>
rect 22549 20961 22583 20995
rect 22293 20893 22327 20927
rect 23673 20757 23707 20791
rect 21741 20553 21775 20587
rect 22385 20553 22419 20587
rect 13645 20349 13679 20383
rect 20361 20349 20395 20383
rect 26065 20349 26099 20383
rect 13553 20281 13587 20315
rect 13890 20281 13924 20315
rect 20269 20281 20303 20315
rect 20606 20281 20640 20315
rect 22753 20281 22787 20315
rect 15025 20213 15059 20247
rect 26249 20213 26283 20247
rect 26709 20213 26743 20247
rect 13645 20009 13679 20043
rect 19717 20009 19751 20043
rect 20453 20009 20487 20043
rect 21557 20009 21591 20043
rect 18582 19941 18616 19975
rect 23745 19873 23779 19907
rect 18337 19805 18371 19839
rect 23489 19805 23523 19839
rect 24869 19669 24903 19703
rect 19257 19329 19291 19363
rect 8585 19261 8619 19295
rect 14565 19261 14599 19295
rect 15117 19261 15151 19295
rect 17417 19261 17451 19295
rect 24869 19261 24903 19295
rect 8493 19193 8527 19227
rect 8830 19193 8864 19227
rect 15362 19193 15396 19227
rect 18613 19193 18647 19227
rect 19165 19193 19199 19227
rect 24777 19193 24811 19227
rect 25114 19193 25148 19227
rect 9965 19125 9999 19159
rect 14933 19125 14967 19159
rect 16497 19125 16531 19159
rect 17877 19125 17911 19159
rect 18705 19125 18739 19159
rect 19073 19125 19107 19159
rect 23857 19125 23891 19159
rect 24317 19125 24351 19159
rect 26249 19125 26283 19159
rect 14105 18921 14139 18955
rect 17877 18921 17911 18955
rect 18797 18921 18831 18955
rect 18889 18921 18923 18955
rect 21281 18921 21315 18955
rect 23949 18921 23983 18955
rect 18337 18853 18371 18887
rect 4333 18785 4367 18819
rect 8677 18785 8711 18819
rect 10241 18785 10275 18819
rect 10497 18785 10531 18819
rect 12981 18785 13015 18819
rect 19257 18785 19291 18819
rect 23213 18785 23247 18819
rect 23305 18785 23339 18819
rect 1777 18717 1811 18751
rect 4077 18717 4111 18751
rect 12725 18717 12759 18751
rect 19349 18717 19383 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 21557 18717 21591 18751
rect 23489 18717 23523 18751
rect 2237 18581 2271 18615
rect 5457 18581 5491 18615
rect 7205 18581 7239 18615
rect 11621 18581 11655 18615
rect 20453 18581 20487 18615
rect 20913 18581 20947 18615
rect 22845 18581 22879 18615
rect 24961 18581 24995 18615
rect 4445 18377 4479 18411
rect 6561 18377 6595 18411
rect 8493 18377 8527 18411
rect 10701 18377 10735 18411
rect 12817 18377 12851 18411
rect 17877 18377 17911 18411
rect 18889 18377 18923 18411
rect 19901 18377 19935 18411
rect 20269 18377 20303 18411
rect 21557 18377 21591 18411
rect 21833 18377 21867 18411
rect 22385 18377 22419 18411
rect 23673 18377 23707 18411
rect 3249 18309 3283 18343
rect 4169 18309 4203 18343
rect 13093 18309 13127 18343
rect 14289 18309 14323 18343
rect 18337 18309 18371 18343
rect 20453 18309 20487 18343
rect 22753 18309 22787 18343
rect 7113 18241 7147 18275
rect 14841 18241 14875 18275
rect 19441 18241 19475 18275
rect 21005 18241 21039 18275
rect 24225 18241 24259 18275
rect 25697 18241 25731 18275
rect 1869 18173 1903 18207
rect 14657 18173 14691 18207
rect 20821 18173 20855 18207
rect 23489 18173 23523 18207
rect 24133 18173 24167 18207
rect 25796 18173 25830 18207
rect 1777 18105 1811 18139
rect 2136 18105 2170 18139
rect 7380 18105 7414 18139
rect 14749 18105 14783 18139
rect 23121 18105 23155 18139
rect 24041 18105 24075 18139
rect 26034 18105 26068 18139
rect 10241 18037 10275 18071
rect 13829 18037 13863 18071
rect 14197 18037 14231 18071
rect 18705 18037 18739 18071
rect 19257 18037 19291 18071
rect 19349 18037 19383 18071
rect 20913 18037 20947 18071
rect 27169 18037 27203 18071
rect 2237 17833 2271 17867
rect 12633 17833 12667 17867
rect 18613 17833 18647 17867
rect 19257 17833 19291 17867
rect 20545 17833 20579 17867
rect 21189 17833 21223 17867
rect 22109 17833 22143 17867
rect 22937 17833 22971 17867
rect 23213 17833 23247 17867
rect 5886 17765 5920 17799
rect 16396 17765 16430 17799
rect 18981 17765 19015 17799
rect 22201 17765 22235 17799
rect 2329 17697 2363 17731
rect 5641 17697 5675 17731
rect 10517 17697 10551 17731
rect 14013 17697 14047 17731
rect 16129 17697 16163 17731
rect 19625 17697 19659 17731
rect 23581 17697 23615 17731
rect 23673 17697 23707 17731
rect 2513 17629 2547 17663
rect 10609 17629 10643 17663
rect 10701 17629 10735 17663
rect 14105 17629 14139 17663
rect 14197 17629 14231 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 23857 17629 23891 17663
rect 1777 17493 1811 17527
rect 1869 17493 1903 17527
rect 2881 17493 2915 17527
rect 4445 17493 4479 17527
rect 4721 17493 4755 17527
rect 7021 17493 7055 17527
rect 9965 17493 9999 17527
rect 10149 17493 10183 17527
rect 13645 17493 13679 17527
rect 14749 17493 14783 17527
rect 17509 17493 17543 17527
rect 24225 17493 24259 17527
rect 25789 17493 25823 17527
rect 1869 17289 1903 17323
rect 2973 17289 3007 17323
rect 3801 17289 3835 17323
rect 5641 17289 5675 17323
rect 13461 17289 13495 17323
rect 15301 17289 15335 17323
rect 16221 17289 16255 17323
rect 18521 17289 18555 17323
rect 18889 17289 18923 17323
rect 19349 17289 19383 17323
rect 19441 17289 19475 17323
rect 24777 17289 24811 17323
rect 4261 17221 4295 17255
rect 13093 17221 13127 17255
rect 14289 17221 14323 17255
rect 23673 17221 23707 17255
rect 2421 17153 2455 17187
rect 2605 17153 2639 17187
rect 4813 17153 4847 17187
rect 4997 17153 5031 17187
rect 6009 17153 6043 17187
rect 9505 17153 9539 17187
rect 10425 17153 10459 17187
rect 10517 17153 10551 17187
rect 14841 17153 14875 17187
rect 16497 17153 16531 17187
rect 19993 17153 20027 17187
rect 22477 17153 22511 17187
rect 22661 17153 22695 17187
rect 24133 17153 24167 17187
rect 24317 17153 24351 17187
rect 25881 17153 25915 17187
rect 2329 17085 2363 17119
rect 9873 17085 9907 17119
rect 11069 17085 11103 17119
rect 22385 17085 22419 17119
rect 25973 17085 26007 17119
rect 26240 17085 26274 17119
rect 4721 17017 4755 17051
rect 9137 17017 9171 17051
rect 10333 17017 10367 17051
rect 13829 17017 13863 17051
rect 20821 17017 20855 17051
rect 21925 17017 21959 17051
rect 23213 17017 23247 17051
rect 24041 17017 24075 17051
rect 25053 17017 25087 17051
rect 1961 16949 1995 16983
rect 3433 16949 3467 16983
rect 4353 16949 4387 16983
rect 9965 16949 9999 16983
rect 14197 16949 14231 16983
rect 14657 16949 14691 16983
rect 14749 16949 14783 16983
rect 19809 16949 19843 16983
rect 19901 16949 19935 16983
rect 20453 16949 20487 16983
rect 22017 16949 22051 16983
rect 27353 16949 27387 16983
rect 1685 16745 1719 16779
rect 1961 16745 1995 16779
rect 2421 16745 2455 16779
rect 4077 16745 4111 16779
rect 10241 16745 10275 16779
rect 10425 16745 10459 16779
rect 10793 16745 10827 16779
rect 13185 16745 13219 16779
rect 14013 16745 14047 16779
rect 19533 16745 19567 16779
rect 22109 16745 22143 16779
rect 23213 16745 23247 16779
rect 24317 16745 24351 16779
rect 11989 16677 12023 16711
rect 23121 16677 23155 16711
rect 2329 16609 2363 16643
rect 4445 16609 4479 16643
rect 7205 16609 7239 16643
rect 13553 16609 13587 16643
rect 14105 16609 14139 16643
rect 18153 16609 18187 16643
rect 18420 16609 18454 16643
rect 20177 16609 20211 16643
rect 23581 16609 23615 16643
rect 26525 16609 26559 16643
rect 2605 16541 2639 16575
rect 4537 16541 4571 16575
rect 4629 16541 4663 16575
rect 7297 16541 7331 16575
rect 7389 16541 7423 16575
rect 10885 16541 10919 16575
rect 10977 16541 11011 16575
rect 14289 16541 14323 16575
rect 23673 16541 23707 16575
rect 23857 16541 23891 16575
rect 3065 16473 3099 16507
rect 3433 16405 3467 16439
rect 6837 16405 6871 16439
rect 8953 16405 8987 16439
rect 13645 16405 13679 16439
rect 14749 16405 14783 16439
rect 21465 16405 21499 16439
rect 25973 16405 26007 16439
rect 26709 16405 26743 16439
rect 2053 16201 2087 16235
rect 4169 16201 4203 16235
rect 6653 16201 6687 16235
rect 7113 16201 7147 16235
rect 8861 16201 8895 16235
rect 10425 16201 10459 16235
rect 11805 16201 11839 16235
rect 13737 16201 13771 16235
rect 17877 16201 17911 16235
rect 18797 16201 18831 16235
rect 19901 16201 19935 16235
rect 21465 16201 21499 16235
rect 22753 16201 22787 16235
rect 23121 16201 23155 16235
rect 23673 16201 23707 16235
rect 26525 16201 26559 16235
rect 3157 16133 3191 16167
rect 4537 16133 4571 16167
rect 13645 16133 13679 16167
rect 15301 16133 15335 16167
rect 24685 16133 24719 16167
rect 3709 16065 3743 16099
rect 7757 16065 7791 16099
rect 7941 16065 7975 16099
rect 8769 16065 8803 16099
rect 9413 16065 9447 16099
rect 10977 16065 11011 16099
rect 11437 16065 11471 16099
rect 13277 16065 13311 16099
rect 14289 16065 14323 16099
rect 15853 16065 15887 16099
rect 18337 16065 18371 16099
rect 20453 16065 20487 16099
rect 22017 16065 22051 16099
rect 24225 16065 24259 16099
rect 1409 15997 1443 16031
rect 3617 15997 3651 16031
rect 8309 15997 8343 16031
rect 9229 15997 9263 16031
rect 14105 15997 14139 16031
rect 18705 15997 18739 16031
rect 18981 15997 19015 16031
rect 20269 15997 20303 16031
rect 9321 15929 9355 15963
rect 9965 15929 9999 15963
rect 10793 15929 10827 15963
rect 12909 15929 12943 15963
rect 14197 15929 14231 15963
rect 20361 15929 20395 15963
rect 21925 15929 21959 15963
rect 23489 15929 23523 15963
rect 24041 15929 24075 15963
rect 1593 15861 1627 15895
rect 2329 15861 2363 15895
rect 3065 15861 3099 15895
rect 3525 15861 3559 15895
rect 4905 15861 4939 15895
rect 7297 15861 7331 15895
rect 7665 15861 7699 15895
rect 10333 15861 10367 15895
rect 10885 15861 10919 15895
rect 14749 15861 14783 15895
rect 15209 15861 15243 15895
rect 15669 15861 15703 15895
rect 15761 15861 15795 15895
rect 19441 15861 19475 15895
rect 19717 15861 19751 15895
rect 21281 15861 21315 15895
rect 21833 15861 21867 15895
rect 24133 15861 24167 15895
rect 4077 15657 4111 15691
rect 6193 15657 6227 15691
rect 8861 15657 8895 15691
rect 9689 15657 9723 15691
rect 10793 15657 10827 15691
rect 11069 15657 11103 15691
rect 13185 15657 13219 15691
rect 15577 15657 15611 15691
rect 19625 15657 19659 15691
rect 22937 15657 22971 15691
rect 24317 15657 24351 15691
rect 4445 15589 4479 15623
rect 6929 15589 6963 15623
rect 7757 15589 7791 15623
rect 16948 15589 16982 15623
rect 23949 15589 23983 15623
rect 1409 15521 1443 15555
rect 1676 15521 1710 15555
rect 10057 15521 10091 15555
rect 14013 15521 14047 15555
rect 16681 15521 16715 15555
rect 20729 15521 20763 15555
rect 23305 15521 23339 15555
rect 26893 15521 26927 15555
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 6285 15453 6319 15487
rect 6469 15453 6503 15487
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 23397 15453 23431 15487
rect 23489 15453 23523 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 2789 15385 2823 15419
rect 3433 15385 3467 15419
rect 5825 15317 5859 15351
rect 7389 15317 7423 15351
rect 13553 15317 13587 15351
rect 13645 15317 13679 15351
rect 18061 15317 18095 15351
rect 19073 15317 19107 15351
rect 19993 15317 20027 15351
rect 20545 15317 20579 15351
rect 21557 15317 21591 15351
rect 26065 15317 26099 15351
rect 26525 15317 26559 15351
rect 1777 15113 1811 15147
rect 2697 15113 2731 15147
rect 4169 15113 4203 15147
rect 4537 15113 4571 15147
rect 4813 15113 4847 15147
rect 5825 15113 5859 15147
rect 10425 15113 10459 15147
rect 13093 15113 13127 15147
rect 13553 15113 13587 15147
rect 15117 15113 15151 15147
rect 16773 15113 16807 15147
rect 19073 15113 19107 15147
rect 20729 15113 20763 15147
rect 22661 15113 22695 15147
rect 12725 15045 12759 15079
rect 17049 15045 17083 15079
rect 19625 15045 19659 15079
rect 3249 14977 3283 15011
rect 5549 14977 5583 15011
rect 6837 14977 6871 15011
rect 14013 14977 14047 15011
rect 14105 14977 14139 15011
rect 15669 14977 15703 15011
rect 20177 14977 20211 15011
rect 24317 14977 24351 15011
rect 25145 14977 25179 15011
rect 3065 14909 3099 14943
rect 14657 14909 14691 14943
rect 15485 14909 15519 14943
rect 19257 14909 19291 14943
rect 20085 14909 20119 14943
rect 23029 14909 23063 14943
rect 24869 14909 24903 14943
rect 25881 14909 25915 14943
rect 26065 14909 26099 14943
rect 2237 14841 2271 14875
rect 3157 14841 3191 14875
rect 6653 14841 6687 14875
rect 7104 14841 7138 14875
rect 13921 14841 13955 14875
rect 14933 14841 14967 14875
rect 15577 14841 15611 14875
rect 18981 14841 19015 14875
rect 19993 14841 20027 14875
rect 24041 14841 24075 14875
rect 24961 14841 24995 14875
rect 26332 14841 26366 14875
rect 2605 14773 2639 14807
rect 3709 14773 3743 14807
rect 6285 14773 6319 14807
rect 8217 14773 8251 14807
rect 9781 14773 9815 14807
rect 10149 14773 10183 14807
rect 13369 14773 13403 14807
rect 23305 14773 23339 14807
rect 24501 14773 24535 14807
rect 27445 14773 27479 14807
rect 2789 14569 2823 14603
rect 6009 14569 6043 14603
rect 7113 14569 7147 14603
rect 9229 14569 9263 14603
rect 13185 14569 13219 14603
rect 13645 14569 13679 14603
rect 26157 14569 26191 14603
rect 27169 14569 27203 14603
rect 5917 14501 5951 14535
rect 10784 14501 10818 14535
rect 14013 14501 14047 14535
rect 1409 14433 1443 14467
rect 1665 14433 1699 14467
rect 6929 14433 6963 14467
rect 7481 14433 7515 14467
rect 9413 14433 9447 14467
rect 9873 14433 9907 14467
rect 10517 14433 10551 14467
rect 13553 14433 13587 14467
rect 15485 14433 15519 14467
rect 16405 14433 16439 14467
rect 17969 14433 18003 14467
rect 18236 14433 18270 14467
rect 22836 14433 22870 14467
rect 6193 14365 6227 14399
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 16497 14365 16531 14399
rect 16589 14365 16623 14399
rect 22569 14365 22603 14399
rect 5549 14229 5583 14263
rect 8125 14229 8159 14263
rect 11897 14229 11931 14263
rect 16037 14229 16071 14263
rect 19349 14229 19383 14263
rect 19993 14229 20027 14263
rect 23949 14229 23983 14263
rect 24593 14229 24627 14263
rect 26801 14229 26835 14263
rect 1593 14025 1627 14059
rect 1961 14025 1995 14059
rect 4445 14025 4479 14059
rect 5273 14025 5307 14059
rect 6653 14025 6687 14059
rect 10517 14025 10551 14059
rect 11713 14025 11747 14059
rect 14473 14025 14507 14059
rect 15577 14025 15611 14059
rect 18613 14025 18647 14059
rect 21557 14025 21591 14059
rect 22661 14025 22695 14059
rect 5641 13957 5675 13991
rect 7481 13957 7515 13991
rect 9137 13957 9171 13991
rect 10701 13957 10735 13991
rect 16037 13957 16071 13991
rect 24593 13957 24627 13991
rect 25789 13957 25823 13991
rect 2973 13889 3007 13923
rect 7941 13889 7975 13923
rect 8125 13889 8159 13923
rect 9597 13889 9631 13923
rect 9781 13889 9815 13923
rect 11253 13889 11287 13923
rect 13737 13889 13771 13923
rect 15853 13889 15887 13923
rect 16589 13889 16623 13923
rect 20085 13889 20119 13923
rect 25237 13889 25271 13923
rect 26065 13889 26099 13923
rect 26893 13889 26927 13923
rect 3065 13821 3099 13855
rect 3332 13821 3366 13855
rect 6285 13821 6319 13855
rect 7205 13821 7239 13855
rect 9045 13821 9079 13855
rect 11161 13821 11195 13855
rect 14105 13821 14139 13855
rect 15209 13821 15243 13855
rect 16497 13821 16531 13855
rect 17141 13821 17175 13855
rect 20177 13821 20211 13855
rect 20444 13821 20478 13855
rect 24225 13821 24259 13855
rect 25145 13821 25179 13855
rect 26709 13821 26743 13855
rect 5733 13753 5767 13787
rect 7849 13753 7883 13787
rect 8677 13753 8711 13787
rect 9505 13753 9539 13787
rect 11069 13753 11103 13787
rect 25053 13753 25087 13787
rect 26617 13753 26651 13787
rect 10241 13685 10275 13719
rect 16405 13685 16439 13719
rect 18245 13685 18279 13719
rect 22937 13685 22971 13719
rect 24685 13685 24719 13719
rect 26249 13685 26283 13719
rect 5641 13481 5675 13515
rect 6285 13481 6319 13515
rect 7205 13481 7239 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 9229 13481 9263 13515
rect 10701 13481 10735 13515
rect 12541 13481 12575 13515
rect 16129 13481 16163 13515
rect 16773 13481 16807 13515
rect 17233 13481 17267 13515
rect 18337 13481 18371 13515
rect 20177 13481 20211 13515
rect 24685 13481 24719 13515
rect 26249 13481 26283 13515
rect 6193 13413 6227 13447
rect 7941 13413 7975 13447
rect 10149 13413 10183 13447
rect 16405 13413 16439 13447
rect 17141 13413 17175 13447
rect 22744 13413 22778 13447
rect 7573 13345 7607 13379
rect 10057 13345 10091 13379
rect 12725 13345 12759 13379
rect 12992 13345 13026 13379
rect 18705 13345 18739 13379
rect 26893 13345 26927 13379
rect 1685 13277 1719 13311
rect 3157 13277 3191 13311
rect 6377 13277 6411 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 10333 13277 10367 13311
rect 17325 13277 17359 13311
rect 18797 13277 18831 13311
rect 18889 13277 18923 13311
rect 22477 13277 22511 13311
rect 26985 13277 27019 13311
rect 27169 13277 27203 13311
rect 9689 13209 9723 13243
rect 25697 13209 25731 13243
rect 4721 13141 4755 13175
rect 5825 13141 5859 13175
rect 7389 13141 7423 13175
rect 11069 13141 11103 13175
rect 14105 13141 14139 13175
rect 14749 13141 14783 13175
rect 23857 13141 23891 13175
rect 26525 13141 26559 13175
rect 5825 12937 5859 12971
rect 6285 12937 6319 12971
rect 6561 12937 6595 12971
rect 7389 12937 7423 12971
rect 8217 12937 8251 12971
rect 9229 12937 9263 12971
rect 9781 12937 9815 12971
rect 13921 12937 13955 12971
rect 15853 12937 15887 12971
rect 17049 12937 17083 12971
rect 19073 12937 19107 12971
rect 22201 12937 22235 12971
rect 22569 12937 22603 12971
rect 27077 12937 27111 12971
rect 7757 12869 7791 12903
rect 15945 12869 15979 12903
rect 17325 12869 17359 12903
rect 25237 12869 25271 12903
rect 4169 12801 4203 12835
rect 5181 12801 5215 12835
rect 8125 12801 8159 12835
rect 9689 12801 9723 12835
rect 10241 12801 10275 12835
rect 10425 12801 10459 12835
rect 11897 12801 11931 12835
rect 13369 12801 13403 12835
rect 14933 12801 14967 12835
rect 15485 12801 15519 12835
rect 16405 12801 16439 12835
rect 16497 12801 16531 12835
rect 24225 12801 24259 12835
rect 24317 12801 24351 12835
rect 25513 12801 25547 12835
rect 26341 12801 26375 12835
rect 27261 12801 27295 12835
rect 1409 12733 1443 12767
rect 1961 12733 1995 12767
rect 4997 12733 5031 12767
rect 8401 12733 8435 12767
rect 12265 12733 12299 12767
rect 13093 12733 13127 12767
rect 13185 12733 13219 12767
rect 14749 12733 14783 12767
rect 14841 12733 14875 12767
rect 16313 12733 16347 12767
rect 18705 12733 18739 12767
rect 23121 12733 23155 12767
rect 24133 12733 24167 12767
rect 26065 12733 26099 12767
rect 26709 12733 26743 12767
rect 4537 12665 4571 12699
rect 5089 12665 5123 12699
rect 10149 12665 10183 12699
rect 23489 12665 23523 12699
rect 1593 12597 1627 12631
rect 4629 12597 4663 12631
rect 8861 12597 8895 12631
rect 10885 12597 10919 12631
rect 12725 12597 12759 12631
rect 14197 12597 14231 12631
rect 14381 12597 14415 12631
rect 18337 12597 18371 12631
rect 23765 12597 23799 12631
rect 25697 12597 25731 12631
rect 26157 12597 26191 12631
rect 1869 12393 1903 12427
rect 6193 12393 6227 12427
rect 7389 12393 7423 12427
rect 8125 12393 8159 12427
rect 12817 12393 12851 12427
rect 13185 12393 13219 12427
rect 16865 12393 16899 12427
rect 23857 12393 23891 12427
rect 24869 12393 24903 12427
rect 25329 12393 25363 12427
rect 27169 12393 27203 12427
rect 16037 12325 16071 12359
rect 21180 12325 21214 12359
rect 25237 12325 25271 12359
rect 4997 12257 5031 12291
rect 13369 12257 13403 12291
rect 17509 12257 17543 12291
rect 20913 12257 20947 12291
rect 26525 12257 26559 12291
rect 5089 12189 5123 12223
rect 5273 12189 5307 12223
rect 17601 12189 17635 12223
rect 17785 12189 17819 12223
rect 25421 12189 25455 12223
rect 4629 12053 4663 12087
rect 8493 12053 8527 12087
rect 9873 12053 9907 12087
rect 10333 12053 10367 12087
rect 14657 12053 14691 12087
rect 17141 12053 17175 12087
rect 19257 12053 19291 12087
rect 22293 12053 22327 12087
rect 26709 12053 26743 12087
rect 4721 11849 4755 11883
rect 5733 11849 5767 11883
rect 11161 11849 11195 11883
rect 17509 11849 17543 11883
rect 21281 11849 21315 11883
rect 24961 11849 24995 11883
rect 25329 11849 25363 11883
rect 25605 11849 25639 11883
rect 27353 11849 27387 11883
rect 12541 11781 12575 11815
rect 14749 11781 14783 11815
rect 1869 11713 1903 11747
rect 5273 11713 5307 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 13829 11713 13863 11747
rect 13921 11713 13955 11747
rect 14381 11713 14415 11747
rect 18061 11713 18095 11747
rect 19257 11713 19291 11747
rect 4629 11645 4663 11679
rect 5089 11645 5123 11679
rect 7297 11645 7331 11679
rect 9321 11645 9355 11679
rect 9781 11645 9815 11679
rect 26433 11645 26467 11679
rect 26985 11645 27019 11679
rect 1777 11577 1811 11611
rect 2136 11577 2170 11611
rect 3893 11577 3927 11611
rect 7205 11577 7239 11611
rect 7542 11577 7576 11611
rect 10026 11577 10060 11611
rect 11897 11577 11931 11611
rect 12909 11577 12943 11611
rect 13737 11577 13771 11611
rect 15209 11577 15243 11611
rect 16865 11577 16899 11611
rect 19165 11577 19199 11611
rect 19502 11577 19536 11611
rect 3249 11509 3283 11543
rect 4261 11509 4295 11543
rect 5181 11509 5215 11543
rect 8677 11509 8711 11543
rect 9597 11509 9631 11543
rect 12173 11509 12207 11543
rect 13369 11509 13403 11543
rect 17141 11509 17175 11543
rect 20637 11509 20671 11543
rect 21649 11509 21683 11543
rect 26617 11509 26651 11543
rect 5181 11305 5215 11339
rect 5457 11305 5491 11339
rect 7665 11305 7699 11339
rect 12541 11305 12575 11339
rect 13093 11305 13127 11339
rect 14013 11305 14047 11339
rect 14105 11305 14139 11339
rect 17325 11305 17359 11339
rect 18429 11305 18463 11339
rect 18797 11305 18831 11339
rect 26709 11305 26743 11339
rect 17233 11237 17267 11271
rect 1409 11169 1443 11203
rect 4445 11169 4479 11203
rect 22017 11169 22051 11203
rect 22284 11169 22318 11203
rect 26525 11169 26559 11203
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 7757 11101 7791 11135
rect 7849 11101 7883 11135
rect 14289 11101 14323 11135
rect 17417 11101 17451 11135
rect 18889 11101 18923 11135
rect 19073 11101 19107 11135
rect 1593 11033 1627 11067
rect 4077 11033 4111 11067
rect 7297 11033 7331 11067
rect 13369 11033 13403 11067
rect 13645 11033 13679 11067
rect 16865 11033 16899 11067
rect 21925 11033 21959 11067
rect 23397 10965 23431 10999
rect 1593 10761 1627 10795
rect 2053 10761 2087 10795
rect 2421 10761 2455 10795
rect 3617 10761 3651 10795
rect 7389 10761 7423 10795
rect 14381 10761 14415 10795
rect 17325 10761 17359 10795
rect 17785 10761 17819 10795
rect 18521 10761 18555 10795
rect 21649 10761 21683 10795
rect 22845 10761 22879 10795
rect 26525 10761 26559 10795
rect 3249 10693 3283 10727
rect 4445 10693 4479 10727
rect 7757 10693 7791 10727
rect 16589 10693 16623 10727
rect 18889 10693 18923 10727
rect 3985 10625 4019 10659
rect 5089 10625 5123 10659
rect 8033 10625 8067 10659
rect 12909 10625 12943 10659
rect 22477 10625 22511 10659
rect 1409 10557 1443 10591
rect 13001 10557 13035 10591
rect 13268 10557 13302 10591
rect 19073 10557 19107 10591
rect 19349 10557 19383 10591
rect 24225 10557 24259 10591
rect 24470 10489 24504 10523
rect 4353 10421 4387 10455
rect 4813 10421 4847 10455
rect 4905 10421 4939 10455
rect 16957 10421 16991 10455
rect 21833 10421 21867 10455
rect 22201 10421 22235 10455
rect 22293 10421 22327 10455
rect 24041 10421 24075 10455
rect 25605 10421 25639 10455
rect 26709 10421 26743 10455
rect 4905 10217 4939 10251
rect 5089 10217 5123 10251
rect 5457 10217 5491 10251
rect 14105 10217 14139 10251
rect 19257 10217 19291 10251
rect 21557 10217 21591 10251
rect 21925 10217 21959 10251
rect 22385 10217 22419 10251
rect 24225 10217 24259 10251
rect 24869 10217 24903 10251
rect 25329 10217 25363 10251
rect 26525 10217 26559 10251
rect 26985 10217 27019 10251
rect 5549 10149 5583 10183
rect 13737 10149 13771 10183
rect 19165 10149 19199 10183
rect 1676 10081 1710 10115
rect 4537 10081 4571 10115
rect 10241 10081 10275 10115
rect 10508 10081 10542 10115
rect 14381 10081 14415 10115
rect 15844 10081 15878 10115
rect 20637 10081 20671 10115
rect 22753 10081 22787 10115
rect 25237 10081 25271 10115
rect 26893 10081 26927 10115
rect 1409 10013 1443 10047
rect 5641 10013 5675 10047
rect 15577 10013 15611 10047
rect 19349 10013 19383 10047
rect 22845 10013 22879 10047
rect 22937 10013 22971 10047
rect 25421 10013 25455 10047
rect 27077 10013 27111 10047
rect 18153 9945 18187 9979
rect 22293 9945 22327 9979
rect 2789 9877 2823 9911
rect 3525 9877 3559 9911
rect 7849 9877 7883 9911
rect 11621 9877 11655 9911
rect 12449 9877 12483 9911
rect 13093 9877 13127 9911
rect 16957 9877 16991 9911
rect 17785 9877 17819 9911
rect 18429 9877 18463 9911
rect 18797 9877 18831 9911
rect 19901 9877 19935 9911
rect 20453 9877 20487 9911
rect 23673 9877 23707 9911
rect 25881 9877 25915 9911
rect 2329 9673 2363 9707
rect 3433 9673 3467 9707
rect 10241 9673 10275 9707
rect 10333 9673 10367 9707
rect 13921 9673 13955 9707
rect 16037 9673 16071 9707
rect 17601 9673 17635 9707
rect 19073 9673 19107 9707
rect 22569 9673 22603 9707
rect 24869 9673 24903 9707
rect 25329 9673 25363 9707
rect 26893 9673 26927 9707
rect 27261 9673 27295 9707
rect 4997 9605 5031 9639
rect 9229 9605 9263 9639
rect 12173 9605 12207 9639
rect 20913 9605 20947 9639
rect 23673 9605 23707 9639
rect 25789 9605 25823 9639
rect 3341 9537 3375 9571
rect 4077 9537 4111 9571
rect 5641 9537 5675 9571
rect 7849 9537 7883 9571
rect 10885 9537 10919 9571
rect 13001 9537 13035 9571
rect 17233 9537 17267 9571
rect 18521 9537 18555 9571
rect 18613 9537 18647 9571
rect 20545 9537 20579 9571
rect 22017 9537 22051 9571
rect 24225 9537 24259 9571
rect 26433 9537 26467 9571
rect 1409 9469 1443 9503
rect 3801 9469 3835 9503
rect 6101 9469 6135 9503
rect 10517 9469 10551 9503
rect 11161 9469 11195 9503
rect 14013 9469 14047 9503
rect 14269 9469 14303 9503
rect 17877 9469 17911 9503
rect 18429 9469 18463 9503
rect 20269 9469 20303 9503
rect 21925 9469 21959 9503
rect 26249 9469 26283 9503
rect 27445 9469 27479 9503
rect 27997 9469 28031 9503
rect 2053 9401 2087 9435
rect 4537 9401 4571 9435
rect 5365 9401 5399 9435
rect 8116 9401 8150 9435
rect 12909 9401 12943 9435
rect 20361 9401 20395 9435
rect 21833 9401 21867 9435
rect 23121 9401 23155 9435
rect 24133 9401 24167 9435
rect 26341 9401 26375 9435
rect 1593 9333 1627 9367
rect 3893 9333 3927 9367
rect 4905 9333 4939 9367
rect 5457 9333 5491 9367
rect 7757 9333 7791 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 15393 9333 15427 9367
rect 16405 9333 16439 9367
rect 17693 9333 17727 9367
rect 18061 9333 18095 9367
rect 19717 9333 19751 9367
rect 19901 9333 19935 9367
rect 21281 9333 21315 9367
rect 21465 9333 21499 9367
rect 23489 9333 23523 9367
rect 24041 9333 24075 9367
rect 25881 9333 25915 9367
rect 27629 9333 27663 9367
rect 2053 9129 2087 9163
rect 2697 9129 2731 9163
rect 3525 9129 3559 9163
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 5089 9129 5123 9163
rect 5549 9129 5583 9163
rect 5917 9129 5951 9163
rect 6929 9129 6963 9163
rect 10885 9129 10919 9163
rect 12541 9129 12575 9163
rect 16497 9129 16531 9163
rect 17877 9129 17911 9163
rect 19257 9129 19291 9163
rect 19717 9129 19751 9163
rect 20361 9129 20395 9163
rect 21557 9129 21591 9163
rect 22477 9129 22511 9163
rect 23029 9129 23063 9163
rect 24961 9129 24995 9163
rect 25973 9129 26007 9163
rect 26709 9129 26743 9163
rect 18797 9061 18831 9095
rect 19625 9061 19659 9095
rect 22753 9061 22787 9095
rect 23489 9061 23523 9095
rect 27077 9061 27111 9095
rect 1409 8993 1443 9027
rect 2513 8993 2547 9027
rect 4445 8993 4479 9027
rect 7288 8993 7322 9027
rect 10609 8993 10643 9027
rect 11805 8993 11839 9027
rect 17785 8993 17819 9027
rect 18521 8993 18555 9027
rect 23397 8993 23431 9027
rect 26525 8993 26559 9027
rect 4721 8925 4755 8959
rect 7021 8925 7055 8959
rect 11897 8925 11931 8959
rect 12081 8925 12115 8959
rect 17969 8925 18003 8959
rect 19809 8925 19843 8959
rect 23581 8925 23615 8959
rect 1593 8789 1627 8823
rect 8401 8789 8435 8823
rect 9045 8789 9079 8823
rect 10425 8789 10459 8823
rect 11437 8789 11471 8823
rect 14013 8789 14047 8823
rect 17417 8789 17451 8823
rect 24133 8789 24167 8823
rect 2053 8585 2087 8619
rect 2421 8585 2455 8619
rect 6653 8585 6687 8619
rect 8861 8585 8895 8619
rect 11805 8585 11839 8619
rect 17877 8585 17911 8619
rect 18245 8585 18279 8619
rect 19257 8585 19291 8619
rect 19717 8585 19751 8619
rect 20085 8585 20119 8619
rect 23673 8585 23707 8619
rect 27537 8585 27571 8619
rect 1593 8517 1627 8551
rect 3433 8517 3467 8551
rect 4169 8517 4203 8551
rect 7389 8517 7423 8551
rect 10609 8517 10643 8551
rect 16405 8517 16439 8551
rect 22753 8517 22787 8551
rect 26985 8517 27019 8551
rect 2789 8449 2823 8483
rect 3801 8449 3835 8483
rect 4997 8449 5031 8483
rect 5089 8449 5123 8483
rect 5917 8449 5951 8483
rect 7297 8449 7331 8483
rect 7941 8449 7975 8483
rect 8493 8449 8527 8483
rect 9597 8449 9631 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 12449 8449 12483 8483
rect 16957 8449 16991 8483
rect 23121 8449 23155 8483
rect 24317 8449 24351 8483
rect 1409 8381 1443 8415
rect 9321 8381 9355 8415
rect 9413 8381 9447 8415
rect 10241 8381 10275 8415
rect 11069 8381 11103 8415
rect 16773 8381 16807 8415
rect 23489 8381 23523 8415
rect 25605 8381 25639 8415
rect 4905 8313 4939 8347
rect 5549 8313 5583 8347
rect 7757 8313 7791 8347
rect 12081 8313 12115 8347
rect 16221 8313 16255 8347
rect 22385 8313 22419 8347
rect 24041 8313 24075 8347
rect 24133 8313 24167 8347
rect 25421 8313 25455 8347
rect 25850 8313 25884 8347
rect 4537 8245 4571 8279
rect 7849 8245 7883 8279
rect 8953 8245 8987 8279
rect 10701 8245 10735 8279
rect 16865 8245 16899 8279
rect 17417 8245 17451 8279
rect 2237 8041 2271 8075
rect 2697 8041 2731 8075
rect 4997 8041 5031 8075
rect 6101 8041 6135 8075
rect 7113 8041 7147 8075
rect 7757 8041 7791 8075
rect 8033 8041 8067 8075
rect 8493 8041 8527 8075
rect 9689 8041 9723 8075
rect 10057 8041 10091 8075
rect 10793 8041 10827 8075
rect 11529 8041 11563 8075
rect 13461 8041 13495 8075
rect 14841 8041 14875 8075
rect 16497 8041 16531 8075
rect 18061 8041 18095 8075
rect 21373 8041 21407 8075
rect 23121 8041 23155 8075
rect 23581 8041 23615 8075
rect 25605 8041 25639 8075
rect 26709 8041 26743 8075
rect 4905 7973 4939 8007
rect 8401 7973 8435 8007
rect 1409 7905 1443 7939
rect 2513 7905 2547 7939
rect 7389 7905 7423 7939
rect 10149 7905 10183 7939
rect 12081 7905 12115 7939
rect 12348 7905 12382 7939
rect 16681 7905 16715 7939
rect 16937 7905 16971 7939
rect 21281 7905 21315 7939
rect 23949 7905 23983 7939
rect 26525 7905 26559 7939
rect 5089 7837 5123 7871
rect 8677 7837 8711 7871
rect 10333 7837 10367 7871
rect 19809 7837 19843 7871
rect 21465 7837 21499 7871
rect 24041 7837 24075 7871
rect 24225 7837 24259 7871
rect 4353 7769 4387 7803
rect 7205 7769 7239 7803
rect 20913 7769 20947 7803
rect 1593 7701 1627 7735
rect 4537 7701 4571 7735
rect 5549 7701 5583 7735
rect 19165 7701 19199 7735
rect 20637 7701 20671 7735
rect 2145 7497 2179 7531
rect 4261 7497 4295 7531
rect 7297 7497 7331 7531
rect 8125 7497 8159 7531
rect 8493 7497 8527 7531
rect 8861 7497 8895 7531
rect 9413 7497 9447 7531
rect 9781 7497 9815 7531
rect 10517 7497 10551 7531
rect 12633 7497 12667 7531
rect 16773 7497 16807 7531
rect 20085 7497 20119 7531
rect 22569 7497 22603 7531
rect 23121 7497 23155 7531
rect 23673 7497 23707 7531
rect 26617 7497 26651 7531
rect 4629 7429 4663 7463
rect 17049 7429 17083 7463
rect 27353 7429 27387 7463
rect 27721 7429 27755 7463
rect 2237 7361 2271 7395
rect 5181 7361 5215 7395
rect 5273 7361 5307 7395
rect 5733 7361 5767 7395
rect 10149 7361 10183 7395
rect 11161 7361 11195 7395
rect 12081 7361 12115 7395
rect 14749 7361 14783 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 24317 7361 24351 7395
rect 1685 7293 1719 7327
rect 5089 7293 5123 7327
rect 6101 7293 6135 7327
rect 11069 7293 11103 7327
rect 18981 7293 19015 7327
rect 20637 7293 20671 7327
rect 24041 7293 24075 7327
rect 26433 7293 26467 7327
rect 26985 7293 27019 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 2504 7225 2538 7259
rect 10977 7225 11011 7259
rect 14657 7225 14691 7259
rect 15016 7225 15050 7259
rect 19441 7225 19475 7259
rect 20904 7225 20938 7259
rect 23489 7225 23523 7259
rect 3617 7157 3651 7191
rect 4721 7157 4755 7191
rect 10609 7157 10643 7191
rect 16129 7157 16163 7191
rect 19073 7157 19107 7191
rect 20453 7157 20487 7191
rect 22017 7157 22051 7191
rect 24133 7157 24167 7191
rect 24685 7157 24719 7191
rect 2329 6953 2363 6987
rect 9965 6953 9999 6987
rect 15669 6953 15703 6987
rect 21281 6953 21315 6987
rect 24041 6953 24075 6987
rect 1409 6817 1443 6851
rect 4905 6817 4939 6851
rect 5172 6817 5206 6851
rect 10609 6817 10643 6851
rect 14013 6817 14047 6851
rect 16405 6817 16439 6851
rect 17325 6817 17359 6851
rect 19165 6817 19199 6851
rect 20729 6817 20763 6851
rect 26525 6817 26559 6851
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 14749 6749 14783 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 17417 6749 17451 6783
rect 17509 6749 17543 6783
rect 21373 6749 21407 6783
rect 21465 6749 21499 6783
rect 13645 6681 13679 6715
rect 20913 6681 20947 6715
rect 26709 6681 26743 6715
rect 1593 6613 1627 6647
rect 2697 6613 2731 6647
rect 4629 6613 4663 6647
rect 6285 6613 6319 6647
rect 8861 6613 8895 6647
rect 15301 6613 15335 6647
rect 16957 6613 16991 6647
rect 23765 6613 23799 6647
rect 24501 6613 24535 6647
rect 1685 6409 1719 6443
rect 5549 6409 5583 6443
rect 10149 6409 10183 6443
rect 13369 6409 13403 6443
rect 15669 6409 15703 6443
rect 17785 6409 17819 6443
rect 21005 6409 21039 6443
rect 21281 6409 21315 6443
rect 25329 6409 25363 6443
rect 27077 6409 27111 6443
rect 27353 6409 27387 6443
rect 5089 6341 5123 6375
rect 10333 6341 10367 6375
rect 17417 6341 17451 6375
rect 26617 6341 26651 6375
rect 2329 6273 2363 6307
rect 2973 6273 3007 6307
rect 3985 6273 4019 6307
rect 4629 6273 4663 6307
rect 9321 6273 9355 6307
rect 9781 6273 9815 6307
rect 10885 6273 10919 6307
rect 14565 6273 14599 6307
rect 15301 6273 15335 6307
rect 16957 6273 16991 6307
rect 18061 6273 18095 6307
rect 2789 6205 2823 6239
rect 3433 6205 3467 6239
rect 4445 6205 4479 6239
rect 8677 6205 8711 6239
rect 9137 6205 9171 6239
rect 10701 6205 10735 6239
rect 15025 6205 15059 6239
rect 16865 6205 16899 6239
rect 23121 6205 23155 6239
rect 23949 6205 23983 6239
rect 26433 6205 26467 6239
rect 9229 6137 9263 6171
rect 10793 6137 10827 6171
rect 15117 6137 15151 6171
rect 16313 6137 16347 6171
rect 16773 6137 16807 6171
rect 24194 6137 24228 6171
rect 2421 6069 2455 6103
rect 2881 6069 2915 6103
rect 4077 6069 4111 6103
rect 4537 6069 4571 6103
rect 7757 6069 7791 6103
rect 8769 6069 8803 6103
rect 13645 6069 13679 6103
rect 14013 6069 14047 6103
rect 14657 6069 14691 6103
rect 16405 6069 16439 6103
rect 21649 6069 21683 6103
rect 23489 6069 23523 6103
rect 2237 5865 2271 5899
rect 3341 5865 3375 5899
rect 4261 5865 4295 5899
rect 4721 5865 4755 5899
rect 10333 5865 10367 5899
rect 12817 5865 12851 5899
rect 15853 5865 15887 5899
rect 16497 5865 16531 5899
rect 17049 5865 17083 5899
rect 17693 5865 17727 5899
rect 19717 5865 19751 5899
rect 20913 5865 20947 5899
rect 23857 5865 23891 5899
rect 2605 5797 2639 5831
rect 6276 5797 6310 5831
rect 17141 5797 17175 5831
rect 19625 5797 19659 5831
rect 22722 5797 22756 5831
rect 6009 5729 6043 5763
rect 11437 5729 11471 5763
rect 11693 5729 11727 5763
rect 21281 5729 21315 5763
rect 22477 5729 22511 5763
rect 26525 5729 26559 5763
rect 2145 5661 2179 5695
rect 2697 5661 2731 5695
rect 2789 5661 2823 5695
rect 17233 5661 17267 5695
rect 19901 5661 19935 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 8861 5593 8895 5627
rect 26709 5593 26743 5627
rect 7389 5525 7423 5559
rect 14657 5525 14691 5559
rect 15485 5525 15519 5559
rect 16681 5525 16715 5559
rect 19257 5525 19291 5559
rect 20729 5525 20763 5559
rect 1593 5321 1627 5355
rect 2513 5321 2547 5355
rect 4721 5321 4755 5355
rect 6101 5321 6135 5355
rect 11897 5321 11931 5355
rect 15577 5321 15611 5355
rect 16773 5321 16807 5355
rect 17417 5321 17451 5355
rect 18981 5321 19015 5355
rect 19717 5321 19751 5355
rect 20453 5321 20487 5355
rect 20637 5321 20671 5355
rect 21649 5321 21683 5355
rect 22109 5321 22143 5355
rect 22937 5321 22971 5355
rect 27353 5321 27387 5355
rect 2329 5253 2363 5287
rect 6377 5253 6411 5287
rect 8493 5253 8527 5287
rect 17141 5253 17175 5287
rect 19349 5253 19383 5287
rect 22477 5253 22511 5287
rect 3157 5185 3191 5219
rect 3893 5185 3927 5219
rect 8125 5185 8159 5219
rect 9045 5185 9079 5219
rect 9229 5185 9263 5219
rect 21281 5185 21315 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 4077 5117 4111 5151
rect 7757 5117 7791 5151
rect 8953 5117 8987 5151
rect 14197 5117 14231 5151
rect 21097 5117 21131 5151
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 14105 5049 14139 5083
rect 14442 5049 14476 5083
rect 20177 5049 20211 5083
rect 2973 4981 3007 5015
rect 3617 4981 3651 5015
rect 4261 4981 4295 5015
rect 8585 4981 8619 5015
rect 11437 4981 11471 5015
rect 21005 4981 21039 5015
rect 26617 4981 26651 5015
rect 1593 4777 1627 4811
rect 2421 4777 2455 4811
rect 2881 4777 2915 4811
rect 3433 4777 3467 4811
rect 4721 4777 4755 4811
rect 7021 4777 7055 4811
rect 7573 4777 7607 4811
rect 8401 4777 8435 4811
rect 10517 4777 10551 4811
rect 12817 4777 12851 4811
rect 14657 4777 14691 4811
rect 20729 4777 20763 4811
rect 20913 4777 20947 4811
rect 11682 4709 11716 4743
rect 16764 4709 16798 4743
rect 21281 4709 21315 4743
rect 2329 4641 2363 4675
rect 2789 4641 2823 4675
rect 4077 4641 4111 4675
rect 11437 4641 11471 4675
rect 14197 4641 14231 4675
rect 16497 4641 16531 4675
rect 26525 4641 26559 4675
rect 3065 4573 3099 4607
rect 7941 4573 7975 4607
rect 8493 4573 8527 4607
rect 8585 4573 8619 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 4261 4437 4295 4471
rect 8033 4437 8067 4471
rect 17877 4437 17911 4471
rect 26709 4437 26743 4471
rect 2697 4233 2731 4267
rect 3709 4233 3743 4267
rect 5641 4233 5675 4267
rect 8953 4233 8987 4267
rect 11897 4233 11931 4267
rect 20913 4233 20947 4267
rect 27353 4233 27387 4267
rect 14473 4165 14507 4199
rect 2605 4097 2639 4131
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 6561 4097 6595 4131
rect 7481 4097 7515 4131
rect 8125 4097 8159 4131
rect 8861 4097 8895 4131
rect 9597 4097 9631 4131
rect 10425 4097 10459 4131
rect 11069 4097 11103 4131
rect 15117 4097 15151 4131
rect 16313 4097 16347 4131
rect 16957 4097 16991 4131
rect 20177 4097 20211 4131
rect 1409 4029 1443 4063
rect 4261 4029 4295 4063
rect 4517 4029 4551 4063
rect 7297 4029 7331 4063
rect 8493 4029 8527 4063
rect 9413 4029 9447 4063
rect 10885 4029 10919 4063
rect 14933 4029 14967 4063
rect 15025 4029 15059 4063
rect 16773 4029 16807 4063
rect 21005 4029 21039 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 4169 3961 4203 3995
rect 7389 3961 7423 3995
rect 9321 3961 9355 3995
rect 10977 3961 11011 3995
rect 15853 3961 15887 3995
rect 16865 3961 16899 3995
rect 20545 3961 20579 3995
rect 21272 3961 21306 3995
rect 1593 3893 1627 3927
rect 2237 3893 2271 3927
rect 3065 3893 3099 3927
rect 6929 3893 6963 3927
rect 10517 3893 10551 3927
rect 11621 3893 11655 3927
rect 14565 3893 14599 3927
rect 16405 3893 16439 3927
rect 17417 3893 17451 3927
rect 22385 3893 22419 3927
rect 26617 3893 26651 3927
rect 1593 3689 1627 3723
rect 2881 3689 2915 3723
rect 3433 3689 3467 3723
rect 4629 3689 4663 3723
rect 7021 3689 7055 3723
rect 9137 3689 9171 3723
rect 10517 3689 10551 3723
rect 12449 3689 12483 3723
rect 14657 3689 14691 3723
rect 16865 3689 16899 3723
rect 20361 3689 20395 3723
rect 20729 3689 20763 3723
rect 20913 3689 20947 3723
rect 21373 3689 21407 3723
rect 7380 3621 7414 3655
rect 16589 3621 16623 3655
rect 18398 3621 18432 3655
rect 21281 3621 21315 3655
rect 2789 3553 2823 3587
rect 4077 3553 4111 3587
rect 5181 3553 5215 3587
rect 7113 3553 7147 3587
rect 11069 3553 11103 3587
rect 11336 3553 11370 3587
rect 18153 3553 18187 3587
rect 25329 3553 25363 3587
rect 26525 3553 26559 3587
rect 2329 3485 2363 3519
rect 3065 3485 3099 3519
rect 21465 3485 21499 3519
rect 5365 3417 5399 3451
rect 8493 3417 8527 3451
rect 19533 3417 19567 3451
rect 25513 3417 25547 3451
rect 2421 3349 2455 3383
rect 3801 3349 3835 3383
rect 4261 3349 4295 3383
rect 26709 3349 26743 3383
rect 1961 3145 1995 3179
rect 3801 3145 3835 3179
rect 4813 3145 4847 3179
rect 5457 3145 5491 3179
rect 7665 3145 7699 3179
rect 8769 3145 8803 3179
rect 10149 3145 10183 3179
rect 11161 3145 11195 3179
rect 11529 3145 11563 3179
rect 18245 3145 18279 3179
rect 20361 3145 20395 3179
rect 21281 3145 21315 3179
rect 21649 3145 21683 3179
rect 24409 3145 24443 3179
rect 25329 3145 25363 3179
rect 27353 3145 27387 3179
rect 8217 3077 8251 3111
rect 18613 3077 18647 3111
rect 27077 3077 27111 3111
rect 4353 3009 4387 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 2421 2941 2455 2975
rect 4905 2941 4939 2975
rect 6653 2941 6687 2975
rect 6929 2941 6963 2975
rect 8677 2941 8711 2975
rect 9137 2941 9171 2975
rect 10333 2941 10367 2975
rect 13645 2941 13679 2975
rect 14381 2941 14415 2975
rect 20453 2941 20487 2975
rect 23673 2941 23707 2975
rect 26433 2941 26467 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 2666 2873 2700 2907
rect 7205 2873 7239 2907
rect 10609 2873 10643 2907
rect 13921 2873 13955 2907
rect 20729 2873 20763 2907
rect 23949 2873 23983 2907
rect 2237 2805 2271 2839
rect 5089 2805 5123 2839
rect 26617 2805 26651 2839
rect 27721 2805 27755 2839
rect 2697 2601 2731 2635
rect 3065 2601 3099 2635
rect 6377 2601 6411 2635
rect 7113 2601 7147 2635
rect 8861 2601 8895 2635
rect 19257 2601 19291 2635
rect 20637 2601 20671 2635
rect 21005 2601 21039 2635
rect 2053 2533 2087 2567
rect 3433 2533 3467 2567
rect 1409 2465 1443 2499
rect 2421 2465 2455 2499
rect 2513 2465 2547 2499
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 5549 2465 5583 2499
rect 7573 2465 7607 2499
rect 8309 2465 8343 2499
rect 9781 2465 9815 2499
rect 10517 2465 10551 2499
rect 11161 2465 11195 2499
rect 11897 2465 11931 2499
rect 14105 2465 14139 2499
rect 14841 2465 14875 2499
rect 16405 2465 16439 2499
rect 17141 2465 17175 2499
rect 18521 2465 18555 2499
rect 19809 2465 19843 2499
rect 22293 2465 22327 2499
rect 23029 2465 23063 2499
rect 24317 2465 24351 2499
rect 25053 2465 25087 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 4353 2397 4387 2431
rect 5825 2397 5859 2431
rect 7849 2397 7883 2431
rect 10057 2397 10091 2431
rect 11437 2397 11471 2431
rect 14381 2397 14415 2431
rect 16681 2397 16715 2431
rect 18797 2397 18831 2431
rect 20085 2397 20119 2431
rect 22569 2397 22603 2431
rect 24593 2397 24627 2431
rect 1593 2261 1627 2295
rect 25881 2261 25915 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3418 22108 3424 22160
rect 3476 22148 3482 22160
rect 10410 22148 10416 22160
rect 3476 22120 10416 22148
rect 3476 22108 3482 22120
rect 10410 22108 10416 22120
rect 10468 22108 10474 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 22537 20995 22595 21001
rect 22537 20992 22549 20995
rect 22428 20964 22549 20992
rect 22428 20952 22434 20964
rect 22537 20961 22549 20964
rect 22583 20961 22595 20995
rect 22537 20955 22595 20961
rect 22278 20924 22284 20936
rect 22239 20896 22284 20924
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 18046 20788 18052 20800
rect 2924 20760 18052 20788
rect 2924 20748 2930 20760
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 23566 20748 23572 20800
rect 23624 20788 23630 20800
rect 23661 20791 23719 20797
rect 23661 20788 23673 20791
rect 23624 20760 23673 20788
rect 23624 20748 23630 20760
rect 23661 20757 23673 20760
rect 23707 20757 23719 20791
rect 23661 20751 23719 20757
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21729 20587 21787 20593
rect 21729 20584 21741 20587
rect 21600 20556 21741 20584
rect 21600 20544 21606 20556
rect 21729 20553 21741 20556
rect 21775 20584 21787 20587
rect 22370 20584 22376 20596
rect 21775 20556 22376 20584
rect 21775 20553 21787 20556
rect 21729 20547 21787 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 13630 20380 13636 20392
rect 13591 20352 13636 20380
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 20349 20383 20407 20389
rect 20349 20349 20361 20383
rect 20395 20380 20407 20383
rect 20438 20380 20444 20392
rect 20395 20352 20444 20380
rect 20395 20349 20407 20352
rect 20349 20343 20407 20349
rect 20438 20340 20444 20352
rect 20496 20380 20502 20392
rect 22278 20380 22284 20392
rect 20496 20352 22284 20380
rect 20496 20340 20502 20352
rect 13541 20315 13599 20321
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 13878 20315 13936 20321
rect 13878 20312 13890 20315
rect 13587 20284 13890 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 13878 20281 13890 20284
rect 13924 20312 13936 20315
rect 14090 20312 14096 20324
rect 13924 20284 14096 20312
rect 13924 20281 13936 20284
rect 13878 20275 13936 20281
rect 14090 20272 14096 20284
rect 14148 20272 14154 20324
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 20257 20315 20315 20321
rect 20257 20312 20269 20315
rect 19760 20284 20269 20312
rect 19760 20272 19766 20284
rect 20257 20281 20269 20284
rect 20303 20312 20315 20315
rect 20594 20315 20652 20321
rect 20594 20312 20606 20315
rect 20303 20284 20606 20312
rect 20303 20281 20315 20284
rect 20257 20275 20315 20281
rect 20594 20281 20606 20284
rect 20640 20281 20652 20315
rect 22112 20312 22140 20352
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 26053 20383 26111 20389
rect 26053 20349 26065 20383
rect 26099 20380 26111 20383
rect 26099 20352 26740 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 22741 20315 22799 20321
rect 22741 20312 22753 20315
rect 22112 20284 22753 20312
rect 20594 20275 20652 20281
rect 22741 20281 22753 20284
rect 22787 20312 22799 20315
rect 23474 20312 23480 20324
rect 22787 20284 23480 20312
rect 22787 20281 22799 20284
rect 22741 20275 22799 20281
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15013 20247 15071 20253
rect 15013 20244 15025 20247
rect 14884 20216 15025 20244
rect 14884 20204 14890 20216
rect 15013 20213 15025 20216
rect 15059 20213 15071 20247
rect 26234 20244 26240 20256
rect 26195 20216 26240 20244
rect 15013 20207 15071 20213
rect 26234 20204 26240 20216
rect 26292 20204 26298 20256
rect 26712 20253 26740 20352
rect 26697 20247 26755 20253
rect 26697 20213 26709 20247
rect 26743 20244 26755 20247
rect 27522 20244 27528 20256
rect 26743 20216 27528 20244
rect 26743 20213 26755 20216
rect 26697 20207 26755 20213
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 13630 20040 13636 20052
rect 13591 20012 13636 20040
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 19702 20040 19708 20052
rect 19663 20012 19708 20040
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 20438 20040 20444 20052
rect 20399 20012 20444 20040
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21545 20043 21603 20049
rect 21545 20009 21557 20043
rect 21591 20040 21603 20043
rect 22462 20040 22468 20052
rect 21591 20012 22468 20040
rect 21591 20009 21603 20012
rect 21545 20003 21603 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 18322 19932 18328 19984
rect 18380 19972 18386 19984
rect 18570 19975 18628 19981
rect 18570 19972 18582 19975
rect 18380 19944 18582 19972
rect 18380 19932 18386 19944
rect 18570 19941 18582 19944
rect 18616 19941 18628 19975
rect 18570 19935 18628 19941
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 23733 19907 23791 19913
rect 23733 19904 23745 19907
rect 23624 19876 23745 19904
rect 23624 19864 23630 19876
rect 23733 19873 23745 19876
rect 23779 19873 23791 19907
rect 23733 19867 23791 19873
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18012 19808 18337 19836
rect 18012 19796 18018 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 23474 19836 23480 19848
rect 23435 19808 23480 19836
rect 18325 19799 18383 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 24857 19703 24915 19709
rect 24857 19669 24869 19703
rect 24903 19700 24915 19703
rect 24946 19700 24952 19712
rect 24903 19672 24952 19700
rect 24903 19669 24915 19672
rect 24857 19663 24915 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 13630 19320 13636 19372
rect 13688 19360 13694 19372
rect 13688 19332 13768 19360
rect 13688 19320 13694 19332
rect 8570 19292 8576 19304
rect 8531 19264 8576 19292
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 13740 19292 13768 19332
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 18380 19332 19257 19360
rect 18380 19320 18386 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 13740 19264 14565 19292
rect 14553 19261 14565 19264
rect 14599 19292 14611 19295
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14599 19264 15117 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 15105 19261 15117 19264
rect 15151 19292 15163 19295
rect 15838 19292 15844 19304
rect 15151 19264 15844 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15838 19252 15844 19264
rect 15896 19292 15902 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 15896 19264 17417 19292
rect 15896 19252 15902 19264
rect 17405 19261 17417 19264
rect 17451 19292 17463 19295
rect 17954 19292 17960 19304
rect 17451 19264 17960 19292
rect 17451 19261 17463 19264
rect 17405 19255 17463 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 23474 19252 23480 19304
rect 23532 19292 23538 19304
rect 24857 19295 24915 19301
rect 24857 19292 24869 19295
rect 23532 19264 24869 19292
rect 23532 19252 23538 19264
rect 8478 19224 8484 19236
rect 8391 19196 8484 19224
rect 8478 19184 8484 19196
rect 8536 19224 8542 19236
rect 8818 19227 8876 19233
rect 8818 19224 8830 19227
rect 8536 19196 8830 19224
rect 8536 19184 8542 19196
rect 8818 19193 8830 19196
rect 8864 19193 8876 19227
rect 15350 19227 15408 19233
rect 15350 19224 15362 19227
rect 8818 19187 8876 19193
rect 14936 19196 15362 19224
rect 9953 19159 10011 19165
rect 9953 19125 9965 19159
rect 9999 19156 10011 19159
rect 10318 19156 10324 19168
rect 9999 19128 10324 19156
rect 9999 19125 10011 19128
rect 9953 19119 10011 19125
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 14936 19165 14964 19196
rect 15350 19193 15362 19196
rect 15396 19193 15408 19227
rect 18598 19224 18604 19236
rect 18559 19196 18604 19224
rect 15350 19187 15408 19193
rect 18598 19184 18604 19196
rect 18656 19224 18662 19236
rect 19153 19227 19211 19233
rect 19153 19224 19165 19227
rect 18656 19196 19165 19224
rect 18656 19184 18662 19196
rect 19153 19193 19165 19196
rect 19199 19193 19211 19227
rect 19153 19187 19211 19193
rect 24412 19168 24440 19264
rect 24857 19261 24869 19264
rect 24903 19261 24915 19295
rect 24857 19255 24915 19261
rect 24765 19227 24823 19233
rect 24765 19193 24777 19227
rect 24811 19224 24823 19227
rect 24946 19224 24952 19236
rect 24811 19196 24952 19224
rect 24811 19193 24823 19196
rect 24765 19187 24823 19193
rect 24946 19184 24952 19196
rect 25004 19224 25010 19236
rect 25102 19227 25160 19233
rect 25102 19224 25114 19227
rect 25004 19196 25114 19224
rect 25004 19184 25010 19196
rect 25102 19193 25114 19196
rect 25148 19193 25160 19227
rect 25102 19187 25160 19193
rect 14921 19159 14979 19165
rect 14921 19156 14933 19159
rect 14884 19128 14933 19156
rect 14884 19116 14890 19128
rect 14921 19125 14933 19128
rect 14967 19125 14979 19159
rect 16482 19156 16488 19168
rect 16443 19128 16488 19156
rect 14921 19119 14979 19125
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 18322 19156 18328 19168
rect 17911 19128 18328 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 18690 19156 18696 19168
rect 18651 19128 18696 19156
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 18840 19128 19073 19156
rect 18840 19116 18846 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19061 19119 19119 19125
rect 23566 19116 23572 19168
rect 23624 19156 23630 19168
rect 23845 19159 23903 19165
rect 23845 19156 23857 19159
rect 23624 19128 23857 19156
rect 23624 19116 23630 19128
rect 23845 19125 23857 19128
rect 23891 19125 23903 19159
rect 23845 19119 23903 19125
rect 24305 19159 24363 19165
rect 24305 19125 24317 19159
rect 24351 19156 24363 19159
rect 24394 19156 24400 19168
rect 24351 19128 24400 19156
rect 24351 19125 24363 19128
rect 24305 19119 24363 19125
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 26237 19159 26295 19165
rect 26237 19156 26249 19159
rect 25740 19128 26249 19156
rect 25740 19116 25746 19128
rect 26237 19125 26249 19128
rect 26283 19125 26295 19159
rect 26237 19119 26295 19125
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 14090 18952 14096 18964
rect 14051 18924 14096 18952
rect 14090 18912 14096 18924
rect 14148 18952 14154 18964
rect 14458 18952 14464 18964
rect 14148 18924 14464 18952
rect 14148 18912 14154 18924
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 17865 18955 17923 18961
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 18782 18952 18788 18964
rect 17911 18924 18788 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 18782 18912 18788 18924
rect 18840 18912 18846 18964
rect 18877 18955 18935 18961
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 18923 18924 21281 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 21269 18921 21281 18924
rect 21315 18952 21327 18955
rect 21818 18952 21824 18964
rect 21315 18924 21824 18952
rect 21315 18921 21327 18924
rect 21269 18915 21327 18921
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 23937 18955 23995 18961
rect 23937 18921 23949 18955
rect 23983 18952 23995 18955
rect 24210 18952 24216 18964
rect 23983 18924 24216 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24210 18912 24216 18924
rect 24268 18952 24274 18964
rect 24946 18952 24952 18964
rect 24268 18924 24952 18952
rect 24268 18912 24274 18924
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 10686 18884 10692 18896
rect 10244 18856 10692 18884
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4321 18819 4379 18825
rect 4321 18816 4333 18819
rect 4212 18788 4333 18816
rect 4212 18776 4218 18788
rect 4321 18785 4333 18788
rect 4367 18785 4379 18819
rect 4321 18779 4379 18785
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 8665 18819 8723 18825
rect 8665 18816 8677 18819
rect 8628 18788 8677 18816
rect 8628 18776 8634 18788
rect 8665 18785 8677 18788
rect 8711 18816 8723 18819
rect 9214 18816 9220 18828
rect 8711 18788 9220 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 9214 18776 9220 18788
rect 9272 18816 9278 18828
rect 10244 18825 10272 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 18322 18884 18328 18896
rect 18283 18856 18328 18884
rect 18322 18844 18328 18856
rect 18380 18844 18386 18896
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 9272 18788 10241 18816
rect 9272 18776 9278 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10485 18819 10543 18825
rect 10485 18816 10497 18819
rect 10376 18788 10497 18816
rect 10376 18776 10382 18788
rect 10485 18785 10497 18788
rect 10531 18785 10543 18819
rect 10485 18779 10543 18785
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 12969 18819 13027 18825
rect 12969 18816 12981 18819
rect 12860 18788 12981 18816
rect 12860 18776 12866 18788
rect 12969 18785 12981 18788
rect 13015 18785 13027 18819
rect 12969 18779 13027 18785
rect 18690 18776 18696 18828
rect 18748 18816 18754 18828
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 18748 18788 19257 18816
rect 18748 18776 18754 18788
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 23198 18816 23204 18828
rect 23159 18788 23204 18816
rect 19245 18779 19303 18785
rect 23198 18776 23204 18788
rect 23256 18776 23262 18828
rect 23290 18776 23296 18828
rect 23348 18816 23354 18828
rect 23348 18788 23393 18816
rect 23348 18776 23354 18788
rect 1762 18748 1768 18760
rect 1723 18720 1768 18748
rect 1762 18708 1768 18720
rect 1820 18708 1826 18760
rect 4062 18748 4068 18760
rect 2240 18720 4068 18748
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 2240 18621 2268 18720
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 19337 18751 19395 18757
rect 19337 18748 19349 18751
rect 18932 18720 19349 18748
rect 18932 18708 18938 18720
rect 19337 18717 19349 18720
rect 19383 18717 19395 18751
rect 19337 18711 19395 18717
rect 19521 18751 19579 18757
rect 19521 18717 19533 18751
rect 19567 18748 19579 18751
rect 19702 18748 19708 18760
rect 19567 18720 19708 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18717 21419 18751
rect 21542 18748 21548 18760
rect 21503 18720 21548 18748
rect 21361 18711 21419 18717
rect 21266 18640 21272 18692
rect 21324 18680 21330 18692
rect 21376 18680 21404 18711
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 22738 18708 22744 18760
rect 22796 18748 22802 18760
rect 23477 18751 23535 18757
rect 23477 18748 23489 18751
rect 22796 18720 23489 18748
rect 22796 18708 22802 18720
rect 23477 18717 23489 18720
rect 23523 18748 23535 18751
rect 24302 18748 24308 18760
rect 23523 18720 24308 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 24302 18708 24308 18720
rect 24360 18748 24366 18760
rect 25682 18748 25688 18760
rect 24360 18720 25688 18748
rect 24360 18708 24366 18720
rect 25682 18708 25688 18720
rect 25740 18708 25746 18760
rect 21324 18652 21404 18680
rect 21324 18640 21330 18652
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 1544 18584 2237 18612
rect 1544 18572 1550 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 5442 18612 5448 18624
rect 5403 18584 5448 18612
rect 2225 18575 2283 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 7193 18615 7251 18621
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 7374 18612 7380 18624
rect 7239 18584 7380 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11609 18615 11667 18621
rect 11609 18612 11621 18615
rect 10928 18584 11621 18612
rect 10928 18572 10934 18584
rect 11609 18581 11621 18584
rect 11655 18612 11667 18615
rect 12710 18612 12716 18624
rect 11655 18584 12716 18612
rect 11655 18581 11667 18584
rect 11609 18575 11667 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 20438 18612 20444 18624
rect 20399 18584 20444 18612
rect 20438 18572 20444 18584
rect 20496 18572 20502 18624
rect 20901 18615 20959 18621
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21358 18612 21364 18624
rect 20947 18584 21364 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 22830 18612 22836 18624
rect 22791 18584 22836 18612
rect 22830 18572 22836 18584
rect 22888 18572 22894 18624
rect 24394 18572 24400 18624
rect 24452 18612 24458 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24452 18584 24961 18612
rect 24452 18572 24458 18584
rect 24949 18581 24961 18584
rect 24995 18612 25007 18615
rect 25774 18612 25780 18624
rect 24995 18584 25780 18612
rect 24995 18581 25007 18584
rect 24949 18575 25007 18581
rect 25774 18572 25780 18584
rect 25832 18572 25838 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 4433 18411 4491 18417
rect 4433 18408 4445 18411
rect 4120 18380 4445 18408
rect 4120 18368 4126 18380
rect 4433 18377 4445 18380
rect 4479 18408 4491 18411
rect 5626 18408 5632 18420
rect 4479 18380 5632 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 5626 18368 5632 18380
rect 5684 18408 5690 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 5684 18380 6561 18408
rect 5684 18368 5690 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 6549 18371 6607 18377
rect 3237 18343 3295 18349
rect 3237 18309 3249 18343
rect 3283 18340 3295 18343
rect 3786 18340 3792 18352
rect 3283 18312 3792 18340
rect 3283 18309 3295 18312
rect 3237 18303 3295 18309
rect 3786 18300 3792 18312
rect 3844 18340 3850 18352
rect 4154 18340 4160 18352
rect 3844 18312 4160 18340
rect 3844 18300 3850 18312
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 6564 18272 6592 18371
rect 8478 18368 8484 18380
rect 8536 18408 8542 18420
rect 9582 18408 9588 18420
rect 8536 18380 9588 18408
rect 8536 18368 8542 18380
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 10686 18408 10692 18420
rect 10647 18380 10692 18408
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 12802 18408 12808 18420
rect 12763 18380 12808 18408
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 17865 18411 17923 18417
rect 17865 18377 17877 18411
rect 17911 18408 17923 18411
rect 18690 18408 18696 18420
rect 17911 18380 18696 18408
rect 17911 18377 17923 18380
rect 17865 18371 17923 18377
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 18874 18408 18880 18420
rect 18835 18380 18880 18408
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 19702 18368 19708 18420
rect 19760 18408 19766 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 19760 18380 19901 18408
rect 19760 18368 19766 18380
rect 19889 18377 19901 18380
rect 19935 18408 19947 18411
rect 20257 18411 20315 18417
rect 20257 18408 20269 18411
rect 19935 18380 20269 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 20257 18377 20269 18380
rect 20303 18377 20315 18411
rect 21542 18408 21548 18420
rect 21503 18380 21548 18408
rect 20257 18371 20315 18377
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 13081 18343 13139 18349
rect 13081 18340 13093 18343
rect 12676 18312 13093 18340
rect 12676 18300 12682 18312
rect 13081 18309 13093 18312
rect 13127 18309 13139 18343
rect 13081 18303 13139 18309
rect 13998 18300 14004 18352
rect 14056 18340 14062 18352
rect 14277 18343 14335 18349
rect 14277 18340 14289 18343
rect 14056 18312 14289 18340
rect 14056 18300 14062 18312
rect 14277 18309 14289 18312
rect 14323 18309 14335 18343
rect 18322 18340 18328 18352
rect 18283 18312 18328 18340
rect 14277 18303 14335 18309
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6564 18244 7113 18272
rect 7101 18241 7113 18244
rect 7147 18241 7159 18275
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 7101 18235 7159 18241
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 18340 18272 18368 18300
rect 19429 18275 19487 18281
rect 19429 18272 19441 18275
rect 18340 18244 19441 18272
rect 19429 18241 19441 18244
rect 19475 18241 19487 18275
rect 20272 18272 20300 18371
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 21818 18408 21824 18420
rect 21779 18380 21824 18408
rect 21818 18368 21824 18380
rect 21876 18368 21882 18420
rect 22373 18411 22431 18417
rect 22373 18377 22385 18411
rect 22419 18408 22431 18411
rect 23198 18408 23204 18420
rect 22419 18380 23204 18408
rect 22419 18377 22431 18380
rect 22373 18371 22431 18377
rect 23198 18368 23204 18380
rect 23256 18408 23262 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23256 18380 23673 18408
rect 23256 18368 23262 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 25222 18368 25228 18420
rect 25280 18408 25286 18420
rect 25498 18408 25504 18420
rect 25280 18380 25504 18408
rect 25280 18368 25286 18380
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 20441 18343 20499 18349
rect 20441 18309 20453 18343
rect 20487 18340 20499 18343
rect 21266 18340 21272 18352
rect 20487 18312 21272 18340
rect 20487 18309 20499 18312
rect 20441 18303 20499 18309
rect 21266 18300 21272 18312
rect 21324 18300 21330 18352
rect 22738 18340 22744 18352
rect 22699 18312 22744 18340
rect 22738 18300 22744 18312
rect 22796 18300 22802 18352
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20272 18244 21005 18272
rect 19429 18235 19487 18241
rect 20993 18241 21005 18244
rect 21039 18241 21051 18275
rect 24210 18272 24216 18284
rect 24171 18244 24216 18272
rect 20993 18235 21051 18241
rect 24210 18232 24216 18244
rect 24268 18232 24274 18284
rect 25682 18272 25688 18284
rect 25643 18244 25688 18272
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 1486 18164 1492 18216
rect 1544 18204 1550 18216
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1544 18176 1869 18204
rect 1544 18164 1550 18176
rect 1857 18173 1869 18176
rect 1903 18173 1915 18207
rect 14645 18207 14703 18213
rect 14645 18204 14657 18207
rect 1857 18167 1915 18173
rect 13832 18176 14657 18204
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 2124 18139 2182 18145
rect 2124 18136 2136 18139
rect 1811 18108 2136 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 2124 18105 2136 18108
rect 2170 18136 2182 18139
rect 2498 18136 2504 18148
rect 2170 18108 2504 18136
rect 2170 18105 2182 18108
rect 2124 18099 2182 18105
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 7374 18145 7380 18148
rect 7368 18136 7380 18145
rect 7335 18108 7380 18136
rect 7368 18099 7380 18108
rect 7374 18096 7380 18099
rect 7432 18096 7438 18148
rect 13832 18080 13860 18176
rect 14645 18173 14657 18176
rect 14691 18173 14703 18207
rect 14645 18167 14703 18173
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 20438 18204 20444 18216
rect 19392 18176 20444 18204
rect 19392 18164 19398 18176
rect 20438 18164 20444 18176
rect 20496 18204 20502 18216
rect 20809 18207 20867 18213
rect 20809 18204 20821 18207
rect 20496 18176 20821 18204
rect 20496 18164 20502 18176
rect 20809 18173 20821 18176
rect 20855 18173 20867 18207
rect 23474 18204 23480 18216
rect 23387 18176 23480 18204
rect 20809 18167 20867 18173
rect 23474 18164 23480 18176
rect 23532 18204 23538 18216
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23532 18176 24133 18204
rect 23532 18164 23538 18176
rect 24121 18173 24133 18176
rect 24167 18204 24179 18207
rect 24762 18204 24768 18216
rect 24167 18176 24768 18204
rect 24167 18173 24179 18176
rect 24121 18167 24179 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 25784 18207 25842 18213
rect 25784 18204 25796 18207
rect 25608 18176 25796 18204
rect 14734 18136 14740 18148
rect 14695 18108 14740 18136
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 19150 18096 19156 18148
rect 19208 18136 19214 18148
rect 19208 18108 19380 18136
rect 19208 18096 19214 18108
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 9824 18040 10241 18068
rect 9824 18028 9830 18040
rect 10229 18037 10241 18040
rect 10275 18068 10287 18071
rect 10318 18068 10324 18080
rect 10275 18040 10324 18068
rect 10275 18037 10287 18040
rect 10229 18031 10287 18037
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14185 18071 14243 18077
rect 14185 18068 14197 18071
rect 13964 18040 14197 18068
rect 13964 18028 13970 18040
rect 14185 18037 14197 18040
rect 14231 18068 14243 18071
rect 14752 18068 14780 18096
rect 14231 18040 14780 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19352 18077 19380 18108
rect 22186 18096 22192 18148
rect 22244 18136 22250 18148
rect 23109 18139 23167 18145
rect 23109 18136 23121 18139
rect 22244 18108 23121 18136
rect 22244 18096 22250 18108
rect 23109 18105 23121 18108
rect 23155 18136 23167 18139
rect 24029 18139 24087 18145
rect 24029 18136 24041 18139
rect 23155 18108 24041 18136
rect 23155 18105 23167 18108
rect 23109 18099 23167 18105
rect 24029 18105 24041 18108
rect 24075 18105 24087 18139
rect 24029 18099 24087 18105
rect 18693 18071 18751 18077
rect 18693 18068 18705 18071
rect 18656 18040 18705 18068
rect 18656 18028 18662 18040
rect 18693 18037 18705 18040
rect 18739 18068 18751 18071
rect 19245 18071 19303 18077
rect 19245 18068 19257 18071
rect 18739 18040 19257 18068
rect 18739 18037 18751 18040
rect 18693 18031 18751 18037
rect 19245 18037 19257 18040
rect 19291 18037 19303 18071
rect 19245 18031 19303 18037
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18037 19395 18071
rect 19337 18031 19395 18037
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20772 18040 20913 18068
rect 20772 18028 20778 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 25608 18068 25636 18176
rect 25784 18173 25796 18176
rect 25830 18173 25842 18207
rect 25784 18167 25842 18173
rect 25682 18096 25688 18148
rect 25740 18136 25746 18148
rect 26022 18139 26080 18145
rect 26022 18136 26034 18139
rect 25740 18108 26034 18136
rect 25740 18096 25746 18108
rect 26022 18105 26034 18108
rect 26068 18105 26080 18139
rect 26022 18099 26080 18105
rect 25774 18068 25780 18080
rect 25608 18040 25780 18068
rect 20901 18031 20959 18037
rect 25774 18028 25780 18040
rect 25832 18028 25838 18080
rect 27154 18068 27160 18080
rect 27115 18040 27160 18068
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2225 17867 2283 17873
rect 2225 17864 2237 17867
rect 1820 17836 2237 17864
rect 1820 17824 1826 17836
rect 2225 17833 2237 17836
rect 2271 17864 2283 17867
rect 2958 17864 2964 17876
rect 2271 17836 2964 17864
rect 2271 17833 2283 17836
rect 2225 17827 2283 17833
rect 2958 17824 2964 17836
rect 3016 17824 3022 17876
rect 12621 17867 12679 17873
rect 12621 17833 12633 17867
rect 12667 17864 12679 17867
rect 13722 17864 13728 17876
rect 12667 17836 13728 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 18601 17867 18659 17873
rect 18601 17833 18613 17867
rect 18647 17864 18659 17867
rect 18874 17864 18880 17876
rect 18647 17836 18880 17864
rect 18647 17833 18659 17836
rect 18601 17827 18659 17833
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 19242 17864 19248 17876
rect 19203 17836 19248 17864
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 20533 17867 20591 17873
rect 20533 17833 20545 17867
rect 20579 17864 20591 17867
rect 20622 17864 20628 17876
rect 20579 17836 20628 17864
rect 20579 17833 20591 17836
rect 20533 17827 20591 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 21177 17867 21235 17873
rect 21177 17833 21189 17867
rect 21223 17864 21235 17867
rect 21266 17864 21272 17876
rect 21223 17836 21272 17864
rect 21223 17833 21235 17836
rect 21177 17827 21235 17833
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17864 22155 17867
rect 22370 17864 22376 17876
rect 22143 17836 22376 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 22370 17824 22376 17836
rect 22428 17864 22434 17876
rect 22830 17864 22836 17876
rect 22428 17836 22836 17864
rect 22428 17824 22434 17836
rect 22830 17824 22836 17836
rect 22888 17824 22894 17876
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17864 22983 17867
rect 23201 17867 23259 17873
rect 23201 17864 23213 17867
rect 22971 17836 23213 17864
rect 22971 17833 22983 17836
rect 22925 17827 22983 17833
rect 23201 17833 23213 17836
rect 23247 17864 23259 17867
rect 23290 17864 23296 17876
rect 23247 17836 23296 17864
rect 23247 17833 23259 17836
rect 23201 17827 23259 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 5442 17756 5448 17808
rect 5500 17796 5506 17808
rect 5874 17799 5932 17805
rect 5874 17796 5886 17799
rect 5500 17768 5886 17796
rect 5500 17756 5506 17768
rect 5874 17765 5886 17768
rect 5920 17765 5932 17799
rect 5874 17759 5932 17765
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 16384 17799 16442 17805
rect 16384 17796 16396 17799
rect 13504 17768 16396 17796
rect 13504 17756 13510 17768
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 5626 17728 5632 17740
rect 5587 17700 5632 17728
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10468 17700 10517 17728
rect 10468 17688 10474 17700
rect 10505 17697 10517 17700
rect 10551 17728 10563 17731
rect 11054 17728 11060 17740
rect 10551 17700 11060 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 13998 17728 14004 17740
rect 13959 17700 14004 17728
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 2498 17660 2504 17672
rect 2459 17632 2504 17660
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10008 17632 10609 17660
rect 10008 17620 10014 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 10689 17623 10747 17629
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 10226 17592 10232 17604
rect 9732 17564 10232 17592
rect 9732 17552 9738 17564
rect 10226 17552 10232 17564
rect 10284 17592 10290 17604
rect 10704 17592 10732 17623
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14200 17669 14228 17768
rect 16384 17765 16396 17768
rect 16430 17796 16442 17799
rect 16482 17796 16488 17808
rect 16430 17768 16488 17796
rect 16430 17765 16442 17768
rect 16384 17759 16442 17765
rect 16482 17756 16488 17768
rect 16540 17756 16546 17808
rect 18969 17799 19027 17805
rect 18969 17765 18981 17799
rect 19015 17796 19027 17799
rect 19150 17796 19156 17808
rect 19015 17768 19156 17796
rect 19015 17765 19027 17768
rect 18969 17759 19027 17765
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 22186 17796 22192 17808
rect 22147 17768 22192 17796
rect 22186 17756 22192 17768
rect 22244 17756 22250 17808
rect 15838 17688 15844 17740
rect 15896 17728 15902 17740
rect 16117 17731 16175 17737
rect 16117 17728 16129 17731
rect 15896 17700 16129 17728
rect 15896 17688 15902 17700
rect 16117 17697 16129 17700
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19613 17731 19671 17737
rect 19613 17728 19625 17731
rect 19392 17700 19625 17728
rect 19392 17688 19398 17700
rect 19613 17697 19625 17700
rect 19659 17697 19671 17731
rect 19613 17691 19671 17697
rect 23198 17688 23204 17740
rect 23256 17728 23262 17740
rect 23569 17731 23627 17737
rect 23569 17728 23581 17731
rect 23256 17700 23581 17728
rect 23256 17688 23262 17700
rect 23569 17697 23581 17700
rect 23615 17697 23627 17731
rect 23569 17691 23627 17697
rect 23658 17688 23664 17740
rect 23716 17728 23722 17740
rect 24762 17728 24768 17740
rect 23716 17700 24768 17728
rect 23716 17688 23722 17700
rect 24762 17688 24768 17700
rect 24820 17688 24826 17740
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17629 14243 17663
rect 19702 17660 19708 17672
rect 19663 17632 19708 17660
rect 14185 17623 14243 17629
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 23842 17660 23848 17672
rect 23755 17632 23848 17660
rect 19797 17623 19855 17629
rect 10284 17564 10732 17592
rect 10284 17552 10290 17564
rect 18322 17552 18328 17604
rect 18380 17592 18386 17604
rect 19812 17592 19840 17623
rect 23842 17620 23848 17632
rect 23900 17660 23906 17672
rect 24210 17660 24216 17672
rect 23900 17632 24216 17660
rect 23900 17620 23906 17632
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 19978 17592 19984 17604
rect 18380 17564 19984 17592
rect 18380 17552 18386 17564
rect 19978 17552 19984 17564
rect 20036 17552 20042 17604
rect 1762 17524 1768 17536
rect 1723 17496 1768 17524
rect 1762 17484 1768 17496
rect 1820 17484 1826 17536
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 2314 17524 2320 17536
rect 1903 17496 2320 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 2314 17484 2320 17496
rect 2372 17524 2378 17536
rect 2869 17527 2927 17533
rect 2869 17524 2881 17527
rect 2372 17496 2881 17524
rect 2372 17484 2378 17496
rect 2869 17493 2881 17496
rect 2915 17493 2927 17527
rect 4430 17524 4436 17536
rect 4391 17496 4436 17524
rect 2869 17487 2927 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 4706 17524 4712 17536
rect 4667 17496 4712 17524
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 7374 17524 7380 17536
rect 7055 17496 7380 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9824 17496 9965 17524
rect 9824 17484 9830 17496
rect 9953 17493 9965 17496
rect 9999 17493 10011 17527
rect 10134 17524 10140 17536
rect 10095 17496 10140 17524
rect 9953 17487 10011 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 13630 17524 13636 17536
rect 13591 17496 13636 17524
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 14734 17524 14740 17536
rect 14695 17496 14740 17524
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 24213 17527 24271 17533
rect 24213 17524 24225 17527
rect 24176 17496 24225 17524
rect 24176 17484 24182 17496
rect 24213 17493 24225 17496
rect 24259 17493 24271 17527
rect 24213 17487 24271 17493
rect 25682 17484 25688 17536
rect 25740 17524 25746 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 25740 17496 25789 17524
rect 25740 17484 25746 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 25777 17487 25835 17493
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1670 17280 1676 17332
rect 1728 17320 1734 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 1728 17292 1869 17320
rect 1728 17280 1734 17292
rect 1857 17289 1869 17292
rect 1903 17320 1915 17323
rect 2222 17320 2228 17332
rect 1903 17292 2228 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 3786 17320 3792 17332
rect 3747 17292 3792 17320
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5500 17292 5641 17320
rect 5500 17280 5506 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 5629 17283 5687 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 15289 17323 15347 17329
rect 15289 17320 15301 17323
rect 14056 17292 15301 17320
rect 14056 17280 14062 17292
rect 15289 17289 15301 17292
rect 15335 17289 15347 17323
rect 15289 17283 15347 17289
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16482 17320 16488 17332
rect 16255 17292 16488 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 18509 17323 18567 17329
rect 18509 17320 18521 17323
rect 18380 17292 18521 17320
rect 18380 17280 18386 17292
rect 18509 17289 18521 17292
rect 18555 17320 18567 17323
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 18555 17292 18889 17320
rect 18555 17289 18567 17292
rect 18509 17283 18567 17289
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 19334 17320 19340 17332
rect 19295 17292 19340 17320
rect 18877 17283 18935 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 20622 17320 20628 17332
rect 19475 17292 20628 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 24762 17320 24768 17332
rect 24723 17292 24768 17320
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 1762 17144 1768 17196
rect 1820 17184 1826 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 1820 17156 2421 17184
rect 1820 17144 1826 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17184 2651 17187
rect 3804 17184 3832 17280
rect 4249 17255 4307 17261
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 4295 17224 5028 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 4154 17184 4160 17196
rect 2639 17156 4160 17184
rect 2639 17153 2651 17156
rect 2593 17147 2651 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 5000 17193 5028 17224
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4488 17156 4813 17184
rect 4488 17144 4494 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17184 5043 17187
rect 5460 17184 5488 17280
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 13081 17255 13139 17261
rect 9824 17224 10548 17252
rect 9824 17212 9830 17224
rect 5031 17156 5488 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 5626 17144 5632 17196
rect 5684 17184 5690 17196
rect 5997 17187 6055 17193
rect 5997 17184 6009 17187
rect 5684 17156 6009 17184
rect 5684 17144 5690 17156
rect 5997 17153 6009 17156
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 10134 17184 10140 17196
rect 9539 17156 10140 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10134 17144 10140 17156
rect 10192 17184 10198 17196
rect 10520 17193 10548 17224
rect 13081 17221 13093 17255
rect 13127 17252 13139 17255
rect 14090 17252 14096 17264
rect 13127 17224 14096 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 14090 17212 14096 17224
rect 14148 17252 14154 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 14148 17224 14289 17252
rect 14148 17212 14154 17224
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 23661 17255 23719 17261
rect 23661 17252 23673 17255
rect 14277 17215 14335 17221
rect 22480 17224 23673 17252
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10192 17156 10425 17184
rect 10192 17144 10198 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 14792 17156 14841 17184
rect 14792 17144 14798 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16485 17187 16543 17193
rect 16485 17184 16497 17187
rect 15896 17156 16497 17184
rect 15896 17144 15902 17156
rect 16485 17153 16497 17156
rect 16531 17184 16543 17187
rect 16666 17184 16672 17196
rect 16531 17156 16672 17184
rect 16531 17153 16543 17156
rect 16485 17147 16543 17153
rect 16666 17144 16672 17156
rect 16724 17184 16730 17196
rect 18138 17184 18144 17196
rect 16724 17156 18144 17184
rect 16724 17144 16730 17156
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 19978 17184 19984 17196
rect 19939 17156 19984 17184
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 22480 17193 22508 17224
rect 23661 17221 23673 17224
rect 23707 17221 23719 17255
rect 23661 17215 23719 17221
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 22152 17156 22477 17184
rect 22152 17144 22158 17156
rect 22465 17153 22477 17156
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 22649 17187 22707 17193
rect 22649 17153 22661 17187
rect 22695 17153 22707 17187
rect 24118 17184 24124 17196
rect 24079 17156 24124 17184
rect 22649 17147 22707 17153
rect 2314 17116 2320 17128
rect 2275 17088 2320 17116
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 9950 17116 9956 17128
rect 9907 17088 9956 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 11054 17116 11060 17128
rect 10967 17088 11060 17116
rect 11054 17076 11060 17088
rect 11112 17116 11118 17128
rect 12986 17116 12992 17128
rect 11112 17088 12992 17116
rect 11112 17076 11118 17088
rect 12986 17076 12992 17088
rect 13044 17076 13050 17128
rect 22370 17116 22376 17128
rect 22331 17088 22376 17116
rect 22370 17076 22376 17088
rect 22428 17076 22434 17128
rect 22664 17116 22692 17147
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 24302 17184 24308 17196
rect 24263 17156 24308 17184
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17184 25927 17187
rect 25915 17156 26096 17184
rect 25915 17153 25927 17156
rect 25869 17147 25927 17153
rect 25884 17116 25912 17147
rect 22664 17088 25912 17116
rect 25961 17119 26019 17125
rect 4706 17048 4712 17060
rect 1964 17020 4712 17048
rect 1964 16989 1992 17020
rect 4706 17008 4712 17020
rect 4764 17008 4770 17060
rect 9125 17051 9183 17057
rect 9125 17017 9137 17051
rect 9171 17048 9183 17051
rect 10321 17051 10379 17057
rect 10321 17048 10333 17051
rect 9171 17020 10333 17048
rect 9171 17017 9183 17020
rect 9125 17011 9183 17017
rect 10321 17017 10333 17020
rect 10367 17048 10379 17051
rect 10410 17048 10416 17060
rect 10367 17020 10416 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 10410 17008 10416 17020
rect 10468 17008 10474 17060
rect 13817 17051 13875 17057
rect 13817 17017 13829 17051
rect 13863 17048 13875 17051
rect 13863 17020 14780 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 1949 16983 2007 16989
rect 1949 16949 1961 16983
rect 1995 16949 2007 16983
rect 1949 16943 2007 16949
rect 3421 16983 3479 16989
rect 3421 16949 3433 16983
rect 3467 16980 3479 16983
rect 3694 16980 3700 16992
rect 3467 16952 3700 16980
rect 3467 16949 3479 16952
rect 3421 16943 3479 16949
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 4338 16980 4344 16992
rect 4299 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 10778 16980 10784 16992
rect 9999 16952 10784 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 14182 16980 14188 16992
rect 14095 16952 14188 16980
rect 14182 16940 14188 16952
rect 14240 16980 14246 16992
rect 14642 16980 14648 16992
rect 14240 16952 14648 16980
rect 14240 16940 14246 16952
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 14752 16989 14780 17020
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20809 17051 20867 17057
rect 20809 17048 20821 17051
rect 19760 17020 20821 17048
rect 19760 17008 19766 17020
rect 20809 17017 20821 17020
rect 20855 17017 20867 17051
rect 20809 17011 20867 17017
rect 21913 17051 21971 17057
rect 21913 17017 21925 17051
rect 21959 17048 21971 17051
rect 22664 17048 22692 17088
rect 25961 17085 25973 17119
rect 26007 17085 26019 17119
rect 26068 17116 26096 17156
rect 26228 17119 26286 17125
rect 26228 17116 26240 17119
rect 26068 17088 26240 17116
rect 25961 17079 26019 17085
rect 26228 17085 26240 17088
rect 26274 17116 26286 17119
rect 27154 17116 27160 17128
rect 26274 17088 27160 17116
rect 26274 17085 26286 17088
rect 26228 17079 26286 17085
rect 23198 17048 23204 17060
rect 21959 17020 22692 17048
rect 23159 17020 23204 17048
rect 21959 17017 21971 17020
rect 21913 17011 21971 17017
rect 23198 17008 23204 17020
rect 23256 17008 23262 17060
rect 24026 17048 24032 17060
rect 23939 17020 24032 17048
rect 24026 17008 24032 17020
rect 24084 17048 24090 17060
rect 25041 17051 25099 17057
rect 25041 17048 25053 17051
rect 24084 17020 25053 17048
rect 24084 17008 24090 17020
rect 25041 17017 25053 17020
rect 25087 17017 25099 17051
rect 25041 17011 25099 17017
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 25976 17048 26004 17079
rect 27154 17076 27160 17088
rect 27212 17076 27218 17128
rect 25740 17020 26004 17048
rect 25740 17008 25746 17020
rect 14737 16983 14795 16989
rect 14737 16949 14749 16983
rect 14783 16980 14795 16983
rect 14826 16980 14832 16992
rect 14783 16952 14832 16980
rect 14783 16949 14795 16952
rect 14737 16943 14795 16949
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 19794 16980 19800 16992
rect 19755 16952 19800 16980
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19944 16952 20453 16980
rect 19944 16940 19950 16952
rect 20441 16949 20453 16952
rect 20487 16949 20499 16983
rect 22002 16980 22008 16992
rect 21963 16952 22008 16980
rect 20441 16943 20499 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 27338 16980 27344 16992
rect 27299 16952 27344 16980
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1820 16748 1961 16776
rect 1820 16736 1826 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 1949 16739 2007 16745
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2682 16776 2688 16788
rect 2455 16748 2688 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16776 4123 16779
rect 4430 16776 4436 16788
rect 4111 16748 4436 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 10226 16776 10232 16788
rect 10187 16748 10232 16776
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10686 16776 10692 16788
rect 10459 16748 10692 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 13173 16779 13231 16785
rect 10836 16748 10881 16776
rect 10836 16736 10842 16748
rect 13173 16745 13185 16779
rect 13219 16776 13231 16779
rect 13630 16776 13636 16788
rect 13219 16748 13636 16776
rect 13219 16745 13231 16748
rect 13173 16739 13231 16745
rect 13630 16736 13636 16748
rect 13688 16776 13694 16788
rect 14001 16779 14059 16785
rect 14001 16776 14013 16779
rect 13688 16748 14013 16776
rect 13688 16736 13694 16748
rect 14001 16745 14013 16748
rect 14047 16745 14059 16779
rect 14001 16739 14059 16745
rect 19521 16779 19579 16785
rect 19521 16745 19533 16779
rect 19567 16776 19579 16779
rect 19978 16776 19984 16788
rect 19567 16748 19984 16776
rect 19567 16745 19579 16748
rect 19521 16739 19579 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 23201 16779 23259 16785
rect 22152 16748 22197 16776
rect 22152 16736 22158 16748
rect 23201 16745 23213 16779
rect 23247 16776 23259 16779
rect 24026 16776 24032 16788
rect 23247 16748 24032 16776
rect 23247 16745 23259 16748
rect 23201 16739 23259 16745
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 24302 16776 24308 16788
rect 24263 16748 24308 16776
rect 24302 16736 24308 16748
rect 24360 16736 24366 16788
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2406 16640 2412 16652
rect 2363 16612 2412 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4890 16640 4896 16652
rect 4479 16612 4896 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 7193 16643 7251 16649
rect 7193 16640 7205 16643
rect 6840 16612 7205 16640
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 2593 16575 2651 16581
rect 2593 16572 2605 16575
rect 2556 16544 2605 16572
rect 2556 16532 2562 16544
rect 2593 16541 2605 16544
rect 2639 16541 2651 16575
rect 4522 16572 4528 16584
rect 4483 16544 4528 16572
rect 2593 16535 2651 16541
rect 2608 16504 2636 16535
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 3053 16507 3111 16513
rect 3053 16504 3065 16507
rect 2608 16476 3065 16504
rect 3053 16473 3065 16476
rect 3099 16504 3111 16507
rect 3694 16504 3700 16516
rect 3099 16476 3700 16504
rect 3099 16473 3111 16476
rect 3053 16467 3111 16473
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 4632 16504 4660 16535
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 6840 16572 6868 16612
rect 7193 16609 7205 16612
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 10796 16640 10824 16736
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 11977 16711 12035 16717
rect 11977 16708 11989 16711
rect 11020 16680 11989 16708
rect 11020 16668 11026 16680
rect 11977 16677 11989 16680
rect 12023 16677 12035 16711
rect 11977 16671 12035 16677
rect 23109 16711 23167 16717
rect 23109 16677 23121 16711
rect 23155 16708 23167 16711
rect 23842 16708 23848 16720
rect 23155 16680 23848 16708
rect 23155 16677 23167 16680
rect 23109 16671 23167 16677
rect 23842 16668 23848 16680
rect 23900 16668 23906 16720
rect 11054 16640 11060 16652
rect 9732 16612 10732 16640
rect 10796 16612 11060 16640
rect 9732 16600 9738 16612
rect 7282 16572 7288 16584
rect 6696 16544 6868 16572
rect 7243 16544 7288 16572
rect 6696 16532 6702 16544
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 10704 16572 10732 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13722 16640 13728 16652
rect 13587 16612 13728 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13832 16612 14105 16640
rect 10870 16572 10876 16584
rect 7432 16544 7477 16572
rect 10704 16544 10876 16572
rect 7432 16532 7438 16544
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 13832 16572 13860 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 18138 16640 18144 16652
rect 18099 16612 18144 16640
rect 14093 16603 14151 16609
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 18414 16649 18420 16652
rect 18408 16640 18420 16649
rect 18375 16612 18420 16640
rect 18408 16603 18420 16612
rect 18414 16600 18420 16603
rect 18472 16600 18478 16652
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 19852 16612 20177 16640
rect 19852 16600 19858 16612
rect 20165 16609 20177 16612
rect 20211 16640 20223 16643
rect 20211 16612 20668 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 10965 16535 11023 16541
rect 13556 16544 13860 16572
rect 14277 16575 14335 16581
rect 4212 16476 4660 16504
rect 4212 16464 4218 16476
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 10980 16504 11008 16535
rect 13556 16516 13584 16544
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14366 16572 14372 16584
rect 14323 16544 14372 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 20640 16572 20668 16612
rect 23474 16600 23480 16652
rect 23532 16640 23538 16652
rect 23569 16643 23627 16649
rect 23569 16640 23581 16643
rect 23532 16612 23581 16640
rect 23532 16600 23538 16612
rect 23569 16609 23581 16612
rect 23615 16609 23627 16643
rect 26510 16640 26516 16652
rect 26471 16612 26516 16640
rect 23569 16603 23627 16609
rect 26510 16600 26516 16612
rect 26568 16600 26574 16652
rect 21450 16572 21456 16584
rect 20640 16544 21456 16572
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23842 16572 23848 16584
rect 23803 16544 23848 16572
rect 23661 16535 23719 16541
rect 10836 16476 11008 16504
rect 10836 16464 10842 16476
rect 13538 16464 13544 16516
rect 13596 16464 13602 16516
rect 22738 16464 22744 16516
rect 22796 16504 22802 16516
rect 23676 16504 23704 16535
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 26418 16504 26424 16516
rect 22796 16476 26424 16504
rect 22796 16464 22802 16476
rect 26418 16464 26424 16476
rect 26476 16464 26482 16516
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 3602 16436 3608 16448
rect 3467 16408 3608 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 6825 16439 6883 16445
rect 6825 16405 6837 16439
rect 6871 16436 6883 16439
rect 7742 16436 7748 16448
rect 6871 16408 7748 16436
rect 6871 16405 6883 16408
rect 6825 16399 6883 16405
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 8938 16436 8944 16448
rect 8899 16408 8944 16436
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 13630 16436 13636 16448
rect 13591 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14734 16436 14740 16448
rect 14695 16408 14740 16436
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 21453 16439 21511 16445
rect 21453 16436 21465 16439
rect 20496 16408 21465 16436
rect 20496 16396 20502 16408
rect 21453 16405 21465 16408
rect 21499 16405 21511 16439
rect 21453 16399 21511 16405
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 25961 16439 26019 16445
rect 25961 16436 25973 16439
rect 25740 16408 25973 16436
rect 25740 16396 25746 16408
rect 25961 16405 25973 16408
rect 26007 16405 26019 16439
rect 26694 16436 26700 16448
rect 26655 16408 26700 16436
rect 25961 16399 26019 16405
rect 26694 16396 26700 16408
rect 26752 16396 26758 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 2041 16235 2099 16241
rect 2041 16201 2053 16235
rect 2087 16232 2099 16235
rect 2406 16232 2412 16244
rect 2087 16204 2412 16232
rect 2087 16201 2099 16204
rect 2041 16195 2099 16201
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7101 16235 7159 16241
rect 7101 16232 7113 16235
rect 6972 16204 7113 16232
rect 6972 16192 6978 16204
rect 7101 16201 7113 16204
rect 7147 16232 7159 16235
rect 7282 16232 7288 16244
rect 7147 16204 7288 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 9674 16232 9680 16244
rect 8895 16204 9680 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10410 16232 10416 16244
rect 10371 16204 10416 16232
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11112 16204 11805 16232
rect 11112 16192 11118 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13596 16204 13737 16232
rect 13596 16192 13602 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 18138 16232 18144 16244
rect 17911 16204 18144 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18138 16192 18144 16204
rect 18196 16232 18202 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18196 16204 18797 16232
rect 18196 16192 18202 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 19886 16232 19892 16244
rect 19847 16204 19892 16232
rect 18785 16195 18843 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 21450 16232 21456 16244
rect 21411 16204 21456 16232
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 22738 16232 22744 16244
rect 22699 16204 22744 16232
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23661 16235 23719 16241
rect 23661 16201 23673 16235
rect 23707 16232 23719 16235
rect 24118 16232 24124 16244
rect 23707 16204 24124 16232
rect 23707 16201 23719 16204
rect 23661 16195 23719 16201
rect 24118 16192 24124 16204
rect 24176 16192 24182 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 25406 16232 25412 16244
rect 25004 16204 25412 16232
rect 25004 16192 25010 16204
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 26510 16232 26516 16244
rect 26471 16204 26516 16232
rect 26510 16192 26516 16204
rect 26568 16192 26574 16244
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16164 3203 16167
rect 4522 16164 4528 16176
rect 3191 16136 4528 16164
rect 3191 16133 3203 16136
rect 3145 16127 3203 16133
rect 4522 16124 4528 16136
rect 4580 16124 4586 16176
rect 13633 16167 13691 16173
rect 13633 16133 13645 16167
rect 13679 16164 13691 16167
rect 14366 16164 14372 16176
rect 13679 16136 14372 16164
rect 13679 16133 13691 16136
rect 13633 16127 13691 16133
rect 14366 16124 14372 16136
rect 14424 16124 14430 16176
rect 15289 16167 15347 16173
rect 15289 16133 15301 16167
rect 15335 16133 15347 16167
rect 15289 16127 15347 16133
rect 3694 16096 3700 16108
rect 3655 16068 3700 16096
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 7742 16096 7748 16108
rect 7703 16068 7748 16096
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 7926 16096 7932 16108
rect 7839 16068 7932 16096
rect 7926 16056 7932 16068
rect 7984 16096 7990 16108
rect 8478 16096 8484 16108
rect 7984 16068 8484 16096
rect 7984 16056 7990 16068
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16096 8815 16099
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 8803 16068 9413 16096
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 9401 16065 9413 16068
rect 9447 16096 9459 16099
rect 9766 16096 9772 16108
rect 9447 16068 9772 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10284 16068 10977 16096
rect 10284 16056 10290 16068
rect 10965 16065 10977 16068
rect 11011 16096 11023 16099
rect 11425 16099 11483 16105
rect 11425 16096 11437 16099
rect 11011 16068 11437 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 11425 16065 11437 16068
rect 11471 16065 11483 16099
rect 11425 16059 11483 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13446 16096 13452 16108
rect 13311 16068 13452 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13446 16056 13452 16068
rect 13504 16096 13510 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 13504 16068 14289 16096
rect 13504 16056 13510 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1670 16028 1676 16040
rect 1443 16000 1676 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 3602 16028 3608 16040
rect 2832 16000 3608 16028
rect 2832 15988 2838 16000
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 7760 16028 7788 16056
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7760 16000 8309 16028
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 8996 16000 9229 16028
rect 8996 15988 9002 16000
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13872 16000 14105 16028
rect 13872 15988 13878 16000
rect 14093 15997 14105 16000
rect 14139 16028 14151 16031
rect 15304 16028 15332 16127
rect 23842 16124 23848 16176
rect 23900 16164 23906 16176
rect 24673 16167 24731 16173
rect 24673 16164 24685 16167
rect 23900 16136 24685 16164
rect 23900 16124 23906 16136
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 14139 16000 15332 16028
rect 15396 16068 15853 16096
rect 14139 15997 14151 16000
rect 14093 15991 14151 15997
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 8812 15932 9321 15960
rect 8812 15920 8818 15932
rect 9309 15929 9321 15932
rect 9355 15929 9367 15963
rect 9309 15923 9367 15929
rect 9953 15963 10011 15969
rect 9953 15929 9965 15963
rect 9999 15960 10011 15963
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 9999 15932 10793 15960
rect 9999 15929 10011 15932
rect 9953 15923 10011 15929
rect 10781 15929 10793 15932
rect 10827 15960 10839 15963
rect 10962 15960 10968 15972
rect 10827 15932 10968 15960
rect 10827 15929 10839 15932
rect 10781 15923 10839 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 13446 15960 13452 15972
rect 12943 15932 13452 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 13446 15920 13452 15932
rect 13504 15960 13510 15972
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 13504 15932 14197 15960
rect 13504 15920 13510 15932
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 15396 15960 15424 16068
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18414 16096 18420 16108
rect 18371 16068 18420 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18414 16056 18420 16068
rect 18472 16096 18478 16108
rect 19978 16096 19984 16108
rect 18472 16068 19984 16096
rect 18472 16056 18478 16068
rect 19978 16056 19984 16068
rect 20036 16096 20042 16108
rect 20438 16096 20444 16108
rect 20036 16068 20444 16096
rect 20036 16056 20042 16068
rect 20438 16056 20444 16068
rect 20496 16096 20502 16108
rect 24228 16105 24256 16136
rect 24673 16133 24685 16136
rect 24719 16133 24731 16167
rect 24673 16127 24731 16133
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 20496 16068 22017 16096
rect 20496 16056 20502 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16096 24271 16099
rect 24259 16068 24293 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 16028 18751 16031
rect 18966 16028 18972 16040
rect 18739 16000 18972 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 19444 16000 20269 16028
rect 14185 15923 14243 15929
rect 14752 15932 15424 15960
rect 14752 15904 14780 15932
rect 19444 15904 19472 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 20349 15963 20407 15969
rect 20349 15960 20361 15963
rect 19720 15932 20361 15960
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1581 15895 1639 15901
rect 1581 15892 1593 15895
rect 1452 15864 1593 15892
rect 1452 15852 1458 15864
rect 1581 15861 1593 15864
rect 1627 15861 1639 15895
rect 1581 15855 1639 15861
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2317 15895 2375 15901
rect 2317 15892 2329 15895
rect 1820 15864 2329 15892
rect 1820 15852 1826 15864
rect 2317 15861 2329 15864
rect 2363 15892 2375 15895
rect 2590 15892 2596 15904
rect 2363 15864 2596 15892
rect 2363 15861 2375 15864
rect 2317 15855 2375 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 3050 15892 3056 15904
rect 3011 15864 3056 15892
rect 3050 15852 3056 15864
rect 3108 15892 3114 15904
rect 3513 15895 3571 15901
rect 3513 15892 3525 15895
rect 3108 15864 3525 15892
rect 3108 15852 3114 15864
rect 3513 15861 3525 15864
rect 3559 15861 3571 15895
rect 4890 15892 4896 15904
rect 4851 15864 4896 15892
rect 3513 15855 3571 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 7282 15892 7288 15904
rect 7243 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7558 15852 7564 15904
rect 7616 15892 7622 15904
rect 7653 15895 7711 15901
rect 7653 15892 7665 15895
rect 7616 15864 7665 15892
rect 7616 15852 7622 15864
rect 7653 15861 7665 15864
rect 7699 15861 7711 15895
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 7653 15855 7711 15861
rect 10318 15852 10324 15864
rect 10376 15892 10382 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10376 15864 10885 15892
rect 10376 15852 10382 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 14734 15892 14740 15904
rect 14695 15864 14740 15892
rect 10873 15855 10931 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 15654 15892 15660 15904
rect 15252 15864 15660 15892
rect 15252 15852 15258 15864
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 19426 15892 19432 15904
rect 15804 15864 15849 15892
rect 19387 15864 19432 15892
rect 15804 15852 15810 15864
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 19720 15901 19748 15932
rect 20349 15929 20361 15932
rect 20395 15929 20407 15963
rect 21913 15963 21971 15969
rect 21913 15960 21925 15963
rect 20349 15923 20407 15929
rect 21284 15932 21925 15960
rect 19705 15895 19763 15901
rect 19705 15892 19717 15895
rect 19668 15864 19717 15892
rect 19668 15852 19674 15864
rect 19705 15861 19717 15864
rect 19751 15861 19763 15895
rect 19705 15855 19763 15861
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21284 15901 21312 15932
rect 21913 15929 21925 15932
rect 21959 15929 21971 15963
rect 21913 15923 21971 15929
rect 23477 15963 23535 15969
rect 23477 15929 23489 15963
rect 23523 15960 23535 15963
rect 23934 15960 23940 15972
rect 23523 15932 23940 15960
rect 23523 15929 23535 15932
rect 23477 15923 23535 15929
rect 23934 15920 23940 15932
rect 23992 15960 23998 15972
rect 24029 15963 24087 15969
rect 24029 15960 24041 15963
rect 23992 15932 24041 15960
rect 23992 15920 23998 15932
rect 24029 15929 24041 15932
rect 24075 15929 24087 15963
rect 24029 15923 24087 15929
rect 21269 15895 21327 15901
rect 21269 15892 21281 15895
rect 20864 15864 21281 15892
rect 20864 15852 20870 15864
rect 21269 15861 21281 15864
rect 21315 15861 21327 15895
rect 21269 15855 21327 15861
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 21784 15864 21833 15892
rect 21784 15852 21790 15864
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 24118 15892 24124 15904
rect 24079 15864 24124 15892
rect 21821 15855 21879 15861
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4890 15688 4896 15700
rect 4111 15660 4896 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 6178 15688 6184 15700
rect 6139 15660 6184 15688
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 8754 15688 8760 15700
rect 7340 15660 8760 15688
rect 7340 15648 7346 15660
rect 8754 15648 8760 15660
rect 8812 15688 8818 15700
rect 8849 15691 8907 15697
rect 8849 15688 8861 15691
rect 8812 15660 8861 15688
rect 8812 15648 8818 15660
rect 8849 15657 8861 15660
rect 8895 15657 8907 15691
rect 8849 15651 8907 15657
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 8996 15660 9689 15688
rect 8996 15648 9002 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 9677 15651 9735 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10928 15660 11069 15688
rect 10928 15648 10934 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15688 13231 15691
rect 13538 15688 13544 15700
rect 13219 15660 13544 15688
rect 13219 15657 13231 15660
rect 13173 15651 13231 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15565 15691 15623 15697
rect 15565 15688 15577 15691
rect 15252 15660 15577 15688
rect 15252 15648 15258 15660
rect 15565 15657 15577 15660
rect 15611 15688 15623 15691
rect 15746 15688 15752 15700
rect 15611 15660 15752 15688
rect 15611 15657 15623 15660
rect 15565 15651 15623 15657
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 19576 15660 19625 15688
rect 19576 15648 19582 15660
rect 19613 15657 19625 15660
rect 19659 15657 19671 15691
rect 19613 15651 19671 15657
rect 22925 15691 22983 15697
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 24118 15688 24124 15700
rect 22971 15660 24124 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 24118 15648 24124 15660
rect 24176 15688 24182 15700
rect 24305 15691 24363 15697
rect 24305 15688 24317 15691
rect 24176 15660 24317 15688
rect 24176 15648 24182 15660
rect 24305 15657 24317 15660
rect 24351 15657 24363 15691
rect 24305 15651 24363 15657
rect 4154 15580 4160 15632
rect 4212 15620 4218 15632
rect 4430 15620 4436 15632
rect 4212 15592 4436 15620
rect 4212 15580 4218 15592
rect 4430 15580 4436 15592
rect 4488 15580 4494 15632
rect 6917 15623 6975 15629
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 7374 15620 7380 15632
rect 6963 15592 7380 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 7374 15580 7380 15592
rect 7432 15580 7438 15632
rect 7745 15623 7803 15629
rect 7745 15589 7757 15623
rect 7791 15620 7803 15623
rect 7926 15620 7932 15632
rect 7791 15592 7932 15620
rect 7791 15589 7803 15592
rect 7745 15583 7803 15589
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 16758 15580 16764 15632
rect 16816 15620 16822 15632
rect 16936 15623 16994 15629
rect 16936 15620 16948 15623
rect 16816 15592 16948 15620
rect 16816 15580 16822 15592
rect 16936 15589 16948 15592
rect 16982 15620 16994 15623
rect 17494 15620 17500 15632
rect 16982 15592 17500 15620
rect 16982 15589 16994 15592
rect 16936 15583 16994 15589
rect 17494 15580 17500 15592
rect 17552 15580 17558 15632
rect 23842 15580 23848 15632
rect 23900 15620 23906 15632
rect 23937 15623 23995 15629
rect 23937 15620 23949 15623
rect 23900 15592 23949 15620
rect 23900 15580 23906 15592
rect 23937 15589 23949 15592
rect 23983 15589 23995 15623
rect 23937 15583 23995 15589
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1486 15552 1492 15564
rect 1443 15524 1492 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 1670 15561 1676 15564
rect 1664 15515 1676 15561
rect 1728 15552 1734 15564
rect 1728 15524 1764 15552
rect 1670 15512 1676 15515
rect 1728 15512 1734 15524
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9824 15524 10057 15552
rect 9824 15512 9830 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 13998 15552 14004 15564
rect 13959 15524 14004 15552
rect 10045 15515 10103 15521
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 16666 15552 16672 15564
rect 16627 15524 16672 15552
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 20714 15552 20720 15564
rect 20675 15524 20720 15552
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 23293 15555 23351 15561
rect 23293 15552 23305 15555
rect 23256 15524 23305 15552
rect 23256 15512 23262 15524
rect 23293 15521 23305 15524
rect 23339 15521 23351 15555
rect 23293 15515 23351 15521
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 26881 15555 26939 15561
rect 26881 15552 26893 15555
rect 26844 15524 26893 15552
rect 26844 15512 26850 15524
rect 26881 15521 26893 15524
rect 26927 15521 26939 15555
rect 26881 15515 26939 15521
rect 4522 15484 4528 15496
rect 4483 15456 4528 15484
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 4798 15484 4804 15496
rect 4755 15456 4804 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 3421 15419 3479 15425
rect 3421 15416 3433 15419
rect 2823 15388 3433 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 3421 15385 3433 15388
rect 3467 15416 3479 15419
rect 3694 15416 3700 15428
rect 3467 15388 3700 15416
rect 3467 15385 3479 15388
rect 3421 15379 3479 15385
rect 3694 15376 3700 15388
rect 3752 15416 3758 15428
rect 4724 15416 4752 15447
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 6270 15484 6276 15496
rect 6231 15456 6276 15484
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 10134 15484 10140 15496
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10284 15456 10329 15484
rect 10284 15444 10290 15456
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13320 15456 14105 15484
rect 13320 15444 13326 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14458 15484 14464 15496
rect 14323 15456 14464 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23566 15484 23572 15496
rect 23523 15456 23572 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 3752 15388 4752 15416
rect 3752 15376 3758 15388
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 23400 15416 23428 15447
rect 23348 15388 23428 15416
rect 23348 15376 23354 15388
rect 5810 15348 5816 15360
rect 5771 15320 5816 15348
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 7377 15351 7435 15357
rect 7377 15317 7389 15351
rect 7423 15348 7435 15351
rect 7558 15348 7564 15360
rect 7423 15320 7564 15348
rect 7423 15317 7435 15320
rect 7377 15311 7435 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 13538 15348 13544 15360
rect 13499 15320 13544 15348
rect 13538 15308 13544 15320
rect 13596 15308 13602 15360
rect 13633 15351 13691 15357
rect 13633 15317 13645 15351
rect 13679 15348 13691 15351
rect 13722 15348 13728 15360
rect 13679 15320 13728 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15348 18107 15351
rect 18230 15348 18236 15360
rect 18095 15320 18236 15348
rect 18095 15317 18107 15320
rect 18049 15311 18107 15317
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 19058 15348 19064 15360
rect 19019 15320 19064 15348
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20162 15308 20168 15360
rect 20220 15348 20226 15360
rect 20533 15351 20591 15357
rect 20533 15348 20545 15351
rect 20220 15320 20545 15348
rect 20220 15308 20226 15320
rect 20533 15317 20545 15320
rect 20579 15317 20591 15351
rect 20533 15311 20591 15317
rect 21545 15351 21603 15357
rect 21545 15317 21557 15351
rect 21591 15348 21603 15351
rect 21726 15348 21732 15360
rect 21591 15320 21732 15348
rect 21591 15317 21603 15320
rect 21545 15311 21603 15317
rect 21726 15308 21732 15320
rect 21784 15308 21790 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 23492 15348 23520 15447
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 26970 15484 26976 15496
rect 26931 15456 26976 15484
rect 26970 15444 26976 15456
rect 27028 15444 27034 15496
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27338 15484 27344 15496
rect 27203 15456 27344 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 27338 15444 27344 15456
rect 27396 15444 27402 15496
rect 22704 15320 23520 15348
rect 22704 15308 22710 15320
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 26053 15351 26111 15357
rect 26053 15348 26065 15351
rect 25740 15320 26065 15348
rect 25740 15308 25746 15320
rect 26053 15317 26065 15320
rect 26099 15317 26111 15351
rect 26053 15311 26111 15317
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 26513 15351 26571 15357
rect 26513 15348 26525 15351
rect 26384 15320 26525 15348
rect 26384 15308 26390 15320
rect 26513 15317 26525 15320
rect 26559 15317 26571 15351
rect 26513 15311 26571 15317
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1728 15116 1777 15144
rect 1728 15104 1734 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 2682 15144 2688 15156
rect 2643 15116 2688 15144
rect 1765 15107 1823 15113
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15144 4215 15147
rect 4430 15144 4436 15156
rect 4203 15116 4436 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 4798 15144 4804 15156
rect 4580 15116 4625 15144
rect 4759 15116 4804 15144
rect 4580 15104 4586 15116
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15144 5871 15147
rect 6362 15144 6368 15156
rect 5859 15116 6368 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10284 15116 10425 15144
rect 10284 15104 10290 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 13078 15144 13084 15156
rect 13039 15116 13084 15144
rect 10413 15107 10471 15113
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 13541 15147 13599 15153
rect 13541 15144 13553 15147
rect 13504 15116 13553 15144
rect 13504 15104 13510 15116
rect 13541 15113 13553 15116
rect 13587 15113 13599 15147
rect 15102 15144 15108 15156
rect 15063 15116 15108 15144
rect 13541 15107 13599 15113
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 16758 15144 16764 15156
rect 16719 15116 16764 15144
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 19024 15116 19073 15144
rect 19024 15104 19030 15116
rect 19061 15113 19073 15116
rect 19107 15144 19119 15147
rect 20714 15144 20720 15156
rect 19107 15116 20720 15144
rect 19107 15113 19119 15116
rect 19061 15107 19119 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 12713 15079 12771 15085
rect 12713 15045 12725 15079
rect 12759 15076 12771 15079
rect 14734 15076 14740 15088
rect 12759 15048 14740 15076
rect 12759 15045 12771 15048
rect 12713 15039 12771 15045
rect 3234 15008 3240 15020
rect 3195 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 15008 5595 15011
rect 6822 15008 6828 15020
rect 5583 14980 6828 15008
rect 5583 14977 5595 14980
rect 5537 14971 5595 14977
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 14108 15017 14136 15048
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 16724 15048 17049 15076
rect 16724 15036 16730 15048
rect 17037 15045 17049 15048
rect 17083 15076 17095 15079
rect 17954 15076 17960 15088
rect 17083 15048 17960 15076
rect 17083 15045 17095 15048
rect 17037 15039 17095 15045
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 19613 15079 19671 15085
rect 19613 15045 19625 15079
rect 19659 15076 19671 15079
rect 19702 15076 19708 15088
rect 19659 15048 19708 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 19702 15036 19708 15048
rect 19760 15036 19766 15088
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13596 14980 14013 15008
rect 13596 14968 13602 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 14977 14151 15011
rect 15654 15008 15660 15020
rect 15615 14980 15660 15008
rect 14093 14971 14151 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 20036 14980 20177 15008
rect 20036 14968 20042 14980
rect 20165 14977 20177 14980
rect 20211 14977 20223 15011
rect 24302 15008 24308 15020
rect 24263 14980 24308 15008
rect 20165 14971 20223 14977
rect 24302 14968 24308 14980
rect 24360 15008 24366 15020
rect 25133 15011 25191 15017
rect 24360 14980 24900 15008
rect 24360 14968 24366 14980
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 2792 14912 3065 14940
rect 2225 14875 2283 14881
rect 2225 14841 2237 14875
rect 2271 14872 2283 14875
rect 2792 14872 2820 14912
rect 3053 14909 3065 14912
rect 3099 14940 3111 14943
rect 4062 14940 4068 14952
rect 3099 14912 4068 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 14550 14900 14556 14952
rect 14608 14940 14614 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14608 14912 14657 14940
rect 14608 14900 14614 14912
rect 14645 14909 14657 14912
rect 14691 14940 14703 14943
rect 15470 14940 15476 14952
rect 14691 14912 15476 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 19058 14900 19064 14952
rect 19116 14940 19122 14952
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 19116 14912 19257 14940
rect 19116 14900 19122 14912
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 20070 14940 20076 14952
rect 19576 14912 20076 14940
rect 19576 14900 19582 14912
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14940 23075 14943
rect 23290 14940 23296 14952
rect 23063 14912 23296 14940
rect 23063 14909 23075 14912
rect 23017 14903 23075 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 24872 14949 24900 14980
rect 25133 14977 25145 15011
rect 25179 15008 25191 15011
rect 25222 15008 25228 15020
rect 25179 14980 25228 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 24857 14943 24915 14949
rect 24857 14909 24869 14943
rect 24903 14909 24915 14943
rect 24857 14903 24915 14909
rect 25774 14900 25780 14952
rect 25832 14940 25838 14952
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25832 14912 25881 14940
rect 25832 14900 25838 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 26050 14940 26056 14952
rect 26011 14912 26056 14940
rect 25869 14903 25927 14909
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 2271 14844 2820 14872
rect 2884 14844 3157 14872
rect 2271 14841 2283 14844
rect 2225 14835 2283 14841
rect 2593 14807 2651 14813
rect 2593 14773 2605 14807
rect 2639 14804 2651 14807
rect 2774 14804 2780 14816
rect 2639 14776 2780 14804
rect 2639 14773 2651 14776
rect 2593 14767 2651 14773
rect 2774 14764 2780 14776
rect 2832 14804 2838 14816
rect 2884 14804 2912 14844
rect 3145 14841 3157 14844
rect 3191 14841 3203 14875
rect 3145 14835 3203 14841
rect 6454 14832 6460 14884
rect 6512 14872 6518 14884
rect 7098 14881 7104 14884
rect 6641 14875 6699 14881
rect 6641 14872 6653 14875
rect 6512 14844 6653 14872
rect 6512 14832 6518 14844
rect 6641 14841 6653 14844
rect 6687 14872 6699 14875
rect 7092 14872 7104 14881
rect 6687 14844 7104 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7092 14835 7104 14844
rect 7098 14832 7104 14835
rect 7156 14832 7162 14884
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 13722 14872 13728 14884
rect 13228 14844 13728 14872
rect 13228 14832 13234 14844
rect 13722 14832 13728 14844
rect 13780 14872 13786 14884
rect 13909 14875 13967 14881
rect 13909 14872 13921 14875
rect 13780 14844 13921 14872
rect 13780 14832 13786 14844
rect 13909 14841 13921 14844
rect 13955 14841 13967 14875
rect 14918 14872 14924 14884
rect 14879 14844 14924 14872
rect 13909 14835 13967 14841
rect 14918 14832 14924 14844
rect 14976 14872 14982 14884
rect 15378 14872 15384 14884
rect 14976 14844 15384 14872
rect 14976 14832 14982 14844
rect 15378 14832 15384 14844
rect 15436 14872 15442 14884
rect 15565 14875 15623 14881
rect 15565 14872 15577 14875
rect 15436 14844 15577 14872
rect 15436 14832 15442 14844
rect 15565 14841 15577 14844
rect 15611 14841 15623 14875
rect 15565 14835 15623 14841
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14872 19027 14875
rect 19886 14872 19892 14884
rect 19015 14844 19892 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 19886 14832 19892 14844
rect 19944 14872 19950 14884
rect 19981 14875 20039 14881
rect 19981 14872 19993 14875
rect 19944 14844 19993 14872
rect 19944 14832 19950 14844
rect 19981 14841 19993 14844
rect 20027 14872 20039 14875
rect 20254 14872 20260 14884
rect 20027 14844 20260 14872
rect 20027 14841 20039 14844
rect 19981 14835 20039 14841
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 24029 14875 24087 14881
rect 24029 14841 24041 14875
rect 24075 14872 24087 14875
rect 24949 14875 25007 14881
rect 24949 14872 24961 14875
rect 24075 14844 24961 14872
rect 24075 14841 24087 14844
rect 24029 14835 24087 14841
rect 24949 14841 24961 14844
rect 24995 14872 25007 14875
rect 26142 14872 26148 14884
rect 24995 14844 26148 14872
rect 24995 14841 25007 14844
rect 24949 14835 25007 14841
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 26326 14881 26332 14884
rect 26320 14872 26332 14881
rect 26287 14844 26332 14872
rect 26320 14835 26332 14844
rect 26326 14832 26332 14835
rect 26384 14832 26390 14884
rect 3694 14804 3700 14816
rect 2832 14776 2925 14804
rect 3655 14776 3700 14804
rect 2832 14764 2838 14776
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 6270 14804 6276 14816
rect 6231 14776 6276 14804
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 9766 14804 9772 14816
rect 9727 14776 9772 14804
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 10134 14804 10140 14816
rect 10095 14776 10140 14804
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 23198 14764 23204 14816
rect 23256 14804 23262 14816
rect 23293 14807 23351 14813
rect 23293 14804 23305 14807
rect 23256 14776 23305 14804
rect 23256 14764 23262 14776
rect 23293 14773 23305 14776
rect 23339 14773 23351 14807
rect 24486 14804 24492 14816
rect 24447 14776 24492 14804
rect 23293 14767 23351 14773
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 27430 14804 27436 14816
rect 27391 14776 27436 14804
rect 27430 14764 27436 14776
rect 27488 14764 27494 14816
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1486 14560 1492 14612
rect 1544 14560 1550 14612
rect 1670 14560 1676 14612
rect 1728 14600 1734 14612
rect 2777 14603 2835 14609
rect 2777 14600 2789 14603
rect 1728 14572 2789 14600
rect 1728 14560 1734 14572
rect 2777 14569 2789 14572
rect 2823 14600 2835 14603
rect 3234 14600 3240 14612
rect 2823 14572 3240 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5868 14572 6009 14600
rect 5868 14560 5874 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14569 7159 14603
rect 9214 14600 9220 14612
rect 9175 14572 9220 14600
rect 7101 14563 7159 14569
rect 1504 14532 1532 14560
rect 3694 14532 3700 14544
rect 1412 14504 3700 14532
rect 1412 14473 1440 14504
rect 3252 14476 3280 14504
rect 3694 14492 3700 14504
rect 3752 14492 3758 14544
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 5905 14535 5963 14541
rect 5905 14532 5917 14535
rect 5684 14504 5917 14532
rect 5684 14492 5690 14504
rect 5905 14501 5917 14504
rect 5951 14532 5963 14535
rect 7116 14532 7144 14563
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13596 14572 13645 14600
rect 13596 14560 13602 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13633 14563 13691 14569
rect 26145 14603 26203 14609
rect 26145 14569 26157 14603
rect 26191 14600 26203 14603
rect 26326 14600 26332 14612
rect 26191 14572 26332 14600
rect 26191 14569 26203 14572
rect 26145 14563 26203 14569
rect 26326 14560 26332 14572
rect 26384 14600 26390 14612
rect 27157 14603 27215 14609
rect 27157 14600 27169 14603
rect 26384 14572 27169 14600
rect 26384 14560 26390 14572
rect 27157 14569 27169 14572
rect 27203 14600 27215 14603
rect 27338 14600 27344 14612
rect 27203 14572 27344 14600
rect 27203 14569 27215 14572
rect 27157 14563 27215 14569
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 9232 14532 9260 14560
rect 10226 14532 10232 14544
rect 5951 14504 7144 14532
rect 7300 14504 7788 14532
rect 9232 14504 10232 14532
rect 5951 14501 5963 14504
rect 5905 14495 5963 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14433 1455 14467
rect 1397 14427 1455 14433
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 1653 14467 1711 14473
rect 1653 14464 1665 14467
rect 1544 14436 1665 14464
rect 1544 14424 1550 14436
rect 1653 14433 1665 14436
rect 1699 14433 1711 14467
rect 1653 14427 1711 14433
rect 3234 14424 3240 14476
rect 3292 14424 3298 14476
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14464 6975 14467
rect 7098 14464 7104 14476
rect 6963 14436 7104 14464
rect 6963 14433 6975 14436
rect 6917 14427 6975 14433
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 7300 14464 7328 14504
rect 7466 14464 7472 14476
rect 7156 14436 7328 14464
rect 7427 14436 7472 14464
rect 7156 14424 7162 14436
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6196 14328 6224 14359
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7760 14405 7788 14504
rect 10226 14492 10232 14504
rect 10284 14532 10290 14544
rect 10772 14535 10830 14541
rect 10284 14504 10548 14532
rect 10284 14492 10290 14504
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 10520 14473 10548 14504
rect 10772 14501 10784 14535
rect 10818 14532 10830 14535
rect 10870 14532 10876 14544
rect 10818 14504 10876 14532
rect 10818 14501 10830 14504
rect 10772 14495 10830 14501
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 14001 14535 14059 14541
rect 14001 14501 14013 14535
rect 14047 14532 14059 14535
rect 14090 14532 14096 14544
rect 14047 14504 14096 14532
rect 14047 14501 14059 14504
rect 14001 14495 14059 14501
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 8168 14436 9413 14464
rect 8168 14424 8174 14436
rect 9401 14433 9413 14436
rect 9447 14464 9459 14467
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9447 14436 9873 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 9861 14433 9873 14436
rect 9907 14433 9919 14467
rect 9861 14427 9919 14433
rect 10505 14467 10563 14473
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 11698 14464 11704 14476
rect 10551 14436 11704 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14458 14464 14464 14476
rect 13587 14436 14464 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7248 14368 7573 14396
rect 7248 14356 7254 14368
rect 7561 14365 7573 14368
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 9030 14396 9036 14408
rect 7791 14368 9036 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 9030 14356 9036 14368
rect 9088 14356 9094 14408
rect 14292 14405 14320 14436
rect 14458 14424 14464 14436
rect 14516 14464 14522 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14516 14436 15485 14464
rect 14516 14424 14522 14436
rect 15473 14433 15485 14436
rect 15519 14464 15531 14467
rect 15654 14464 15660 14476
rect 15519 14436 15660 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16390 14464 16396 14476
rect 16351 14436 16396 14464
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 17954 14464 17960 14476
rect 17915 14436 17960 14464
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18230 14473 18236 14476
rect 18224 14464 18236 14473
rect 18191 14436 18236 14464
rect 18224 14427 18236 14436
rect 18230 14424 18236 14427
rect 18288 14424 18294 14476
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 22824 14467 22882 14473
rect 22824 14464 22836 14467
rect 22704 14436 22836 14464
rect 22704 14424 22710 14436
rect 22824 14433 22836 14436
rect 22870 14464 22882 14467
rect 22870 14436 24624 14464
rect 22870 14433 22882 14436
rect 22824 14427 22882 14433
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 14323 14368 14357 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 6270 14328 6276 14340
rect 6183 14300 6276 14328
rect 6270 14288 6276 14300
rect 6328 14328 6334 14340
rect 8202 14328 8208 14340
rect 6328 14300 8208 14328
rect 6328 14288 6334 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 7926 14220 7932 14272
rect 7984 14260 7990 14272
rect 8113 14263 8171 14269
rect 8113 14260 8125 14263
rect 7984 14232 8125 14260
rect 7984 14220 7990 14232
rect 8113 14229 8125 14232
rect 8159 14229 8171 14263
rect 11882 14260 11888 14272
rect 11843 14232 11888 14260
rect 8113 14223 8171 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 14108 14260 14136 14359
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 15896 14368 16497 14396
rect 15896 14356 15902 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 22554 14396 22560 14408
rect 22515 14368 22560 14396
rect 16577 14359 16635 14365
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 16592 14328 16620 14359
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 15620 14300 16620 14328
rect 15620 14288 15626 14300
rect 16500 14272 16528 14300
rect 14182 14260 14188 14272
rect 14108 14232 14188 14260
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16390 14260 16396 14272
rect 16071 14232 16396 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 19334 14260 19340 14272
rect 19295 14232 19340 14260
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19978 14260 19984 14272
rect 19939 14232 19984 14260
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 23937 14263 23995 14269
rect 23937 14229 23949 14263
rect 23983 14260 23995 14263
rect 24026 14260 24032 14272
rect 23983 14232 24032 14260
rect 23983 14229 23995 14232
rect 23937 14223 23995 14229
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 24596 14269 24624 14436
rect 24581 14263 24639 14269
rect 24581 14229 24593 14263
rect 24627 14260 24639 14263
rect 25222 14260 25228 14272
rect 24627 14232 25228 14260
rect 24627 14229 24639 14232
rect 24581 14223 24639 14229
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 26786 14260 26792 14272
rect 26747 14232 26792 14260
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1544 14028 1593 14056
rect 1544 14016 1550 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1949 14059 2007 14065
rect 1949 14056 1961 14059
rect 1728 14028 1961 14056
rect 1728 14016 1734 14028
rect 1949 14025 1961 14028
rect 1995 14025 2007 14059
rect 4430 14056 4436 14068
rect 4391 14028 4436 14056
rect 1949 14019 2007 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5261 14059 5319 14065
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 5810 14056 5816 14068
rect 5307 14028 5816 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 7098 14056 7104 14068
rect 6687 14028 7104 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 10502 14056 10508 14068
rect 10463 14028 10508 14056
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11698 14056 11704 14068
rect 11659 14028 11704 14056
rect 11698 14016 11704 14028
rect 11756 14056 11762 14068
rect 12434 14056 12440 14068
rect 11756 14028 12440 14056
rect 11756 14016 11762 14028
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18601 14059 18659 14065
rect 18601 14056 18613 14059
rect 18012 14028 18613 14056
rect 18012 14016 18018 14028
rect 18601 14025 18613 14028
rect 18647 14025 18659 14059
rect 18601 14019 18659 14025
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 20036 14028 21557 14056
rect 20036 14016 20042 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 22646 14056 22652 14068
rect 22607 14028 22652 14056
rect 21545 14019 21603 14025
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 25222 14016 25228 14068
rect 25280 14056 25286 14068
rect 25280 14028 25820 14056
rect 25280 14016 25286 14028
rect 5629 13991 5687 13997
rect 5629 13957 5641 13991
rect 5675 13988 5687 13991
rect 6270 13988 6276 14000
rect 5675 13960 6276 13988
rect 5675 13957 5687 13960
rect 5629 13951 5687 13957
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3007 13892 3188 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13821 3111 13855
rect 3160 13852 3188 13892
rect 3320 13855 3378 13861
rect 3320 13852 3332 13855
rect 3160 13824 3332 13852
rect 3053 13815 3111 13821
rect 3320 13821 3332 13824
rect 3366 13852 3378 13855
rect 5644 13852 5672 13951
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 7469 13991 7527 13997
rect 7469 13988 7481 13991
rect 6880 13960 7481 13988
rect 6880 13948 6886 13960
rect 7469 13957 7481 13960
rect 7515 13957 7527 13991
rect 9125 13991 9183 13997
rect 9125 13988 9137 13991
rect 7469 13951 7527 13957
rect 7944 13960 9137 13988
rect 7944 13932 7972 13960
rect 9125 13957 9137 13960
rect 9171 13957 9183 13991
rect 10689 13991 10747 13997
rect 10689 13988 10701 13991
rect 9125 13951 9183 13957
rect 9600 13960 10701 13988
rect 7926 13920 7932 13932
rect 7887 13892 7932 13920
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8202 13920 8208 13932
rect 8159 13892 8208 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9600 13929 9628 13960
rect 10689 13957 10701 13960
rect 10735 13957 10747 13991
rect 11882 13988 11888 14000
rect 10689 13951 10747 13957
rect 10796 13960 11888 13988
rect 9585 13923 9643 13929
rect 9585 13920 9597 13923
rect 9272 13892 9597 13920
rect 9272 13880 9278 13892
rect 9585 13889 9597 13892
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10796 13920 10824 13960
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 16025 13991 16083 13997
rect 16025 13988 16037 13991
rect 15252 13960 16037 13988
rect 15252 13948 15258 13960
rect 16025 13957 16037 13960
rect 16071 13957 16083 13991
rect 16025 13951 16083 13957
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 24026 13988 24032 14000
rect 23532 13960 24032 13988
rect 23532 13948 23538 13960
rect 24026 13948 24032 13960
rect 24084 13988 24090 14000
rect 25792 13997 25820 14028
rect 24581 13991 24639 13997
rect 24581 13988 24593 13991
rect 24084 13960 24593 13988
rect 24084 13948 24090 13960
rect 24581 13957 24593 13960
rect 24627 13988 24639 13991
rect 25777 13991 25835 13997
rect 24627 13960 25268 13988
rect 24627 13957 24639 13960
rect 24581 13951 24639 13957
rect 25240 13932 25268 13960
rect 25777 13957 25789 13991
rect 25823 13988 25835 13991
rect 25823 13960 26924 13988
rect 25823 13957 25835 13960
rect 25777 13951 25835 13957
rect 9815 13892 10824 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 3366 13824 5672 13852
rect 6273 13855 6331 13861
rect 3366 13821 3378 13824
rect 3320 13815 3378 13821
rect 6273 13821 6285 13855
rect 6319 13852 6331 13855
rect 7190 13852 7196 13864
rect 6319 13824 6868 13852
rect 7151 13824 7196 13852
rect 6319 13821 6331 13824
rect 6273 13815 6331 13821
rect 3068 13784 3096 13815
rect 3234 13784 3240 13796
rect 3068 13756 3240 13784
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 5721 13787 5779 13793
rect 5721 13753 5733 13787
rect 5767 13784 5779 13787
rect 6840 13784 6868 13824
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 9030 13852 9036 13864
rect 8943 13824 9036 13852
rect 9030 13812 9036 13824
rect 9088 13852 9094 13864
rect 9784 13852 9812 13883
rect 10870 13880 10876 13932
rect 10928 13920 10934 13932
rect 11241 13923 11299 13929
rect 11241 13920 11253 13923
rect 10928 13892 11253 13920
rect 10928 13880 10934 13892
rect 11241 13889 11253 13892
rect 11287 13889 11299 13923
rect 11241 13883 11299 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 14182 13920 14188 13932
rect 13771 13892 14188 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 16264 13892 16589 13920
rect 16264 13880 16270 13892
rect 16577 13889 16589 13892
rect 16623 13889 16635 13923
rect 16577 13883 16635 13889
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20119 13892 20300 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 9088 13824 9812 13852
rect 9088 13812 9094 13824
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10502 13852 10508 13864
rect 10284 13824 10508 13852
rect 10284 13812 10290 13824
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 10652 13824 11161 13852
rect 10652 13812 10658 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 14090 13852 14096 13864
rect 14051 13824 14096 13852
rect 11149 13815 11207 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13852 15255 13855
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 15243 13824 16497 13852
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 16485 13815 16543 13821
rect 16868 13824 17141 13852
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 5767 13756 6776 13784
rect 6840 13756 7849 13784
rect 5767 13753 5779 13756
rect 5721 13747 5779 13753
rect 6748 13716 6776 13756
rect 7837 13753 7849 13756
rect 7883 13784 7895 13787
rect 8018 13784 8024 13796
rect 7883 13756 8024 13784
rect 7883 13753 7895 13756
rect 7837 13747 7895 13753
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 8665 13787 8723 13793
rect 8665 13753 8677 13787
rect 8711 13784 8723 13787
rect 9493 13787 9551 13793
rect 9493 13784 9505 13787
rect 8711 13756 9505 13784
rect 8711 13753 8723 13756
rect 8665 13747 8723 13753
rect 9493 13753 9505 13756
rect 9539 13784 9551 13787
rect 9766 13784 9772 13796
rect 9539 13756 9772 13784
rect 9539 13753 9551 13756
rect 9493 13747 9551 13753
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 10410 13744 10416 13796
rect 10468 13784 10474 13796
rect 11057 13787 11115 13793
rect 11057 13784 11069 13787
rect 10468 13756 11069 13784
rect 10468 13744 10474 13756
rect 11057 13753 11069 13756
rect 11103 13784 11115 13787
rect 11698 13784 11704 13796
rect 11103 13756 11704 13784
rect 11103 13753 11115 13756
rect 11057 13747 11115 13753
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 16500 13784 16528 13815
rect 16758 13784 16764 13796
rect 16500 13756 16764 13784
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 7466 13716 7472 13728
rect 6748 13688 7472 13716
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 10226 13716 10232 13728
rect 10187 13688 10232 13716
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 16393 13719 16451 13725
rect 16393 13685 16405 13719
rect 16439 13716 16451 13719
rect 16868 13716 16896 13824
rect 17129 13821 17141 13824
rect 17175 13852 17187 13855
rect 17862 13852 17868 13864
rect 17175 13824 17868 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20272 13852 20300 13892
rect 24486 13880 24492 13932
rect 24544 13920 24550 13932
rect 25222 13920 25228 13932
rect 24544 13892 24992 13920
rect 25183 13892 25228 13920
rect 24544 13880 24550 13892
rect 20438 13861 20444 13864
rect 20432 13852 20444 13861
rect 20272 13824 20444 13852
rect 20432 13815 20444 13824
rect 20438 13812 20444 13815
rect 20496 13812 20502 13864
rect 24213 13855 24271 13861
rect 24213 13821 24225 13855
rect 24259 13852 24271 13855
rect 24964 13852 24992 13892
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 26050 13920 26056 13932
rect 26011 13892 26056 13920
rect 26050 13880 26056 13892
rect 26108 13920 26114 13932
rect 26326 13920 26332 13932
rect 26108 13892 26332 13920
rect 26108 13880 26114 13892
rect 26326 13880 26332 13892
rect 26384 13880 26390 13932
rect 26896 13929 26924 13960
rect 26881 13923 26939 13929
rect 26881 13889 26893 13923
rect 26927 13920 26939 13923
rect 27430 13920 27436 13932
rect 26927 13892 27436 13920
rect 26927 13889 26939 13892
rect 26881 13883 26939 13889
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 25133 13855 25191 13861
rect 25133 13852 25145 13855
rect 24259 13824 24900 13852
rect 24964 13824 25145 13852
rect 24259 13821 24271 13824
rect 24213 13815 24271 13821
rect 24872 13784 24900 13824
rect 25133 13821 25145 13824
rect 25179 13821 25191 13855
rect 25133 13815 25191 13821
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26292 13824 26709 13852
rect 26292 13812 26298 13824
rect 26697 13821 26709 13824
rect 26743 13821 26755 13855
rect 26697 13815 26755 13821
rect 25041 13787 25099 13793
rect 25041 13784 25053 13787
rect 24872 13756 25053 13784
rect 25041 13753 25053 13756
rect 25087 13784 25099 13787
rect 25087 13756 26188 13784
rect 25087 13753 25099 13756
rect 25041 13747 25099 13753
rect 16439 13688 16896 13716
rect 16439 13685 16451 13688
rect 16393 13679 16451 13685
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 18230 13716 18236 13728
rect 17368 13688 18236 13716
rect 17368 13676 17374 13688
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 22554 13716 22560 13728
rect 22244 13688 22560 13716
rect 22244 13676 22250 13688
rect 22554 13676 22560 13688
rect 22612 13716 22618 13728
rect 22925 13719 22983 13725
rect 22925 13716 22937 13719
rect 22612 13688 22937 13716
rect 22612 13676 22618 13688
rect 22925 13685 22937 13688
rect 22971 13685 22983 13719
rect 24670 13716 24676 13728
rect 24631 13688 24676 13716
rect 22925 13679 22983 13685
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 26160 13716 26188 13756
rect 26326 13744 26332 13796
rect 26384 13784 26390 13796
rect 26605 13787 26663 13793
rect 26605 13784 26617 13787
rect 26384 13756 26617 13784
rect 26384 13744 26390 13756
rect 26605 13753 26617 13756
rect 26651 13784 26663 13787
rect 27154 13784 27160 13796
rect 26651 13756 27160 13784
rect 26651 13753 26663 13756
rect 26605 13747 26663 13753
rect 27154 13744 27160 13756
rect 27212 13744 27218 13796
rect 26237 13719 26295 13725
rect 26237 13716 26249 13719
rect 26160 13688 26249 13716
rect 26237 13685 26249 13688
rect 26283 13685 26295 13719
rect 26237 13679 26295 13685
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6270 13512 6276 13524
rect 6183 13484 6276 13512
rect 6270 13472 6276 13484
rect 6328 13512 6334 13524
rect 6822 13512 6828 13524
rect 6328 13484 6828 13512
rect 6328 13472 6334 13484
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7466 13512 7472 13524
rect 7239 13484 7472 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10468 13484 10701 13512
rect 10468 13472 10474 13484
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 10689 13475 10747 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 12492 13484 12541 13512
rect 12492 13472 12498 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16298 13512 16304 13524
rect 16163 13484 16304 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5592 13416 6193 13444
rect 5592 13404 5598 13416
rect 6181 13413 6193 13416
rect 6227 13444 6239 13447
rect 6546 13444 6552 13456
rect 6227 13416 6552 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 6546 13404 6552 13416
rect 6604 13404 6610 13456
rect 7929 13447 7987 13453
rect 7929 13413 7941 13447
rect 7975 13444 7987 13447
rect 8202 13444 8208 13456
rect 7975 13416 8208 13444
rect 7975 13413 7987 13416
rect 7929 13407 7987 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 8754 13404 8760 13456
rect 8812 13444 8818 13456
rect 10137 13447 10195 13453
rect 10137 13444 10149 13447
rect 8812 13416 10149 13444
rect 8812 13404 8818 13416
rect 10137 13413 10149 13416
rect 10183 13413 10195 13447
rect 10137 13407 10195 13413
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 8110 13376 8116 13388
rect 7607 13348 8116 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 10042 13376 10048 13388
rect 8904 13348 10048 13376
rect 8904 13336 8910 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 12544 13376 12572 13475
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16758 13512 16764 13524
rect 16719 13484 16764 13512
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 18325 13515 18383 13521
rect 18325 13512 18337 13515
rect 17920 13484 18337 13512
rect 17920 13472 17926 13484
rect 18325 13481 18337 13484
rect 18371 13481 18383 13515
rect 20162 13512 20168 13524
rect 20123 13484 20168 13512
rect 18325 13475 18383 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24673 13515 24731 13521
rect 24673 13512 24685 13515
rect 24544 13484 24685 13512
rect 24544 13472 24550 13484
rect 24673 13481 24685 13484
rect 24719 13481 24731 13515
rect 24673 13475 24731 13481
rect 25130 13472 25136 13524
rect 25188 13472 25194 13524
rect 26234 13512 26240 13524
rect 26195 13484 26240 13512
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16393 13447 16451 13453
rect 16393 13444 16405 13447
rect 16264 13416 16405 13444
rect 16264 13404 16270 13416
rect 16393 13413 16405 13416
rect 16439 13413 16451 13447
rect 17126 13444 17132 13456
rect 17087 13416 17132 13444
rect 16393 13407 16451 13413
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 22554 13404 22560 13456
rect 22612 13444 22618 13456
rect 22732 13447 22790 13453
rect 22732 13444 22744 13447
rect 22612 13416 22744 13444
rect 22612 13404 22618 13416
rect 22732 13413 22744 13416
rect 22778 13444 22790 13447
rect 23382 13444 23388 13456
rect 22778 13416 23388 13444
rect 22778 13413 22790 13416
rect 22732 13407 22790 13413
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12544 13348 12725 13376
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 12980 13379 13038 13385
rect 12980 13345 12992 13379
rect 13026 13376 13038 13379
rect 13354 13376 13360 13388
rect 13026 13348 13360 13376
rect 13026 13345 13038 13348
rect 12980 13339 13038 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 18690 13376 18696 13388
rect 18651 13348 18696 13376
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1854 13308 1860 13320
rect 1719 13280 1860 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1854 13268 1860 13280
rect 1912 13308 1918 13320
rect 3145 13311 3203 13317
rect 3145 13308 3157 13311
rect 1912 13280 3157 13308
rect 1912 13268 1918 13280
rect 3145 13277 3157 13280
rect 3191 13308 3203 13311
rect 3234 13308 3240 13320
rect 3191 13280 3240 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 6365 13311 6423 13317
rect 6365 13308 6377 13311
rect 5776 13280 6377 13308
rect 5776 13268 5782 13280
rect 6365 13277 6377 13280
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 9030 13308 9036 13320
rect 8711 13280 9036 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8496 13240 8524 13271
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10321 13311 10379 13317
rect 10321 13308 10333 13311
rect 10284 13280 10333 13308
rect 10284 13268 10290 13280
rect 10321 13277 10333 13280
rect 10367 13308 10379 13311
rect 10367 13280 10916 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 9677 13243 9735 13249
rect 9677 13240 9689 13243
rect 8260 13212 9689 13240
rect 8260 13200 8266 13212
rect 9677 13209 9689 13212
rect 9723 13209 9735 13243
rect 9677 13203 9735 13209
rect 10888 13184 10916 13280
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 17310 13308 17316 13320
rect 16632 13280 17316 13308
rect 16632 13268 16638 13280
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 18322 13268 18328 13320
rect 18380 13308 18386 13320
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18380 13280 18797 13308
rect 18380 13268 18386 13280
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18877 13311 18935 13317
rect 18877 13277 18889 13311
rect 18923 13277 18935 13311
rect 18877 13271 18935 13277
rect 18230 13200 18236 13252
rect 18288 13240 18294 13252
rect 18892 13240 18920 13271
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22244 13280 22477 13308
rect 22244 13268 22250 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 25148 13308 25176 13472
rect 26878 13376 26884 13388
rect 26839 13348 26884 13376
rect 26878 13336 26884 13348
rect 26936 13336 26942 13388
rect 25222 13308 25228 13320
rect 25148 13280 25228 13308
rect 22465 13271 22523 13277
rect 25222 13268 25228 13280
rect 25280 13268 25286 13320
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 26973 13311 27031 13317
rect 26973 13308 26985 13311
rect 26752 13280 26985 13308
rect 26752 13268 26758 13280
rect 26973 13277 26985 13280
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13308 27215 13311
rect 27430 13308 27436 13320
rect 27203 13280 27436 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 18966 13240 18972 13252
rect 18288 13212 18972 13240
rect 18288 13200 18294 13212
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 24854 13200 24860 13252
rect 24912 13240 24918 13252
rect 25682 13240 25688 13252
rect 24912 13212 25688 13240
rect 24912 13200 24918 13212
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 5810 13172 5816 13184
rect 5771 13144 5816 13172
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 10870 13132 10876 13184
rect 10928 13172 10934 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10928 13144 11069 13172
rect 10928 13132 10934 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 13964 13144 14105 13172
rect 13964 13132 13970 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14734 13172 14740 13184
rect 14695 13144 14740 13172
rect 14093 13135 14151 13141
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 23474 13132 23480 13184
rect 23532 13172 23538 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 23532 13144 23857 13172
rect 23532 13132 23538 13144
rect 23845 13141 23857 13144
rect 23891 13172 23903 13175
rect 24302 13172 24308 13184
rect 23891 13144 24308 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 26513 13175 26571 13181
rect 26513 13172 26525 13175
rect 26384 13144 26525 13172
rect 26384 13132 26390 13144
rect 26513 13141 26525 13144
rect 26559 13141 26571 13175
rect 26513 13135 26571 13141
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5776 12940 5825 12968
rect 5776 12928 5782 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 6270 12968 6276 12980
rect 6231 12940 6276 12968
rect 5813 12931 5871 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7377 12971 7435 12977
rect 7377 12937 7389 12971
rect 7423 12968 7435 12971
rect 8110 12968 8116 12980
rect 7423 12940 8116 12968
rect 7423 12937 7435 12940
rect 7377 12931 7435 12937
rect 8110 12928 8116 12940
rect 8168 12968 8174 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 8168 12940 8217 12968
rect 8168 12928 8174 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8812 12940 9229 12968
rect 8812 12928 8818 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9766 12968 9772 12980
rect 9727 12940 9772 12968
rect 9217 12931 9275 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 15102 12968 15108 12980
rect 13955 12940 15108 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15841 12971 15899 12977
rect 15841 12937 15853 12971
rect 15887 12968 15899 12971
rect 16482 12968 16488 12980
rect 15887 12940 16488 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 16224 12912 16252 12940
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17037 12971 17095 12977
rect 17037 12937 17049 12971
rect 17083 12968 17095 12971
rect 17218 12968 17224 12980
rect 17083 12940 17224 12968
rect 17083 12937 17095 12940
rect 17037 12931 17095 12937
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 19024 12940 19073 12968
rect 19024 12928 19030 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 22186 12968 22192 12980
rect 22147 12940 22192 12968
rect 19061 12931 19119 12937
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 22554 12968 22560 12980
rect 22515 12940 22560 12968
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 26878 12928 26884 12980
rect 26936 12968 26942 12980
rect 27065 12971 27123 12977
rect 27065 12968 27077 12971
rect 26936 12940 27077 12968
rect 26936 12928 26942 12940
rect 27065 12937 27077 12940
rect 27111 12968 27123 12971
rect 27111 12940 27292 12968
rect 27111 12937 27123 12940
rect 27065 12931 27123 12937
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 9030 12900 9036 12912
rect 7791 12872 9036 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 15933 12903 15991 12909
rect 15933 12900 15945 12903
rect 14792 12872 15945 12900
rect 14792 12860 14798 12872
rect 15933 12869 15945 12872
rect 15979 12869 15991 12903
rect 15933 12863 15991 12869
rect 16206 12860 16212 12912
rect 16264 12860 16270 12912
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 16356 12872 16528 12900
rect 16356 12860 16362 12872
rect 16500 12844 16528 12872
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17313 12903 17371 12909
rect 17313 12900 17325 12903
rect 17184 12872 17325 12900
rect 17184 12860 17190 12872
rect 17313 12869 17325 12872
rect 17359 12869 17371 12903
rect 24670 12900 24676 12912
rect 17313 12863 17371 12869
rect 24228 12872 24676 12900
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12832 4215 12835
rect 5166 12832 5172 12844
rect 4203 12804 5172 12832
rect 4203 12801 4215 12804
rect 4157 12795 4215 12801
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12832 8171 12835
rect 8294 12832 8300 12844
rect 8159 12804 8300 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9858 12832 9864 12844
rect 9723 12804 9864 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 9858 12792 9864 12804
rect 9916 12832 9922 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9916 12804 10241 12832
rect 9916 12792 9922 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10870 12832 10876 12844
rect 10459 12804 10876 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 13354 12832 13360 12844
rect 11931 12804 13360 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14200 12804 14933 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1946 12764 1952 12776
rect 1443 12736 1952 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 4985 12767 5043 12773
rect 4985 12764 4997 12767
rect 4764 12736 4997 12764
rect 4764 12724 4770 12736
rect 4985 12733 4997 12736
rect 5031 12764 5043 12767
rect 5534 12764 5540 12776
rect 5031 12736 5540 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 8478 12764 8484 12776
rect 8435 12736 8484 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12124 12736 12265 12764
rect 12124 12724 12130 12736
rect 12253 12733 12265 12736
rect 12299 12764 12311 12767
rect 12894 12764 12900 12776
rect 12299 12736 12900 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13078 12764 13084 12776
rect 13039 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13446 12764 13452 12776
rect 13219 12736 13452 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 5077 12699 5135 12705
rect 5077 12696 5089 12699
rect 4571 12668 5089 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 5077 12665 5089 12668
rect 5123 12696 5135 12699
rect 5350 12696 5356 12708
rect 5123 12668 5356 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 10134 12696 10140 12708
rect 10095 12668 10140 12696
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 1762 12628 1768 12640
rect 1627 12600 1768 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 4890 12628 4896 12640
rect 4663 12600 4896 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 12710 12628 12716 12640
rect 12671 12600 12716 12628
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 13188 12628 13216 12727
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 12952 12600 13216 12628
rect 12952 12588 12958 12600
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14200 12637 14228 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 16390 12832 16396 12844
rect 15519 12804 16396 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 16540 12804 16633 12832
rect 16540 12792 16546 12804
rect 23842 12792 23848 12844
rect 23900 12832 23906 12844
rect 24228 12841 24256 12872
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 25225 12903 25283 12909
rect 25225 12869 25237 12903
rect 25271 12900 25283 12903
rect 25271 12872 26372 12900
rect 25271 12869 25283 12872
rect 25225 12863 25283 12869
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23900 12804 24225 12832
rect 23900 12792 23906 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 25498 12832 25504 12844
rect 24360 12804 24405 12832
rect 25459 12804 25504 12832
rect 24360 12792 24366 12804
rect 25498 12792 25504 12804
rect 25556 12832 25562 12844
rect 26344 12841 26372 12872
rect 27264 12841 27292 12940
rect 26329 12835 26387 12841
rect 25556 12804 26096 12832
rect 25556 12792 25562 12804
rect 14734 12764 14740 12776
rect 14695 12736 14740 12764
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15102 12764 15108 12776
rect 14875 12736 15108 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 16264 12736 16313 12764
rect 16264 12724 16270 12736
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 16942 12724 16948 12776
rect 17000 12764 17006 12776
rect 18690 12764 18696 12776
rect 17000 12736 18696 12764
rect 17000 12724 17006 12736
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 23109 12767 23167 12773
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 24121 12767 24179 12773
rect 24121 12764 24133 12767
rect 23155 12736 24133 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 24121 12733 24133 12736
rect 24167 12764 24179 12767
rect 24854 12764 24860 12776
rect 24167 12736 24860 12764
rect 24167 12733 24179 12736
rect 24121 12727 24179 12733
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 25682 12724 25688 12776
rect 25740 12724 25746 12776
rect 26068 12773 26096 12804
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 27249 12835 27307 12841
rect 26375 12804 26832 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26053 12767 26111 12773
rect 26053 12733 26065 12767
rect 26099 12764 26111 12767
rect 26418 12764 26424 12776
rect 26099 12736 26424 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 26694 12764 26700 12776
rect 26655 12736 26700 12764
rect 26694 12724 26700 12736
rect 26752 12724 26758 12776
rect 26804 12764 26832 12804
rect 27249 12801 27261 12835
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27430 12764 27436 12776
rect 26804 12736 27436 12764
rect 27430 12724 27436 12736
rect 27488 12724 27494 12776
rect 23474 12696 23480 12708
rect 23435 12668 23480 12696
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 24302 12696 24308 12708
rect 23768 12668 24308 12696
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 13964 12600 14197 12628
rect 13964 12588 13970 12600
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14366 12628 14372 12640
rect 14327 12600 14372 12628
rect 14185 12591 14243 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 18322 12628 18328 12640
rect 18283 12600 18328 12628
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 23768 12637 23796 12668
rect 24302 12656 24308 12668
rect 24360 12656 24366 12708
rect 25700 12696 25728 12724
rect 25700 12668 25820 12696
rect 23753 12631 23811 12637
rect 23753 12597 23765 12631
rect 23799 12597 23811 12631
rect 25682 12628 25688 12640
rect 25643 12600 25688 12628
rect 23753 12591 23811 12597
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 25792 12628 25820 12668
rect 25866 12656 25872 12708
rect 25924 12696 25930 12708
rect 27522 12696 27528 12708
rect 25924 12668 27528 12696
rect 25924 12656 25930 12668
rect 27522 12656 27528 12668
rect 27580 12656 27586 12708
rect 26145 12631 26203 12637
rect 26145 12628 26157 12631
rect 25792 12600 26157 12628
rect 26145 12597 26157 12600
rect 26191 12597 26203 12631
rect 26145 12591 26203 12597
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 5592 12396 6193 12424
rect 5592 12384 5598 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 6181 12387 6239 12393
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 8113 12427 8171 12433
rect 8113 12393 8125 12427
rect 8159 12424 8171 12427
rect 8202 12424 8208 12436
rect 8159 12396 8208 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 13078 12424 13084 12436
rect 12851 12396 13084 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13173 12427 13231 12433
rect 13173 12393 13185 12427
rect 13219 12424 13231 12427
rect 13354 12424 13360 12436
rect 13219 12396 13360 12424
rect 13219 12393 13231 12396
rect 13173 12387 13231 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 16853 12427 16911 12433
rect 16853 12393 16865 12427
rect 16899 12424 16911 12427
rect 17310 12424 17316 12436
rect 16899 12396 17316 12424
rect 16899 12393 16911 12396
rect 16853 12387 16911 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 23842 12424 23848 12436
rect 23803 12396 23848 12424
rect 23842 12384 23848 12396
rect 23900 12384 23906 12436
rect 24854 12424 24860 12436
rect 24815 12396 24860 12424
rect 24854 12384 24860 12396
rect 24912 12384 24918 12436
rect 25314 12424 25320 12436
rect 25227 12396 25320 12424
rect 25314 12384 25320 12396
rect 25372 12424 25378 12436
rect 25682 12424 25688 12436
rect 25372 12396 25688 12424
rect 25372 12384 25378 12396
rect 25682 12384 25688 12396
rect 25740 12384 25746 12436
rect 27157 12427 27215 12433
rect 27157 12393 27169 12427
rect 27203 12424 27215 12427
rect 27430 12424 27436 12436
rect 27203 12396 27436 12424
rect 27203 12393 27215 12396
rect 27157 12387 27215 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16482 12356 16488 12368
rect 16071 12328 16488 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 21168 12359 21226 12365
rect 21168 12325 21180 12359
rect 21214 12356 21226 12359
rect 21266 12356 21272 12368
rect 21214 12328 21272 12356
rect 21214 12325 21226 12328
rect 21168 12319 21226 12325
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 25225 12359 25283 12365
rect 25225 12325 25237 12359
rect 25271 12356 25283 12359
rect 25590 12356 25596 12368
rect 25271 12328 25596 12356
rect 25271 12325 25283 12328
rect 25225 12319 25283 12325
rect 25590 12316 25596 12328
rect 25648 12356 25654 12368
rect 26142 12356 26148 12368
rect 25648 12328 26148 12356
rect 25648 12316 25654 12328
rect 26142 12316 26148 12328
rect 26200 12316 26206 12368
rect 4982 12288 4988 12300
rect 4895 12260 4988 12288
rect 4982 12248 4988 12260
rect 5040 12288 5046 12300
rect 5442 12288 5448 12300
rect 5040 12260 5448 12288
rect 5040 12248 5046 12260
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 13446 12288 13452 12300
rect 13403 12260 13452 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 17494 12288 17500 12300
rect 17455 12260 17500 12288
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 21910 12288 21916 12300
rect 20947 12260 21916 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 22738 12248 22744 12300
rect 22796 12288 22802 12300
rect 23842 12288 23848 12300
rect 22796 12260 23848 12288
rect 22796 12248 22802 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 26510 12288 26516 12300
rect 26471 12260 26516 12288
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 5074 12220 5080 12232
rect 5035 12192 5080 12220
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5258 12220 5264 12232
rect 5219 12192 5264 12220
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17586 12220 17592 12232
rect 17184 12192 17592 12220
rect 17184 12180 17190 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 24946 12180 24952 12232
rect 25004 12220 25010 12232
rect 25130 12220 25136 12232
rect 25004 12192 25136 12220
rect 25004 12180 25010 12192
rect 25130 12180 25136 12192
rect 25188 12220 25194 12232
rect 25409 12223 25467 12229
rect 25409 12220 25421 12223
rect 25188 12192 25421 12220
rect 25188 12180 25194 12192
rect 25409 12189 25421 12192
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 4614 12084 4620 12096
rect 4575 12056 4620 12084
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 8478 12084 8484 12096
rect 8439 12056 8484 12084
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 9732 12056 9873 12084
rect 9732 12044 9738 12056
rect 9861 12053 9873 12056
rect 9907 12084 9919 12087
rect 10134 12084 10140 12096
rect 9907 12056 10140 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 10321 12087 10379 12093
rect 10321 12053 10333 12087
rect 10367 12084 10379 12087
rect 10870 12084 10876 12096
rect 10367 12056 10876 12084
rect 10367 12053 10379 12056
rect 10321 12047 10379 12053
rect 10870 12044 10876 12056
rect 10928 12084 10934 12096
rect 11146 12084 11152 12096
rect 10928 12056 11152 12084
rect 10928 12044 10934 12056
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 14642 12084 14648 12096
rect 14603 12056 14648 12084
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 17129 12087 17187 12093
rect 17129 12053 17141 12087
rect 17175 12084 17187 12087
rect 17218 12084 17224 12096
rect 17175 12056 17224 12084
rect 17175 12053 17187 12056
rect 17129 12047 17187 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 21818 12044 21824 12096
rect 21876 12084 21882 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 21876 12056 22293 12084
rect 21876 12044 21882 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 26326 12044 26332 12096
rect 26384 12084 26390 12096
rect 26697 12087 26755 12093
rect 26697 12084 26709 12087
rect 26384 12056 26709 12084
rect 26384 12044 26390 12056
rect 26697 12053 26709 12056
rect 26743 12053 26755 12087
rect 26697 12047 26755 12053
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 5074 11880 5080 11892
rect 4755 11852 5080 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 5074 11840 5080 11852
rect 5132 11880 5138 11892
rect 5721 11883 5779 11889
rect 5721 11880 5733 11883
rect 5132 11852 5733 11880
rect 5132 11840 5138 11852
rect 5721 11849 5733 11852
rect 5767 11849 5779 11883
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 5721 11843 5779 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 17494 11880 17500 11892
rect 12768 11852 13860 11880
rect 17455 11852 17500 11880
rect 12768 11840 12774 11852
rect 12529 11815 12587 11821
rect 12529 11781 12541 11815
rect 12575 11812 12587 11815
rect 13832 11812 13860 11852
rect 17494 11840 17500 11852
rect 17552 11880 17558 11892
rect 21266 11880 21272 11892
rect 17552 11852 18092 11880
rect 21227 11852 21272 11880
rect 17552 11840 17558 11852
rect 14737 11815 14795 11821
rect 14737 11812 14749 11815
rect 12575 11784 13768 11812
rect 12575 11781 12587 11784
rect 12529 11775 12587 11781
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 5224 11716 5273 11744
rect 5224 11704 5230 11716
rect 5261 11713 5273 11716
rect 5307 11713 5319 11747
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 5261 11707 5319 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13354 11744 13360 11756
rect 13219 11716 13360 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4522 11676 4528 11688
rect 4304 11648 4528 11676
rect 4304 11636 4310 11648
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 5074 11676 5080 11688
rect 4663 11648 5080 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7374 11676 7380 11688
rect 7331 11648 7380 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9355 11648 9781 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9769 11645 9781 11648
rect 9815 11676 9827 11679
rect 10502 11676 10508 11688
rect 9815 11648 10508 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 2124 11611 2182 11617
rect 2124 11608 2136 11611
rect 1811 11580 2136 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 2124 11577 2136 11580
rect 2170 11608 2182 11611
rect 2682 11608 2688 11620
rect 2170 11580 2688 11608
rect 2170 11577 2182 11580
rect 2124 11571 2182 11577
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 3881 11611 3939 11617
rect 3881 11608 3893 11611
rect 3252 11580 3893 11608
rect 3252 11549 3280 11580
rect 3881 11577 3893 11580
rect 3927 11608 3939 11611
rect 3970 11608 3976 11620
rect 3927 11580 3976 11608
rect 3927 11577 3939 11580
rect 3881 11571 3939 11577
rect 3970 11568 3976 11580
rect 4028 11608 4034 11620
rect 5258 11608 5264 11620
rect 4028 11580 5264 11608
rect 4028 11568 4034 11580
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 7190 11608 7196 11620
rect 7103 11580 7196 11608
rect 7190 11568 7196 11580
rect 7248 11608 7254 11620
rect 7530 11611 7588 11617
rect 7530 11608 7542 11611
rect 7248 11580 7542 11608
rect 7248 11568 7254 11580
rect 7530 11577 7542 11580
rect 7576 11577 7588 11611
rect 10014 11611 10072 11617
rect 10014 11608 10026 11611
rect 7530 11571 7588 11577
rect 9600 11580 10026 11608
rect 3237 11543 3295 11549
rect 3237 11509 3249 11543
rect 3283 11509 3295 11543
rect 4246 11540 4252 11552
rect 4159 11512 4252 11540
rect 3237 11503 3295 11509
rect 4246 11500 4252 11512
rect 4304 11540 4310 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 4304 11512 5181 11540
rect 4304 11500 4310 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 9600 11549 9628 11580
rect 10014 11577 10026 11580
rect 10060 11577 10072 11611
rect 10014 11571 10072 11577
rect 11885 11611 11943 11617
rect 11885 11577 11897 11611
rect 11931 11608 11943 11611
rect 12342 11608 12348 11620
rect 11931 11580 12348 11608
rect 11931 11577 11943 11580
rect 11885 11571 11943 11577
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 13740 11617 13768 11784
rect 13832 11784 14749 11812
rect 13832 11753 13860 11784
rect 14737 11781 14749 11784
rect 14783 11781 14795 11815
rect 14737 11775 14795 11781
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 18064 11753 18092 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 24946 11880 24952 11892
rect 24907 11852 24952 11880
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25314 11880 25320 11892
rect 25275 11852 25320 11880
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 25590 11880 25596 11892
rect 25551 11852 25596 11880
rect 25590 11840 25596 11852
rect 25648 11840 25654 11892
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 26568 11852 27353 11880
rect 26568 11840 26574 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 14369 11747 14427 11753
rect 14369 11744 14381 11747
rect 13964 11716 14381 11744
rect 13964 11704 13970 11716
rect 14369 11713 14381 11716
rect 14415 11713 14427 11747
rect 14369 11707 14427 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 18049 11707 18107 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 19260 11676 19288 11704
rect 26418 11676 26424 11688
rect 18012 11648 19288 11676
rect 26379 11648 26424 11676
rect 18012 11636 18018 11648
rect 26418 11636 26424 11648
rect 26476 11676 26482 11688
rect 26973 11679 27031 11685
rect 26973 11676 26985 11679
rect 26476 11648 26985 11676
rect 26476 11636 26482 11648
rect 26973 11645 26985 11648
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12400 11580 12909 11608
rect 12400 11568 12406 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 13725 11611 13783 11617
rect 13725 11577 13737 11611
rect 13771 11608 13783 11611
rect 15197 11611 15255 11617
rect 15197 11608 15209 11611
rect 13771 11580 15209 11608
rect 13771 11577 13783 11580
rect 13725 11571 13783 11577
rect 15197 11577 15209 11580
rect 15243 11577 15255 11611
rect 15197 11571 15255 11577
rect 16853 11611 16911 11617
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 17770 11608 17776 11620
rect 16899 11580 17776 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 19150 11608 19156 11620
rect 19111 11580 19156 11608
rect 19150 11568 19156 11580
rect 19208 11608 19214 11620
rect 19490 11611 19548 11617
rect 19490 11608 19502 11611
rect 19208 11580 19502 11608
rect 19208 11568 19214 11580
rect 19490 11577 19502 11580
rect 19536 11577 19548 11611
rect 19490 11571 19548 11577
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 7892 11512 8677 11540
rect 7892 11500 7898 11512
rect 8665 11509 8677 11512
rect 8711 11540 8723 11543
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 8711 11512 9597 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 9585 11503 9643 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11388 11512 12173 11540
rect 11388 11500 11394 11512
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12986 11540 12992 11552
rect 12207 11512 12992 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13357 11543 13415 11549
rect 13357 11509 13369 11543
rect 13403 11540 13415 11543
rect 13630 11540 13636 11552
rect 13403 11512 13636 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 17126 11540 17132 11552
rect 17087 11512 17132 11540
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 19116 11512 20637 11540
rect 19116 11500 19122 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 21637 11543 21695 11549
rect 21637 11509 21649 11543
rect 21683 11540 21695 11543
rect 21910 11540 21916 11552
rect 21683 11512 21916 11540
rect 21683 11509 21695 11512
rect 21637 11503 21695 11509
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 26602 11540 26608 11552
rect 26563 11512 26608 11540
rect 26602 11500 26608 11512
rect 26660 11500 26666 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 5166 11336 5172 11348
rect 5127 11308 5172 11336
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 7650 11336 7656 11348
rect 7611 11308 7656 11336
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 12400 11308 12541 11336
rect 12400 11296 12406 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11336 13139 11339
rect 13354 11336 13360 11348
rect 13127 11308 13360 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 13998 11336 14004 11348
rect 13688 11308 14004 11336
rect 13688 11296 13694 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11336 14151 11339
rect 14366 11336 14372 11348
rect 14139 11308 14372 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 17310 11336 17316 11348
rect 17223 11308 17316 11336
rect 17310 11296 17316 11308
rect 17368 11336 17374 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 17368 11308 18429 11336
rect 17368 11296 17374 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18417 11299 18475 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 17218 11268 17224 11280
rect 17179 11240 17224 11268
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2038 11200 2044 11212
rect 1443 11172 2044 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 22005 11203 22063 11209
rect 22005 11200 22017 11203
rect 21968 11172 22017 11200
rect 21968 11160 21974 11172
rect 22005 11169 22017 11172
rect 22051 11169 22063 11203
rect 22005 11163 22063 11169
rect 22272 11203 22330 11209
rect 22272 11169 22284 11203
rect 22318 11200 22330 11203
rect 22830 11200 22836 11212
rect 22318 11172 22836 11200
rect 22318 11169 22330 11172
rect 22272 11163 22330 11169
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4212 11104 4537 11132
rect 4212 11092 4218 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5258 11132 5264 11144
rect 4755 11104 5264 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 7742 11132 7748 11144
rect 7703 11104 7748 11132
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 14274 11132 14280 11144
rect 7892 11104 7937 11132
rect 14235 11104 14280 11132
rect 7892 11092 7898 11104
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 16942 11092 16948 11144
rect 17000 11132 17006 11144
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17000 11104 17417 11132
rect 17000 11092 17006 11104
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18564 11104 18889 11132
rect 18564 11092 18570 11104
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 19058 11132 19064 11144
rect 19019 11104 19064 11132
rect 18877 11095 18935 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 4062 11064 4068 11076
rect 4023 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 7558 11064 7564 11076
rect 7331 11036 7564 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 13354 11064 13360 11076
rect 13315 11036 13360 11064
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13722 11064 13728 11076
rect 13679 11036 13728 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 16850 11064 16856 11076
rect 16811 11036 16856 11064
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 17770 11024 17776 11076
rect 17828 11064 17834 11076
rect 19076 11064 19104 11092
rect 17828 11036 19104 11064
rect 21913 11067 21971 11073
rect 17828 11024 17834 11036
rect 21913 11033 21925 11067
rect 21959 11064 21971 11067
rect 21959 11036 22048 11064
rect 21959 11033 21971 11036
rect 21913 11027 21971 11033
rect 22020 10996 22048 11036
rect 22186 10996 22192 11008
rect 22020 10968 22192 10996
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 23382 10996 23388 11008
rect 23343 10968 23388 10996
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1544 10764 1593 10792
rect 1544 10752 1550 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 2038 10792 2044 10804
rect 1999 10764 2044 10792
rect 1581 10755 1639 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3476 10764 3617 10792
rect 3476 10752 3482 10764
rect 3605 10761 3617 10764
rect 3651 10792 3663 10795
rect 4062 10792 4068 10804
rect 3651 10764 4068 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7834 10792 7840 10804
rect 7423 10764 7840 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 14332 10764 14381 10792
rect 14332 10752 14338 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 17310 10792 17316 10804
rect 17271 10764 17316 10792
rect 14369 10755 14427 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17770 10792 17776 10804
rect 17731 10764 17776 10792
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18782 10792 18788 10804
rect 18555 10764 18788 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21637 10795 21695 10801
rect 21637 10792 21649 10795
rect 20772 10764 21649 10792
rect 20772 10752 20778 10764
rect 21637 10761 21649 10764
rect 21683 10761 21695 10795
rect 22830 10792 22836 10804
rect 22791 10764 22836 10792
rect 21637 10755 21695 10761
rect 3237 10727 3295 10733
rect 3237 10693 3249 10727
rect 3283 10724 3295 10727
rect 4430 10724 4436 10736
rect 3283 10696 4436 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 7742 10724 7748 10736
rect 7703 10696 7748 10724
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 16577 10727 16635 10733
rect 16577 10693 16589 10727
rect 16623 10724 16635 10727
rect 17218 10724 17224 10736
rect 16623 10696 17224 10724
rect 16623 10693 16635 10696
rect 16577 10687 16635 10693
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 18877 10727 18935 10733
rect 18877 10724 18889 10727
rect 17920 10696 18889 10724
rect 17920 10684 17926 10696
rect 18877 10693 18889 10696
rect 18923 10724 18935 10727
rect 20622 10724 20628 10736
rect 18923 10696 20628 10724
rect 18923 10693 18935 10696
rect 18877 10687 18935 10693
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 3970 10656 3976 10668
rect 3931 10628 3976 10656
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5166 10656 5172 10668
rect 5123 10628 5172 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5166 10616 5172 10628
rect 5224 10616 5230 10668
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7708 10628 8033 10656
rect 7708 10616 7714 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 21652 10656 21680 10755
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 26510 10792 26516 10804
rect 26471 10764 26516 10792
rect 26510 10752 26516 10764
rect 26568 10752 26574 10804
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 12943 10628 13124 10656
rect 21652 10628 22477 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2406 10588 2412 10600
rect 1443 10560 2412 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 12986 10588 12992 10600
rect 12947 10560 12992 10588
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13096 10588 13124 10628
rect 22465 10625 22477 10628
rect 22511 10656 22523 10659
rect 23382 10656 23388 10668
rect 22511 10628 23388 10656
rect 22511 10625 22523 10628
rect 22465 10619 22523 10625
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 13256 10591 13314 10597
rect 13256 10588 13268 10591
rect 13096 10560 13268 10588
rect 13256 10557 13268 10560
rect 13302 10588 13314 10591
rect 13630 10588 13636 10600
rect 13302 10560 13636 10588
rect 13302 10557 13314 10560
rect 13256 10551 13314 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 18932 10560 19073 10588
rect 18932 10548 18938 10560
rect 19061 10557 19073 10560
rect 19107 10588 19119 10591
rect 19337 10591 19395 10597
rect 19337 10588 19349 10591
rect 19107 10560 19349 10588
rect 19107 10557 19119 10560
rect 19061 10551 19119 10557
rect 19337 10557 19349 10560
rect 19383 10557 19395 10591
rect 24210 10588 24216 10600
rect 24171 10560 24216 10588
rect 19337 10551 19395 10557
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 24458 10523 24516 10529
rect 24458 10520 24470 10523
rect 24044 10492 24470 10520
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4798 10452 4804 10464
rect 4387 10424 4804 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 16942 10452 16948 10464
rect 4948 10424 4993 10452
rect 16903 10424 16948 10452
rect 4948 10412 4954 10424
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 20772 10424 21833 10452
rect 20772 10412 20778 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 22186 10452 22192 10464
rect 22147 10424 22192 10452
rect 21821 10415 21879 10421
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22336 10424 22381 10452
rect 22336 10412 22342 10424
rect 23566 10412 23572 10464
rect 23624 10452 23630 10464
rect 24044 10461 24072 10492
rect 24458 10489 24470 10492
rect 24504 10489 24516 10523
rect 24458 10483 24516 10489
rect 24029 10455 24087 10461
rect 24029 10452 24041 10455
rect 23624 10424 24041 10452
rect 23624 10412 23630 10424
rect 24029 10421 24041 10424
rect 24075 10421 24087 10455
rect 25590 10452 25596 10464
rect 25551 10424 25596 10452
rect 24029 10415 24087 10421
rect 25590 10412 25596 10424
rect 25648 10412 25654 10464
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 26697 10455 26755 10461
rect 26697 10452 26709 10455
rect 26660 10424 26709 10452
rect 26660 10412 26666 10424
rect 26697 10421 26709 10424
rect 26743 10421 26755 10455
rect 26697 10415 26755 10421
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2682 10208 2688 10260
rect 2740 10248 2746 10260
rect 2774 10248 2780 10260
rect 2740 10220 2780 10248
rect 2740 10208 2746 10220
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 4890 10208 4896 10220
rect 4948 10248 4954 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4948 10220 5089 10248
rect 4948 10208 4954 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5077 10211 5135 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 14366 10248 14372 10260
rect 14139 10220 14372 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 18966 10208 18972 10260
rect 19024 10248 19030 10260
rect 19245 10251 19303 10257
rect 19245 10248 19257 10251
rect 19024 10220 19257 10248
rect 19024 10208 19030 10220
rect 19245 10217 19257 10220
rect 19291 10217 19303 10251
rect 19245 10211 19303 10217
rect 21545 10251 21603 10257
rect 21545 10217 21557 10251
rect 21591 10248 21603 10251
rect 21818 10248 21824 10260
rect 21591 10220 21824 10248
rect 21591 10217 21603 10220
rect 21545 10211 21603 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 21913 10251 21971 10257
rect 21913 10217 21925 10251
rect 21959 10248 21971 10251
rect 22278 10248 22284 10260
rect 21959 10220 22284 10248
rect 21959 10217 21971 10220
rect 21913 10211 21971 10217
rect 22278 10208 22284 10220
rect 22336 10248 22342 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22336 10220 22385 10248
rect 22336 10208 22342 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 24210 10248 24216 10260
rect 24171 10220 24216 10248
rect 22373 10211 22431 10217
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 24854 10248 24860 10260
rect 24815 10220 24860 10248
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 25314 10248 25320 10260
rect 25227 10220 25320 10248
rect 25314 10208 25320 10220
rect 25372 10248 25378 10260
rect 26513 10251 26571 10257
rect 26513 10248 26525 10251
rect 25372 10220 26525 10248
rect 25372 10208 25378 10220
rect 26513 10217 26525 10220
rect 26559 10217 26571 10251
rect 26970 10248 26976 10260
rect 26931 10220 26976 10248
rect 26513 10211 26571 10217
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 5537 10183 5595 10189
rect 5537 10180 5549 10183
rect 5040 10152 5549 10180
rect 5040 10140 5046 10152
rect 5537 10149 5549 10152
rect 5583 10149 5595 10183
rect 12986 10180 12992 10192
rect 5537 10143 5595 10149
rect 10244 10152 12992 10180
rect 10244 10124 10272 10152
rect 12986 10140 12992 10152
rect 13044 10180 13050 10192
rect 13725 10183 13783 10189
rect 13044 10152 13124 10180
rect 13044 10140 13050 10152
rect 1664 10115 1722 10121
rect 1664 10081 1676 10115
rect 1710 10112 1722 10115
rect 2222 10112 2228 10124
rect 1710 10084 2228 10112
rect 1710 10081 1722 10084
rect 1664 10075 1722 10081
rect 2222 10072 2228 10084
rect 2280 10072 2286 10124
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4120 10084 4537 10112
rect 4120 10072 4126 10084
rect 4525 10081 4537 10084
rect 4571 10112 4583 10115
rect 5166 10112 5172 10124
rect 4571 10084 5172 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 10226 10112 10232 10124
rect 10139 10084 10232 10112
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10496 10115 10554 10121
rect 10496 10081 10508 10115
rect 10542 10112 10554 10115
rect 10870 10112 10876 10124
rect 10542 10084 10876 10112
rect 10542 10081 10554 10084
rect 10496 10075 10554 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1412 9908 1440 10007
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5500 10016 5641 10044
rect 5500 10004 5506 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 2332 9948 5212 9976
rect 2130 9908 2136 9920
rect 1412 9880 2136 9908
rect 2130 9868 2136 9880
rect 2188 9908 2194 9920
rect 2332 9908 2360 9948
rect 2188 9880 2360 9908
rect 2188 9868 2194 9880
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 3510 9908 3516 9920
rect 2832 9880 2877 9908
rect 3471 9880 3516 9908
rect 2832 9868 2838 9880
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 5184 9908 5212 9948
rect 6914 9908 6920 9920
rect 5184 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9908 6978 9920
rect 7834 9908 7840 9920
rect 6972 9880 7840 9908
rect 6972 9868 6978 9880
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 11606 9908 11612 9920
rect 11567 9880 11612 9908
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13096 9917 13124 10152
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 13906 10180 13912 10192
rect 13771 10152 13912 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 13906 10140 13912 10152
rect 13964 10180 13970 10192
rect 14274 10180 14280 10192
rect 13964 10152 14280 10180
rect 13964 10140 13970 10152
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 18782 10180 18788 10192
rect 18472 10152 18788 10180
rect 18472 10140 18478 10152
rect 18782 10140 18788 10152
rect 18840 10180 18846 10192
rect 19153 10183 19211 10189
rect 19153 10180 19165 10183
rect 18840 10152 19165 10180
rect 18840 10140 18846 10152
rect 19153 10149 19165 10152
rect 19199 10149 19211 10183
rect 19153 10143 19211 10149
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 15838 10121 15844 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 14056 10084 14381 10112
rect 14056 10072 14062 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 15832 10112 15844 10121
rect 15799 10084 15844 10112
rect 14369 10075 14427 10081
rect 15832 10075 15844 10084
rect 15838 10072 15844 10075
rect 15896 10072 15902 10124
rect 20622 10112 20628 10124
rect 20583 10084 20628 10112
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 22738 10112 22744 10124
rect 22699 10084 22744 10112
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 25225 10115 25283 10121
rect 25225 10081 25237 10115
rect 25271 10112 25283 10115
rect 25682 10112 25688 10124
rect 25271 10084 25688 10112
rect 25271 10081 25283 10084
rect 25225 10075 25283 10081
rect 25682 10072 25688 10084
rect 25740 10072 25746 10124
rect 26878 10112 26884 10124
rect 26839 10084 26884 10112
rect 26878 10072 26884 10084
rect 26936 10072 26942 10124
rect 15562 10044 15568 10056
rect 15523 10016 15568 10044
rect 15562 10004 15568 10016
rect 15620 10004 15626 10056
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 19208 10016 19349 10044
rect 19208 10004 19214 10016
rect 19337 10013 19349 10016
rect 19383 10013 19395 10047
rect 22830 10044 22836 10056
rect 22791 10016 22836 10044
rect 19337 10007 19395 10013
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 22922 10004 22928 10056
rect 22980 10044 22986 10056
rect 22980 10016 23025 10044
rect 22980 10004 22986 10016
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25409 10047 25467 10053
rect 25409 10044 25421 10047
rect 24912 10016 25421 10044
rect 24912 10004 24918 10016
rect 25409 10013 25421 10016
rect 25455 10044 25467 10047
rect 25590 10044 25596 10056
rect 25455 10016 25596 10044
rect 25455 10013 25467 10016
rect 25409 10007 25467 10013
rect 25590 10004 25596 10016
rect 25648 10004 25654 10056
rect 27065 10047 27123 10053
rect 27065 10013 27077 10047
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 18138 9976 18144 9988
rect 18099 9948 18144 9976
rect 18138 9936 18144 9948
rect 18196 9936 18202 9988
rect 22281 9979 22339 9985
rect 22281 9945 22293 9979
rect 22327 9976 22339 9979
rect 24210 9976 24216 9988
rect 22327 9948 24216 9976
rect 22327 9945 22339 9948
rect 22281 9939 22339 9945
rect 13081 9911 13139 9917
rect 12492 9880 12537 9908
rect 12492 9868 12498 9880
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13630 9908 13636 9920
rect 13127 9880 13636 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 16942 9908 16948 9920
rect 16855 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9908 17006 9920
rect 17402 9908 17408 9920
rect 17000 9880 17408 9908
rect 17000 9868 17006 9880
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 17773 9911 17831 9917
rect 17773 9877 17785 9911
rect 17819 9908 17831 9911
rect 17862 9908 17868 9920
rect 17819 9880 17868 9908
rect 17819 9877 17831 9880
rect 17773 9871 17831 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18564 9880 18797 9908
rect 18564 9868 18570 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18785 9871 18843 9877
rect 19794 9868 19800 9920
rect 19852 9908 19858 9920
rect 19889 9911 19947 9917
rect 19889 9908 19901 9911
rect 19852 9880 19901 9908
rect 19852 9868 19858 9880
rect 19889 9877 19901 9880
rect 19935 9908 19947 9911
rect 20162 9908 20168 9920
rect 19935 9880 20168 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 20438 9908 20444 9920
rect 20399 9880 20444 9908
rect 20438 9868 20444 9880
rect 20496 9908 20502 9920
rect 21910 9908 21916 9920
rect 20496 9880 21916 9908
rect 20496 9868 20502 9880
rect 21910 9868 21916 9880
rect 21968 9908 21974 9920
rect 22296 9908 22324 9939
rect 24210 9936 24216 9948
rect 24268 9936 24274 9988
rect 27080 9976 27108 10007
rect 26436 9948 27108 9976
rect 26436 9920 26464 9948
rect 21968 9880 22324 9908
rect 21968 9868 21974 9880
rect 23566 9868 23572 9920
rect 23624 9908 23630 9920
rect 23661 9911 23719 9917
rect 23661 9908 23673 9911
rect 23624 9880 23673 9908
rect 23624 9868 23630 9880
rect 23661 9877 23673 9880
rect 23707 9908 23719 9911
rect 25869 9911 25927 9917
rect 25869 9908 25881 9911
rect 23707 9880 25881 9908
rect 23707 9877 23719 9880
rect 23661 9871 23719 9877
rect 25869 9877 25881 9880
rect 25915 9908 25927 9911
rect 26418 9908 26424 9920
rect 25915 9880 26424 9908
rect 25915 9877 25927 9880
rect 25869 9871 25927 9877
rect 26418 9868 26424 9880
rect 26476 9868 26482 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 2317 9707 2375 9713
rect 2317 9704 2329 9707
rect 2280 9676 2329 9704
rect 2280 9664 2286 9676
rect 2317 9673 2329 9676
rect 2363 9673 2375 9707
rect 3418 9704 3424 9716
rect 3379 9676 3424 9704
rect 2317 9667 2375 9673
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 4706 9664 4712 9716
rect 4764 9664 4770 9716
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 10226 9664 10232 9676
rect 10284 9704 10290 9716
rect 10321 9707 10379 9713
rect 10321 9704 10333 9707
rect 10284 9676 10333 9704
rect 10284 9664 10290 9676
rect 10321 9673 10333 9676
rect 10367 9673 10379 9707
rect 13906 9704 13912 9716
rect 13867 9676 13912 9704
rect 10321 9667 10379 9673
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 16025 9707 16083 9713
rect 16025 9704 16037 9707
rect 15896 9676 16037 9704
rect 15896 9664 15902 9676
rect 16025 9673 16037 9676
rect 16071 9704 16083 9707
rect 17589 9707 17647 9713
rect 17589 9704 17601 9707
rect 16071 9676 17601 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 17589 9673 17601 9676
rect 17635 9704 17647 9707
rect 17770 9704 17776 9716
rect 17635 9676 17776 9704
rect 17635 9673 17647 9676
rect 17589 9667 17647 9673
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 19024 9676 19073 9704
rect 19024 9664 19030 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19061 9667 19119 9673
rect 20622 9664 20628 9716
rect 20680 9664 20686 9716
rect 22557 9707 22615 9713
rect 22557 9673 22569 9707
rect 22603 9704 22615 9707
rect 22922 9704 22928 9716
rect 22603 9676 22928 9704
rect 22603 9673 22615 9676
rect 22557 9667 22615 9673
rect 22922 9664 22928 9676
rect 22980 9704 22986 9716
rect 24854 9704 24860 9716
rect 22980 9676 24860 9704
rect 22980 9664 22986 9676
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 25314 9704 25320 9716
rect 25275 9676 25320 9704
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 26878 9704 26884 9716
rect 26839 9676 26884 9704
rect 26878 9664 26884 9676
rect 26936 9664 26942 9716
rect 26970 9664 26976 9716
rect 27028 9704 27034 9716
rect 27249 9707 27307 9713
rect 27249 9704 27261 9707
rect 27028 9676 27261 9704
rect 27028 9664 27034 9676
rect 27249 9673 27261 9676
rect 27295 9673 27307 9707
rect 27249 9667 27307 9673
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 2832 9540 3341 9568
rect 2832 9528 2838 9540
rect 3329 9537 3341 9540
rect 3375 9568 3387 9571
rect 4062 9568 4068 9580
rect 3375 9540 4068 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 1412 9432 1440 9463
rect 3510 9460 3516 9512
rect 3568 9500 3574 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 3568 9472 3801 9500
rect 3568 9460 3574 9472
rect 3789 9469 3801 9472
rect 3835 9500 3847 9503
rect 4614 9500 4620 9512
rect 3835 9472 4620 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 2038 9432 2044 9444
rect 1412 9404 2044 9432
rect 2038 9392 2044 9404
rect 2096 9392 2102 9444
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 4525 9435 4583 9441
rect 3660 9404 4200 9432
rect 3660 9392 3666 9404
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3881 9367 3939 9373
rect 3881 9333 3893 9367
rect 3927 9364 3939 9367
rect 4062 9364 4068 9376
rect 3927 9336 4068 9364
rect 3927 9333 3939 9336
rect 3881 9327 3939 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4172 9364 4200 9404
rect 4525 9401 4537 9435
rect 4571 9432 4583 9435
rect 4724 9432 4752 9664
rect 4798 9596 4804 9648
rect 4856 9636 4862 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4856 9608 4997 9636
rect 4856 9596 4862 9608
rect 4985 9605 4997 9608
rect 5031 9605 5043 9639
rect 4985 9599 5043 9605
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9605 9275 9639
rect 12158 9636 12164 9648
rect 12119 9608 12164 9636
rect 9217 9599 9275 9605
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5500 9540 5641 9568
rect 5500 9528 5506 9540
rect 5629 9537 5641 9540
rect 5675 9568 5687 9571
rect 5902 9568 5908 9580
rect 5675 9540 5908 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5902 9528 5908 9540
rect 5960 9568 5966 9580
rect 7834 9568 7840 9580
rect 5960 9540 6132 9568
rect 7795 9540 7840 9568
rect 5960 9528 5966 9540
rect 6104 9509 6132 9540
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 9232 9500 9260 9599
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 10870 9568 10876 9580
rect 10783 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9568 10934 9580
rect 12434 9568 12440 9580
rect 10928 9540 12440 9568
rect 10928 9528 10934 9540
rect 12434 9528 12440 9540
rect 12492 9568 12498 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12492 9540 13001 9568
rect 12492 9528 12498 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 13924 9568 13952 9664
rect 17788 9636 17816 9664
rect 20640 9636 20668 9664
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 17788 9608 18644 9636
rect 20640 9608 20913 9636
rect 17221 9571 17279 9577
rect 13924 9540 14136 9568
rect 12989 9531 13047 9537
rect 6135 9472 9260 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10468 9472 10517 9500
rect 10468 9460 10474 9472
rect 10505 9469 10517 9472
rect 10551 9500 10563 9503
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10551 9472 11161 9500
rect 10551 9469 10563 9472
rect 10505 9463 10563 9469
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 11149 9463 11207 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14108 9500 14136 9540
rect 17221 9537 17233 9571
rect 17267 9568 17279 9571
rect 18506 9568 18512 9580
rect 17267 9540 18512 9568
rect 17267 9537 17279 9540
rect 17221 9531 17279 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18616 9577 18644 9608
rect 20901 9605 20913 9608
rect 20947 9605 20959 9639
rect 20901 9599 20959 9605
rect 22738 9596 22744 9648
rect 22796 9636 22802 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 22796 9608 23673 9636
rect 22796 9596 22802 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 25774 9636 25780 9648
rect 25735 9608 25780 9636
rect 23661 9599 23719 9605
rect 25774 9596 25780 9608
rect 25832 9596 25838 9648
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9568 18659 9571
rect 19058 9568 19064 9580
rect 18647 9540 19064 9568
rect 18647 9537 18659 9540
rect 18601 9531 18659 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 20346 9568 20352 9580
rect 19208 9540 20352 9568
rect 19208 9528 19214 9540
rect 20346 9528 20352 9540
rect 20404 9568 20410 9580
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 20404 9540 20545 9568
rect 20404 9528 20410 9540
rect 20533 9537 20545 9540
rect 20579 9568 20591 9571
rect 21818 9568 21824 9580
rect 20579 9540 21824 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 21818 9528 21824 9540
rect 21876 9568 21882 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21876 9540 22017 9568
rect 21876 9528 21882 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 24213 9571 24271 9577
rect 24213 9568 24225 9571
rect 23624 9540 24225 9568
rect 23624 9528 23630 9540
rect 24213 9537 24225 9540
rect 24259 9537 24271 9571
rect 26418 9568 26424 9580
rect 26379 9540 26424 9568
rect 24213 9531 24271 9537
rect 26418 9528 26424 9540
rect 26476 9528 26482 9580
rect 14257 9503 14315 9509
rect 14257 9500 14269 9503
rect 14108 9472 14269 9500
rect 14257 9469 14269 9472
rect 14303 9469 14315 9503
rect 17862 9500 17868 9512
rect 17823 9472 17868 9500
rect 14257 9463 14315 9469
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 18196 9472 18429 9500
rect 18196 9460 18202 9472
rect 18417 9469 18429 9472
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 19794 9460 19800 9512
rect 19852 9500 19858 9512
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19852 9472 20269 9500
rect 19852 9460 19858 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 21913 9503 21971 9509
rect 21913 9500 21925 9503
rect 20257 9463 20315 9469
rect 21284 9472 21925 9500
rect 5350 9432 5356 9444
rect 4571 9404 5356 9432
rect 4571 9401 4583 9404
rect 4525 9395 4583 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 8104 9435 8162 9441
rect 8104 9401 8116 9435
rect 8150 9401 8162 9435
rect 8104 9395 8162 9401
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4172 9336 4905 9364
rect 4893 9333 4905 9336
rect 4939 9364 4951 9367
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4939 9336 5457 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 5445 9333 5457 9336
rect 5491 9364 5503 9367
rect 5718 9364 5724 9376
rect 5491 9336 5724 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 8128 9364 8156 9395
rect 12158 9392 12164 9444
rect 12216 9432 12222 9444
rect 12894 9432 12900 9444
rect 12216 9404 12900 9432
rect 12216 9392 12222 9404
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 20349 9435 20407 9441
rect 20349 9432 20361 9435
rect 15068 9404 15608 9432
rect 15068 9392 15074 9404
rect 15580 9376 15608 9404
rect 19720 9404 20361 9432
rect 19720 9376 19748 9404
rect 20349 9401 20361 9404
rect 20395 9432 20407 9435
rect 20530 9432 20536 9444
rect 20395 9404 20536 9432
rect 20395 9401 20407 9404
rect 20349 9395 20407 9401
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 21284 9376 21312 9472
rect 21913 9469 21925 9472
rect 21959 9469 21971 9503
rect 23842 9500 23848 9512
rect 21913 9463 21971 9469
rect 23032 9472 23848 9500
rect 21542 9392 21548 9444
rect 21600 9432 21606 9444
rect 21821 9435 21879 9441
rect 21821 9432 21833 9435
rect 21600 9404 21833 9432
rect 21600 9392 21606 9404
rect 21821 9401 21833 9404
rect 21867 9432 21879 9435
rect 23032 9432 23060 9472
rect 23842 9460 23848 9472
rect 23900 9460 23906 9512
rect 25958 9460 25964 9512
rect 26016 9500 26022 9512
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 26016 9472 26249 9500
rect 26016 9460 26022 9472
rect 26237 9469 26249 9472
rect 26283 9500 26295 9503
rect 26602 9500 26608 9512
rect 26283 9472 26608 9500
rect 26283 9469 26295 9472
rect 26237 9463 26295 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 26878 9460 26884 9512
rect 26936 9500 26942 9512
rect 27433 9503 27491 9509
rect 27433 9500 27445 9503
rect 26936 9472 27445 9500
rect 26936 9460 26942 9472
rect 27433 9469 27445 9472
rect 27479 9500 27491 9503
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 27479 9472 27997 9500
rect 27479 9469 27491 9472
rect 27433 9463 27491 9469
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 21867 9404 23060 9432
rect 23109 9435 23167 9441
rect 21867 9401 21879 9404
rect 21821 9395 21879 9401
rect 23109 9401 23121 9435
rect 23155 9432 23167 9435
rect 23658 9432 23664 9444
rect 23155 9404 23664 9432
rect 23155 9401 23167 9404
rect 23109 9395 23167 9401
rect 23658 9392 23664 9404
rect 23716 9432 23722 9444
rect 24121 9435 24179 9441
rect 24121 9432 24133 9435
rect 23716 9404 24133 9432
rect 23716 9392 23722 9404
rect 24121 9401 24133 9404
rect 24167 9401 24179 9435
rect 24121 9395 24179 9401
rect 25774 9392 25780 9444
rect 25832 9432 25838 9444
rect 26329 9435 26387 9441
rect 26329 9432 26341 9435
rect 25832 9404 26341 9432
rect 25832 9392 25838 9404
rect 26329 9401 26341 9404
rect 26375 9401 26387 9435
rect 26329 9395 26387 9401
rect 8386 9364 8392 9376
rect 7791 9336 8392 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12308 9336 12449 9364
rect 12308 9324 12314 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 12584 9336 12817 9364
rect 12584 9324 12590 9336
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 12805 9327 12863 9333
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15381 9367 15439 9373
rect 15381 9364 15393 9367
rect 15160 9336 15393 9364
rect 15160 9324 15166 9336
rect 15381 9333 15393 9336
rect 15427 9333 15439 9367
rect 15381 9327 15439 9333
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 15620 9336 16405 9364
rect 15620 9324 15626 9336
rect 16393 9333 16405 9336
rect 16439 9364 16451 9367
rect 16666 9364 16672 9376
rect 16439 9336 16672 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16666 9324 16672 9336
rect 16724 9364 16730 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 16724 9336 17693 9364
rect 16724 9324 16730 9336
rect 17681 9333 17693 9336
rect 17727 9364 17739 9367
rect 17862 9364 17868 9376
rect 17727 9336 17868 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18230 9364 18236 9376
rect 18095 9336 18236 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 19702 9364 19708 9376
rect 19663 9336 19708 9364
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19886 9364 19892 9376
rect 19847 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21450 9364 21456 9376
rect 21411 9336 21456 9364
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9364 23814 9376
rect 24029 9367 24087 9373
rect 24029 9364 24041 9367
rect 23808 9336 24041 9364
rect 23808 9324 23814 9336
rect 24029 9333 24041 9336
rect 24075 9364 24087 9367
rect 24210 9364 24216 9376
rect 24075 9336 24216 9364
rect 24075 9333 24087 9336
rect 24029 9327 24087 9333
rect 24210 9324 24216 9336
rect 24268 9324 24274 9376
rect 25682 9324 25688 9376
rect 25740 9364 25746 9376
rect 25869 9367 25927 9373
rect 25869 9364 25881 9367
rect 25740 9336 25881 9364
rect 25740 9324 25746 9336
rect 25869 9333 25881 9336
rect 25915 9333 25927 9367
rect 27614 9364 27620 9376
rect 27575 9336 27620 9364
rect 25869 9327 25927 9333
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2130 9160 2136 9172
rect 2087 9132 2136 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 4062 9160 4068 9172
rect 3559 9132 4068 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4488 9132 4537 9160
rect 4488 9120 4494 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 4982 9120 4988 9172
rect 5040 9160 5046 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 5040 9132 5089 9160
rect 5040 9120 5046 9132
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5077 9123 5135 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5902 9160 5908 9172
rect 5863 9132 5908 9160
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 6914 9160 6920 9172
rect 6875 9132 6920 9160
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10836 9132 10885 9160
rect 10836 9120 10842 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 10873 9123 10931 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 16485 9163 16543 9169
rect 16485 9129 16497 9163
rect 16531 9160 16543 9163
rect 16850 9160 16856 9172
rect 16531 9132 16856 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17862 9160 17868 9172
rect 17775 9132 17868 9160
rect 17862 9120 17868 9132
rect 17920 9160 17926 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 17920 9132 19257 9160
rect 17920 9120 17926 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 19245 9123 19303 9129
rect 19705 9163 19763 9169
rect 19705 9129 19717 9163
rect 19751 9160 19763 9163
rect 19886 9160 19892 9172
rect 19751 9132 19892 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 20346 9160 20352 9172
rect 20307 9132 20352 9160
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 21542 9160 21548 9172
rect 21503 9132 21548 9160
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 22465 9163 22523 9169
rect 22465 9129 22477 9163
rect 22511 9160 22523 9163
rect 22830 9160 22836 9172
rect 22511 9132 22836 9160
rect 22511 9129 22523 9132
rect 22465 9123 22523 9129
rect 22830 9120 22836 9132
rect 22888 9160 22894 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22888 9132 23029 9160
rect 22888 9120 22894 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23017 9123 23075 9129
rect 24949 9163 25007 9169
rect 24949 9129 24961 9163
rect 24995 9160 25007 9163
rect 25682 9160 25688 9172
rect 24995 9132 25688 9160
rect 24995 9129 25007 9132
rect 24949 9123 25007 9129
rect 25682 9120 25688 9132
rect 25740 9120 25746 9172
rect 25958 9160 25964 9172
rect 25919 9132 25964 9160
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 2406 9092 2412 9104
rect 1412 9064 2412 9092
rect 1412 9033 1440 9064
rect 2406 9052 2412 9064
rect 2464 9052 2470 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 1397 8987 1455 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 9024 4491 9027
rect 4614 9024 4620 9036
rect 4479 8996 4620 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 7276 9027 7334 9033
rect 7276 9024 7288 9027
rect 6696 8996 7288 9024
rect 6696 8984 6702 8996
rect 7276 8993 7288 8996
rect 7322 9024 7334 9027
rect 8110 9024 8116 9036
rect 7322 8996 8116 9024
rect 7322 8993 7334 8996
rect 7276 8987 7334 8993
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10796 9024 10824 9120
rect 18782 9092 18788 9104
rect 18743 9064 18788 9092
rect 18782 9052 18788 9064
rect 18840 9052 18846 9104
rect 19613 9095 19671 9101
rect 19613 9061 19625 9095
rect 19659 9092 19671 9095
rect 20070 9092 20076 9104
rect 19659 9064 20076 9092
rect 19659 9061 19671 9064
rect 19613 9055 19671 9061
rect 20070 9052 20076 9064
rect 20128 9092 20134 9104
rect 21450 9092 21456 9104
rect 20128 9064 21456 9092
rect 20128 9052 20134 9064
rect 21450 9052 21456 9064
rect 21508 9052 21514 9104
rect 22738 9092 22744 9104
rect 22699 9064 22744 9092
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 23198 9052 23204 9104
rect 23256 9092 23262 9104
rect 23477 9095 23535 9101
rect 23477 9092 23489 9095
rect 23256 9064 23489 9092
rect 23256 9052 23262 9064
rect 23477 9061 23489 9064
rect 23523 9061 23535 9095
rect 23477 9055 23535 9061
rect 26418 9052 26424 9104
rect 26476 9092 26482 9104
rect 26970 9092 26976 9104
rect 26476 9064 26976 9092
rect 26476 9052 26482 9064
rect 26970 9052 26976 9064
rect 27028 9092 27034 9104
rect 27065 9095 27123 9101
rect 27065 9092 27077 9095
rect 27028 9064 27077 9092
rect 27028 9052 27034 9064
rect 27065 9061 27077 9064
rect 27111 9061 27123 9095
rect 27065 9055 27123 9061
rect 11790 9024 11796 9036
rect 10643 8996 10824 9024
rect 11751 8996 11796 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 17773 9027 17831 9033
rect 17773 8993 17785 9027
rect 17819 9024 17831 9027
rect 18230 9024 18236 9036
rect 17819 8996 18236 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 9024 18567 9027
rect 19150 9024 19156 9036
rect 18555 8996 19156 9024
rect 18555 8993 18567 8996
rect 18509 8987 18567 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 23382 9024 23388 9036
rect 23343 8996 23388 9024
rect 23382 8984 23388 8996
rect 23440 8984 23446 9036
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 24026 9024 24032 9036
rect 23900 8996 24032 9024
rect 23900 8984 23906 8996
rect 24026 8984 24032 8996
rect 24084 8984 24090 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 3476 8928 4721 8956
rect 3476 8916 3482 8928
rect 4709 8925 4721 8928
rect 4755 8956 4767 8959
rect 5442 8956 5448 8968
rect 4755 8928 5448 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6972 8928 7021 8956
rect 6972 8916 6978 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 11974 8956 11980 8968
rect 11931 8928 11980 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8956 12127 8959
rect 12434 8956 12440 8968
rect 12115 8928 12440 8956
rect 12115 8925 12127 8928
rect 12069 8919 12127 8925
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17460 8928 17969 8956
rect 17460 8916 17466 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19797 8959 19855 8965
rect 19797 8956 19809 8959
rect 19116 8928 19809 8956
rect 19116 8916 19122 8928
rect 19797 8925 19809 8928
rect 19843 8925 19855 8959
rect 23566 8956 23572 8968
rect 23527 8928 23572 8956
rect 19797 8919 19855 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9398 8820 9404 8832
rect 9079 8792 9404 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9398 8780 9404 8792
rect 9456 8820 9462 8832
rect 9674 8820 9680 8832
rect 9456 8792 9680 8820
rect 9456 8780 9462 8792
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10410 8820 10416 8832
rect 10371 8792 10416 8820
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 11204 8792 11437 8820
rect 11204 8780 11210 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 13998 8820 14004 8832
rect 13688 8792 14004 8820
rect 13688 8780 13694 8792
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 17000 8792 17417 8820
rect 17000 8780 17006 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 24118 8820 24124 8832
rect 24079 8792 24124 8820
rect 17405 8783 17463 8789
rect 24118 8780 24124 8792
rect 24176 8780 24182 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 6638 8616 6644 8628
rect 6599 8588 6644 8616
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 9122 8616 9128 8628
rect 8895 8588 9128 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18230 8616 18236 8628
rect 18191 8588 18236 8616
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 19116 8588 19257 8616
rect 19116 8576 19122 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 19245 8579 19303 8585
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 19886 8616 19892 8628
rect 19751 8588 19892 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20070 8616 20076 8628
rect 20031 8588 20076 8616
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27525 8619 27583 8625
rect 27525 8616 27537 8619
rect 26568 8588 27537 8616
rect 26568 8576 26574 8588
rect 27525 8585 27537 8588
rect 27571 8585 27583 8619
rect 27525 8579 27583 8585
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 1581 8551 1639 8557
rect 1581 8548 1593 8551
rect 1452 8520 1593 8548
rect 1452 8508 1458 8520
rect 1581 8517 1593 8520
rect 1627 8517 1639 8551
rect 1581 8511 1639 8517
rect 2222 8508 2228 8560
rect 2280 8548 2286 8560
rect 3418 8548 3424 8560
rect 2280 8520 3424 8548
rect 2280 8508 2286 8520
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 4430 8548 4436 8560
rect 4203 8520 4436 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 5442 8548 5448 8560
rect 4488 8520 5448 8548
rect 4488 8508 4494 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6914 8508 6920 8560
rect 6972 8548 6978 8560
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 6972 8520 7389 8548
rect 6972 8508 6978 8520
rect 7377 8517 7389 8520
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 10597 8551 10655 8557
rect 10597 8548 10609 8551
rect 9548 8520 10609 8548
rect 9548 8508 9554 8520
rect 10597 8517 10609 8520
rect 10643 8548 10655 8551
rect 10643 8520 11376 8548
rect 10643 8517 10655 8520
rect 10597 8511 10655 8517
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 2556 8452 2789 8480
rect 2556 8440 2562 8452
rect 2777 8449 2789 8452
rect 2823 8480 2835 8483
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 2823 8452 3801 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 3789 8449 3801 8452
rect 3835 8480 3847 8483
rect 4982 8480 4988 8492
rect 3835 8452 4988 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5132 8452 5917 8480
rect 5132 8440 5138 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7331 8452 7941 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 7929 8449 7941 8452
rect 7975 8480 7987 8483
rect 8386 8480 8392 8492
rect 7975 8452 8392 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 9582 8480 9588 8492
rect 8527 8452 9588 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 11146 8480 11152 8492
rect 11107 8452 11152 8480
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11348 8489 11376 8520
rect 16298 8508 16304 8560
rect 16356 8548 16362 8560
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 16356 8520 16405 8548
rect 16356 8508 16362 8520
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 22741 8551 22799 8557
rect 22741 8517 22753 8551
rect 22787 8548 22799 8551
rect 23566 8548 23572 8560
rect 22787 8520 23572 8548
rect 22787 8517 22799 8520
rect 22741 8511 22799 8517
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 26970 8548 26976 8560
rect 26931 8520 26976 8548
rect 26970 8508 26976 8520
rect 27028 8508 27034 8560
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11606 8480 11612 8492
rect 11379 8452 11612 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12526 8480 12532 8492
rect 12483 8452 12532 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16224 8452 16957 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 2038 8412 2044 8424
rect 1443 8384 2044 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 9180 8384 9321 8412
rect 9180 8372 9186 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 10229 8415 10287 8421
rect 9456 8384 9501 8412
rect 9456 8372 9462 8384
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 11057 8415 11115 8421
rect 11057 8412 11069 8415
rect 10275 8384 11069 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 11057 8381 11069 8384
rect 11103 8412 11115 8415
rect 12250 8412 12256 8424
rect 11103 8384 12256 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 16224 8356 16252 8452
rect 16945 8449 16957 8452
rect 16991 8480 17003 8483
rect 17862 8480 17868 8492
rect 16991 8452 17868 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 22646 8440 22652 8492
rect 22704 8480 22710 8492
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 22704 8452 23121 8480
rect 22704 8440 22710 8452
rect 23109 8449 23121 8452
rect 23155 8480 23167 8483
rect 23934 8480 23940 8492
rect 23155 8452 23940 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 24118 8440 24124 8492
rect 24176 8480 24182 8492
rect 24305 8483 24363 8489
rect 24305 8480 24317 8483
rect 24176 8452 24317 8480
rect 24176 8440 24182 8452
rect 24305 8449 24317 8452
rect 24351 8480 24363 8483
rect 24351 8452 24716 8480
rect 24351 8449 24363 8452
rect 24305 8443 24363 8449
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 16850 8412 16856 8424
rect 16807 8384 16856 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 23477 8415 23535 8421
rect 23477 8381 23489 8415
rect 23523 8412 23535 8415
rect 23523 8384 24164 8412
rect 23523 8381 23535 8384
rect 23477 8375 23535 8381
rect 4893 8347 4951 8353
rect 4893 8313 4905 8347
rect 4939 8344 4951 8347
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 4939 8316 5549 8344
rect 4939 8313 4951 8316
rect 4893 8307 4951 8313
rect 5537 8313 5549 8316
rect 5583 8344 5595 8347
rect 6086 8344 6092 8356
rect 5583 8316 6092 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 7156 8316 7757 8344
rect 7156 8304 7162 8316
rect 7745 8313 7757 8316
rect 7791 8344 7803 8347
rect 7791 8316 10732 8344
rect 7791 8313 7803 8316
rect 7745 8307 7803 8313
rect 4522 8276 4528 8288
rect 4483 8248 4528 8276
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8938 8276 8944 8288
rect 7892 8248 7937 8276
rect 8899 8248 8944 8276
rect 7892 8236 7898 8248
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 10704 8285 10732 8316
rect 11974 8304 11980 8356
rect 12032 8344 12038 8356
rect 12069 8347 12127 8353
rect 12069 8344 12081 8347
rect 12032 8316 12081 8344
rect 12032 8304 12038 8316
rect 12069 8313 12081 8316
rect 12115 8313 12127 8347
rect 16206 8344 16212 8356
rect 16167 8316 16212 8344
rect 12069 8307 12127 8313
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 16482 8304 16488 8356
rect 16540 8344 16546 8356
rect 16942 8344 16948 8356
rect 16540 8316 16948 8344
rect 16540 8304 16546 8316
rect 16868 8285 16896 8316
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 22373 8347 22431 8353
rect 22373 8313 22385 8347
rect 22419 8344 22431 8347
rect 22419 8316 23520 8344
rect 22419 8313 22431 8316
rect 22373 8307 22431 8313
rect 23492 8288 23520 8316
rect 23934 8304 23940 8356
rect 23992 8344 23998 8356
rect 24136 8353 24164 8384
rect 24688 8356 24716 8452
rect 25590 8412 25596 8424
rect 25551 8384 25596 8412
rect 25590 8372 25596 8384
rect 25648 8372 25654 8424
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23992 8316 24041 8344
rect 23992 8304 23998 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 24029 8307 24087 8313
rect 24121 8347 24179 8353
rect 24121 8313 24133 8347
rect 24167 8344 24179 8347
rect 24578 8344 24584 8356
rect 24167 8316 24584 8344
rect 24167 8313 24179 8316
rect 24121 8307 24179 8313
rect 24578 8304 24584 8316
rect 24636 8304 24642 8356
rect 24670 8304 24676 8356
rect 24728 8344 24734 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 24728 8316 25421 8344
rect 24728 8304 24734 8316
rect 25409 8313 25421 8316
rect 25455 8344 25467 8347
rect 25838 8347 25896 8353
rect 25838 8344 25850 8347
rect 25455 8316 25850 8344
rect 25455 8313 25467 8316
rect 25409 8307 25467 8313
rect 25838 8313 25850 8316
rect 25884 8313 25896 8347
rect 25838 8307 25896 8313
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8245 10747 8279
rect 10689 8239 10747 8245
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8245 16911 8279
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 16853 8239 16911 8245
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 23474 8236 23480 8288
rect 23532 8236 23538 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2225 8035 2283 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 4982 8072 4988 8084
rect 4943 8044 4988 8072
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 6086 8072 6092 8084
rect 6047 8044 6092 8072
rect 6086 8032 6092 8044
rect 6144 8032 6150 8084
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 7834 8072 7840 8084
rect 7791 8044 7840 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 7834 8032 7840 8044
rect 7892 8072 7898 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7892 8044 8033 8072
rect 7892 8032 7898 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8478 8072 8484 8084
rect 8391 8044 8484 8072
rect 8021 8035 8079 8041
rect 8478 8032 8484 8044
rect 8536 8072 8542 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 8536 8044 9689 8072
rect 8536 8032 8542 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9916 8044 10057 8072
rect 9916 8032 9922 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 10045 8035 10103 8041
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 12434 8072 12440 8084
rect 11563 8044 12440 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 4890 8004 4896 8016
rect 4851 7976 4896 8004
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 8938 8004 8944 8016
rect 8435 7976 8944 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 8938 7964 8944 7976
rect 8996 7964 9002 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1670 7936 1676 7948
rect 1443 7908 1676 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 7340 7908 7389 7936
rect 7340 7896 7346 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10594 7936 10600 7948
rect 10183 7908 10600 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5132 7840 5177 7868
rect 5132 7828 5138 7840
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 8168 7840 8677 7868
rect 8168 7828 8174 7840
rect 8665 7837 8677 7840
rect 8711 7868 8723 7871
rect 9490 7868 9496 7880
rect 8711 7840 9496 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 9640 7840 10333 7868
rect 9640 7828 9646 7840
rect 10321 7837 10333 7840
rect 10367 7868 10379 7871
rect 11532 7868 11560 8035
rect 12434 8032 12440 8044
rect 12492 8072 12498 8084
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12492 8044 13461 8072
rect 12492 8032 12498 8044
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14792 8044 14841 8072
rect 14792 8032 14798 8044
rect 14829 8041 14841 8044
rect 14875 8072 14887 8075
rect 15010 8072 15016 8084
rect 14875 8044 15016 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 18012 8044 18061 8072
rect 18012 8032 18018 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 18049 8035 18107 8041
rect 20070 8032 20076 8084
rect 20128 8072 20134 8084
rect 21361 8075 21419 8081
rect 21361 8072 21373 8075
rect 20128 8044 21373 8072
rect 20128 8032 20134 8044
rect 21361 8041 21373 8044
rect 21407 8041 21419 8075
rect 21361 8035 21419 8041
rect 23109 8075 23167 8081
rect 23109 8041 23121 8075
rect 23155 8072 23167 8075
rect 23198 8072 23204 8084
rect 23155 8044 23204 8072
rect 23155 8041 23167 8044
rect 23109 8035 23167 8041
rect 23198 8032 23204 8044
rect 23256 8072 23262 8084
rect 23569 8075 23627 8081
rect 23569 8072 23581 8075
rect 23256 8044 23581 8072
rect 23256 8032 23262 8044
rect 23569 8041 23581 8044
rect 23615 8041 23627 8075
rect 23569 8035 23627 8041
rect 24762 8032 24768 8084
rect 24820 8072 24826 8084
rect 25590 8072 25596 8084
rect 24820 8044 25596 8072
rect 24820 8032 24826 8044
rect 25590 8032 25596 8044
rect 25648 8032 25654 8084
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 12618 8004 12624 8016
rect 12084 7976 12624 8004
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12084 7945 12112 7976
rect 12618 7964 12624 7976
rect 12676 8004 12682 8016
rect 13630 8004 13636 8016
rect 12676 7976 13636 8004
rect 12676 7964 12682 7976
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 12342 7945 12348 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11940 7908 12081 7936
rect 11940 7896 11946 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12336 7936 12348 7945
rect 12303 7908 12348 7936
rect 12069 7899 12127 7905
rect 12336 7899 12348 7908
rect 12342 7896 12348 7899
rect 12400 7896 12406 7948
rect 16666 7936 16672 7948
rect 16627 7908 16672 7936
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 16758 7896 16764 7948
rect 16816 7936 16822 7948
rect 16925 7939 16983 7945
rect 16925 7936 16937 7939
rect 16816 7908 16937 7936
rect 16816 7896 16822 7908
rect 16925 7905 16937 7908
rect 16971 7936 16983 7939
rect 17402 7936 17408 7948
rect 16971 7908 17408 7936
rect 16971 7905 16983 7908
rect 16925 7899 16983 7905
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 20438 7896 20444 7948
rect 20496 7936 20502 7948
rect 21266 7936 21272 7948
rect 20496 7908 21272 7936
rect 20496 7896 20502 7908
rect 21266 7896 21272 7908
rect 21324 7896 21330 7948
rect 23106 7896 23112 7948
rect 23164 7936 23170 7948
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23164 7908 23949 7936
rect 23164 7896 23170 7908
rect 23937 7905 23949 7908
rect 23983 7905 23995 7939
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 23937 7899 23995 7905
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 19794 7868 19800 7880
rect 10367 7840 11560 7868
rect 19755 7840 19800 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 21450 7868 21456 7880
rect 21411 7840 21456 7868
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 23290 7828 23296 7880
rect 23348 7868 23354 7880
rect 23842 7868 23848 7880
rect 23348 7840 23848 7868
rect 23348 7828 23354 7840
rect 23842 7828 23848 7840
rect 23900 7868 23906 7880
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 23900 7840 24041 7868
rect 23900 7828 23906 7840
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7868 24271 7871
rect 24670 7868 24676 7880
rect 24259 7840 24676 7868
rect 24259 7837 24271 7840
rect 24213 7831 24271 7837
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 4341 7803 4399 7809
rect 4341 7769 4353 7803
rect 4387 7800 4399 7803
rect 4614 7800 4620 7812
rect 4387 7772 4620 7800
rect 4387 7769 4399 7772
rect 4341 7763 4399 7769
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7193 7803 7251 7809
rect 7193 7800 7205 7803
rect 7064 7772 7205 7800
rect 7064 7760 7070 7772
rect 7193 7769 7205 7772
rect 7239 7769 7251 7803
rect 7193 7763 7251 7769
rect 19518 7760 19524 7812
rect 19576 7800 19582 7812
rect 20901 7803 20959 7809
rect 20901 7800 20913 7803
rect 19576 7772 20913 7800
rect 19576 7760 19582 7772
rect 20901 7769 20913 7772
rect 20947 7769 20959 7803
rect 20901 7763 20959 7769
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 5166 7732 5172 7744
rect 4571 7704 5172 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 5166 7692 5172 7704
rect 5224 7732 5230 7744
rect 5537 7735 5595 7741
rect 5537 7732 5549 7735
rect 5224 7704 5549 7732
rect 5224 7692 5230 7704
rect 5537 7701 5549 7704
rect 5583 7701 5595 7735
rect 19150 7732 19156 7744
rect 19111 7704 19156 7732
rect 5537 7695 5595 7701
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 20346 7692 20352 7744
rect 20404 7732 20410 7744
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 20404 7704 20637 7732
rect 20404 7692 20410 7704
rect 20625 7701 20637 7704
rect 20671 7701 20683 7735
rect 20625 7695 20683 7701
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21542 7732 21548 7744
rect 20864 7704 21548 7732
rect 20864 7692 20870 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2498 7528 2504 7540
rect 2179 7500 2504 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 4246 7528 4252 7540
rect 4159 7500 4252 7528
rect 4246 7488 4252 7500
rect 4304 7528 4310 7540
rect 4982 7528 4988 7540
rect 4304 7500 4988 7528
rect 4304 7488 4310 7500
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 7282 7528 7288 7540
rect 7243 7500 7288 7528
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8478 7528 8484 7540
rect 8439 7500 8484 7528
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 8849 7531 8907 7537
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 8938 7528 8944 7540
rect 8895 7500 8944 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9582 7528 9588 7540
rect 9447 7500 9588 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 9858 7528 9864 7540
rect 9815 7500 9864 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10502 7528 10508 7540
rect 10463 7500 10508 7528
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 16758 7528 16764 7540
rect 16719 7500 16764 7528
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 20070 7528 20076 7540
rect 20031 7500 20076 7528
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 21652 7500 22569 7528
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 4890 7460 4896 7472
rect 4663 7432 4896 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 17037 7463 17095 7469
rect 17037 7460 17049 7463
rect 16724 7432 17049 7460
rect 16724 7420 16730 7432
rect 17037 7429 17049 7432
rect 17083 7429 17095 7463
rect 17037 7423 17095 7429
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 2188 7364 2237 7392
rect 2188 7352 2194 7364
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 2225 7355 2283 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5316 7364 5733 7392
rect 5316 7352 5322 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10183 7364 11161 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 11149 7361 11161 7364
rect 11195 7392 11207 7395
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 11195 7364 12081 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 12069 7361 12081 7364
rect 12115 7392 12127 7395
rect 12342 7392 12348 7404
rect 12115 7364 12348 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 12342 7352 12348 7364
rect 12400 7392 12406 7404
rect 12434 7392 12440 7404
rect 12400 7364 12440 7392
rect 12400 7352 12406 7364
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 14734 7392 14740 7404
rect 14695 7364 14740 7392
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19659 7364 20760 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 4580 7296 5089 7324
rect 4580 7284 4586 7296
rect 5077 7293 5089 7296
rect 5123 7324 5135 7327
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5123 7296 6101 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10560 7296 11069 7324
rect 10560 7284 10566 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19628 7324 19656 7355
rect 19015 7296 19656 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 20346 7284 20352 7336
rect 20404 7324 20410 7336
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 20404 7296 20637 7324
rect 20404 7284 20410 7296
rect 20625 7293 20637 7296
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 2498 7265 2504 7268
rect 2492 7256 2504 7265
rect 2459 7228 2504 7256
rect 2492 7219 2504 7228
rect 2498 7216 2504 7219
rect 2556 7216 2562 7268
rect 10318 7216 10324 7268
rect 10376 7256 10382 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 10376 7228 10977 7256
rect 10376 7216 10382 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 10965 7219 11023 7225
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 14332 7228 14657 7256
rect 14332 7216 14338 7228
rect 14645 7225 14657 7228
rect 14691 7256 14703 7259
rect 15004 7259 15062 7265
rect 15004 7256 15016 7259
rect 14691 7228 15016 7256
rect 14691 7225 14703 7228
rect 14645 7219 14703 7225
rect 15004 7225 15016 7228
rect 15050 7256 15062 7259
rect 15102 7256 15108 7268
rect 15050 7228 15108 7256
rect 15050 7225 15062 7228
rect 15004 7219 15062 7225
rect 15102 7216 15108 7228
rect 15160 7216 15166 7268
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19429 7259 19487 7265
rect 19429 7256 19441 7259
rect 19208 7228 19441 7256
rect 19208 7216 19214 7228
rect 19429 7225 19441 7228
rect 19475 7256 19487 7259
rect 19475 7228 20668 7256
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 20640 7200 20668 7228
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 10594 7188 10600 7200
rect 10555 7160 10600 7188
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 19061 7191 19119 7197
rect 19061 7157 19073 7191
rect 19107 7188 19119 7191
rect 19242 7188 19248 7200
rect 19107 7160 19248 7188
rect 19107 7157 19119 7160
rect 19061 7151 19119 7157
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 20438 7188 20444 7200
rect 20399 7160 20444 7188
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20622 7148 20628 7200
rect 20680 7148 20686 7200
rect 20732 7188 20760 7364
rect 21652 7324 21680 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 23106 7528 23112 7540
rect 23067 7500 23112 7528
rect 22557 7491 22615 7497
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 23474 7488 23480 7540
rect 23532 7528 23538 7540
rect 23661 7531 23719 7537
rect 23661 7528 23673 7531
rect 23532 7500 23673 7528
rect 23532 7488 23538 7500
rect 23661 7497 23673 7500
rect 23707 7497 23719 7531
rect 26602 7528 26608 7540
rect 26563 7500 26608 7528
rect 23661 7491 23719 7497
rect 26602 7488 26608 7500
rect 26660 7488 26666 7540
rect 26510 7420 26516 7472
rect 26568 7460 26574 7472
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26568 7432 27353 7460
rect 26568 7420 26574 7432
rect 27341 7429 27353 7432
rect 27387 7429 27399 7463
rect 27706 7460 27712 7472
rect 27667 7432 27712 7460
rect 27341 7423 27399 7429
rect 27706 7420 27712 7432
rect 27764 7420 27770 7472
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7392 24363 7395
rect 24670 7392 24676 7404
rect 24351 7364 24676 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 24670 7352 24676 7364
rect 24728 7352 24734 7404
rect 24026 7324 24032 7336
rect 21376 7296 21680 7324
rect 23987 7296 24032 7324
rect 21376 7268 21404 7296
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 26418 7284 26424 7296
rect 26476 7324 26482 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26476 7296 26985 7324
rect 26476 7284 26482 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 27522 7324 27528 7336
rect 27483 7296 27528 7324
rect 26973 7287 27031 7293
rect 27522 7284 27528 7296
rect 27580 7324 27586 7336
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27580 7296 28089 7324
rect 27580 7284 27586 7296
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 20892 7259 20950 7265
rect 20892 7225 20904 7259
rect 20938 7256 20950 7259
rect 21358 7256 21364 7268
rect 20938 7228 21364 7256
rect 20938 7225 20950 7228
rect 20892 7219 20950 7225
rect 21358 7216 21364 7228
rect 21416 7216 21422 7268
rect 23477 7259 23535 7265
rect 23477 7225 23489 7259
rect 23523 7256 23535 7259
rect 23842 7256 23848 7268
rect 23523 7228 23848 7256
rect 23523 7225 23535 7228
rect 23477 7219 23535 7225
rect 23842 7216 23848 7228
rect 23900 7256 23906 7268
rect 25130 7256 25136 7268
rect 23900 7228 25136 7256
rect 23900 7216 23906 7228
rect 25130 7216 25136 7228
rect 25188 7216 25194 7268
rect 21450 7188 21456 7200
rect 20732 7160 21456 7188
rect 21450 7148 21456 7160
rect 21508 7188 21514 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 21508 7160 22017 7188
rect 21508 7148 21514 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 22005 7151 22063 7157
rect 23750 7148 23756 7200
rect 23808 7188 23814 7200
rect 24121 7191 24179 7197
rect 24121 7188 24133 7191
rect 23808 7160 24133 7188
rect 23808 7148 23814 7160
rect 24121 7157 24133 7160
rect 24167 7157 24179 7191
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24121 7151 24179 7157
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 2317 6987 2375 6993
rect 2317 6953 2329 6987
rect 2363 6984 2375 6987
rect 2498 6984 2504 6996
rect 2363 6956 2504 6984
rect 2363 6953 2375 6956
rect 2317 6947 2375 6953
rect 2498 6944 2504 6956
rect 2556 6984 2562 6996
rect 5074 6984 5080 6996
rect 2556 6956 5080 6984
rect 2556 6944 2562 6956
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 9953 6987 10011 6993
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10594 6984 10600 6996
rect 9999 6956 10600 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 15654 6984 15660 6996
rect 15615 6956 15660 6984
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 19794 6944 19800 6996
rect 19852 6984 19858 6996
rect 21266 6984 21272 6996
rect 19852 6956 21272 6984
rect 19852 6944 19858 6956
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 24026 6984 24032 6996
rect 23987 6956 24032 6984
rect 24026 6944 24032 6956
rect 24084 6944 24090 6996
rect 7006 6916 7012 6928
rect 5000 6888 5304 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1854 6848 1860 6860
rect 1443 6820 1860 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5000 6848 5028 6888
rect 5166 6857 5172 6860
rect 5160 6848 5172 6857
rect 4939 6820 5028 6848
rect 5127 6820 5172 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 5160 6811 5172 6820
rect 5166 6808 5172 6811
rect 5224 6808 5230 6860
rect 5276 6848 5304 6888
rect 6840 6888 7012 6916
rect 5534 6848 5540 6860
rect 5276 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6848 5598 6860
rect 6840 6848 6868 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 19518 6916 19524 6928
rect 15304 6888 15792 6916
rect 5592 6820 6868 6848
rect 5592 6808 5598 6820
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10376 6820 10609 6848
rect 10376 6808 10382 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 13998 6848 14004 6860
rect 13959 6820 14004 6848
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14182 6848 14188 6860
rect 14108 6820 14188 6848
rect 13648 6780 13676 6808
rect 14108 6789 14136 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 15304 6792 15332 6888
rect 15764 6848 15792 6888
rect 19352 6888 19524 6916
rect 16114 6848 16120 6860
rect 15764 6820 16120 6848
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13648 6752 14105 6780
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 14093 6743 14151 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6780 14795 6783
rect 15286 6780 15292 6792
rect 14783 6752 15292 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 15746 6780 15752 6792
rect 15707 6752 15752 6780
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15856 6789 15884 6820
rect 16114 6808 16120 6820
rect 16172 6848 16178 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 16172 6820 16405 6848
rect 16172 6808 16178 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 17310 6848 17316 6860
rect 17271 6820 17316 6848
rect 16393 6811 16451 6817
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 13633 6715 13691 6721
rect 13633 6681 13645 6715
rect 13679 6712 13691 6715
rect 16408 6712 16436 6811
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 19153 6851 19211 6857
rect 19153 6817 19165 6851
rect 19199 6848 19211 6851
rect 19352 6848 19380 6888
rect 19518 6876 19524 6888
rect 19576 6876 19582 6928
rect 21358 6876 21364 6928
rect 21416 6876 21422 6928
rect 19199 6820 19380 6848
rect 20717 6851 20775 6857
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 20717 6817 20729 6851
rect 20763 6848 20775 6851
rect 21174 6848 21180 6860
rect 20763 6820 21180 6848
rect 20763 6817 20775 6820
rect 20717 6811 20775 6817
rect 21174 6808 21180 6820
rect 21232 6848 21238 6860
rect 21376 6848 21404 6876
rect 21232 6820 21496 6848
rect 21232 6808 21238 6820
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 21468 6789 21496 6820
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 26513 6851 26571 6857
rect 26513 6848 26525 6851
rect 26384 6820 26525 6848
rect 26384 6808 26390 6820
rect 26513 6817 26525 6820
rect 26559 6848 26571 6851
rect 27338 6848 27344 6860
rect 26559 6820 27344 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 27338 6808 27344 6820
rect 27396 6808 27402 6860
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 17276 6752 17417 6780
rect 17276 6740 17282 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 17512 6712 17540 6743
rect 17678 6712 17684 6724
rect 13679 6684 15700 6712
rect 16408 6684 17684 6712
rect 13679 6681 13691 6684
rect 13633 6675 13691 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5074 6644 5080 6656
rect 4663 6616 5080 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5074 6604 5080 6616
rect 5132 6644 5138 6656
rect 5258 6644 5264 6656
rect 5132 6616 5264 6644
rect 5132 6604 5138 6616
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 8849 6647 8907 6653
rect 8849 6613 8861 6647
rect 8895 6644 8907 6647
rect 9306 6644 9312 6656
rect 8895 6616 9312 6644
rect 8895 6613 8907 6616
rect 8849 6607 8907 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 15068 6616 15301 6644
rect 15068 6604 15074 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15672 6644 15700 6684
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 20901 6715 20959 6721
rect 20901 6712 20913 6715
rect 20772 6684 20913 6712
rect 20772 6672 20778 6684
rect 20901 6681 20913 6684
rect 20947 6681 20959 6715
rect 20901 6675 20959 6681
rect 20990 6672 20996 6724
rect 21048 6712 21054 6724
rect 21376 6712 21404 6743
rect 21818 6712 21824 6724
rect 21048 6684 21824 6712
rect 21048 6672 21054 6684
rect 21818 6672 21824 6684
rect 21876 6672 21882 6724
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 15746 6644 15752 6656
rect 15672 6616 15752 6644
rect 15289 6607 15347 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 23750 6644 23756 6656
rect 23711 6616 23756 6644
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 24489 6647 24547 6653
rect 24489 6613 24501 6647
rect 24535 6644 24547 6647
rect 24670 6644 24676 6656
rect 24535 6616 24676 6644
rect 24535 6613 24547 6616
rect 24489 6607 24547 6613
rect 24670 6604 24676 6616
rect 24728 6644 24734 6656
rect 25314 6644 25320 6656
rect 24728 6616 25320 6644
rect 24728 6604 24734 6616
rect 25314 6604 25320 6616
rect 25372 6604 25378 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1854 6440 1860 6452
rect 1719 6412 1860 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 14274 6440 14280 6452
rect 13403 6412 14280 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 15654 6440 15660 6452
rect 15615 6412 15660 6440
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17368 6412 17785 6440
rect 17368 6400 17374 6412
rect 17773 6409 17785 6412
rect 17819 6440 17831 6443
rect 20990 6440 20996 6452
rect 17819 6412 18092 6440
rect 20951 6412 20996 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 5077 6375 5135 6381
rect 5077 6372 5089 6375
rect 3620 6344 5089 6372
rect 3620 6316 3648 6344
rect 5077 6341 5089 6344
rect 5123 6372 5135 6375
rect 5166 6372 5172 6384
rect 5123 6344 5172 6372
rect 5123 6341 5135 6344
rect 5077 6335 5135 6341
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10321 6375 10379 6381
rect 10321 6372 10333 6375
rect 9732 6344 10333 6372
rect 9732 6332 9738 6344
rect 10321 6341 10333 6344
rect 10367 6341 10379 6375
rect 10321 6335 10379 6341
rect 17218 6332 17224 6384
rect 17276 6372 17282 6384
rect 17405 6375 17463 6381
rect 17405 6372 17417 6375
rect 17276 6344 17417 6372
rect 17276 6332 17282 6344
rect 17405 6341 17417 6344
rect 17451 6341 17463 6375
rect 17405 6335 17463 6341
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2363 6276 2973 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2961 6273 2973 6276
rect 3007 6304 3019 6307
rect 3602 6304 3608 6316
rect 3007 6276 3608 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4019 6276 4629 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4617 6273 4629 6276
rect 4663 6304 4675 6307
rect 6270 6304 6276 6316
rect 4663 6276 6276 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 9306 6304 9312 6316
rect 9267 6276 9312 6304
rect 9306 6264 9312 6276
rect 9364 6304 9370 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9364 6276 9781 6304
rect 9364 6264 9370 6276
rect 9769 6273 9781 6276
rect 9815 6304 9827 6307
rect 10502 6304 10508 6316
rect 9815 6276 10508 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 10502 6264 10508 6276
rect 10560 6304 10566 6316
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10560 6276 10885 6304
rect 10560 6264 10566 6276
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 15102 6304 15108 6316
rect 14599 6276 15108 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 2832 6208 3433 6236
rect 2832 6196 2838 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3421 6199 3479 6205
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4706 6236 4712 6248
rect 4479 6208 4712 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 8662 6236 8668 6248
rect 8575 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6236 8726 6248
rect 9122 6236 9128 6248
rect 8720 6208 9128 6236
rect 8720 6196 8726 6208
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 15028 6245 15056 6276
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15286 6304 15292 6316
rect 15247 6276 15292 6304
rect 15286 6264 15292 6276
rect 15344 6304 15350 6316
rect 18064 6313 18092 6412
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21266 6440 21272 6452
rect 21227 6412 21272 6440
rect 21266 6400 21272 6412
rect 21324 6400 21330 6452
rect 25314 6440 25320 6452
rect 25275 6412 25320 6440
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 27065 6443 27123 6449
rect 27065 6409 27077 6443
rect 27111 6440 27123 6443
rect 27154 6440 27160 6452
rect 27111 6412 27160 6440
rect 27111 6409 27123 6412
rect 27065 6403 27123 6409
rect 26602 6372 26608 6384
rect 26563 6344 26608 6372
rect 26602 6332 26608 6344
rect 26660 6332 26666 6384
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 15344 6276 16957 6304
rect 15344 6264 15350 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 10376 6208 10701 6236
rect 10376 6196 10382 6208
rect 10689 6205 10701 6208
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 16850 6236 16856 6248
rect 16811 6208 16856 6236
rect 15013 6199 15071 6205
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 22922 6196 22928 6248
rect 22980 6236 22986 6248
rect 23109 6239 23167 6245
rect 23109 6236 23121 6239
rect 22980 6208 23121 6236
rect 22980 6196 22986 6208
rect 23109 6205 23121 6208
rect 23155 6236 23167 6239
rect 23937 6239 23995 6245
rect 23937 6236 23949 6239
rect 23155 6208 23949 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 23937 6205 23949 6208
rect 23983 6236 23995 6239
rect 24762 6236 24768 6248
rect 23983 6208 24768 6236
rect 23983 6205 23995 6208
rect 23937 6199 23995 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6236 26479 6239
rect 27080 6236 27108 6403
rect 27154 6400 27160 6412
rect 27212 6400 27218 6452
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 26467 6208 27108 6236
rect 26467 6205 26479 6208
rect 26421 6199 26479 6205
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 9217 6171 9275 6177
rect 9217 6168 9229 6171
rect 8904 6140 9229 6168
rect 8904 6128 8910 6140
rect 9217 6137 9229 6140
rect 9263 6137 9275 6171
rect 9217 6131 9275 6137
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10781 6171 10839 6177
rect 10781 6168 10793 6171
rect 10192 6140 10793 6168
rect 10192 6128 10198 6140
rect 10781 6137 10793 6140
rect 10827 6137 10839 6171
rect 10781 6131 10839 6137
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 15105 6171 15163 6177
rect 15105 6168 15117 6171
rect 14608 6140 15117 6168
rect 14608 6128 14614 6140
rect 15105 6137 15117 6140
rect 15151 6137 15163 6171
rect 15105 6131 15163 6137
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16758 6168 16764 6180
rect 16347 6140 16764 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 24182 6171 24240 6177
rect 24182 6168 24194 6171
rect 23492 6140 24194 6168
rect 23492 6112 23520 6140
rect 24182 6137 24194 6140
rect 24228 6137 24240 6171
rect 24182 6131 24240 6137
rect 2406 6100 2412 6112
rect 2367 6072 2412 6100
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2740 6072 2881 6100
rect 2740 6060 2746 6072
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 2869 6063 2927 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4246 6060 4252 6112
rect 4304 6100 4310 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4304 6072 4537 6100
rect 4304 6060 4310 6072
rect 4525 6069 4537 6072
rect 4571 6069 4583 6103
rect 7742 6100 7748 6112
rect 7703 6072 7748 6100
rect 4525 6063 4583 6069
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8754 6100 8760 6112
rect 8715 6072 8760 6100
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 13630 6100 13636 6112
rect 13591 6072 13636 6100
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13998 6100 14004 6112
rect 13959 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14642 6100 14648 6112
rect 14603 6072 14648 6100
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 21637 6103 21695 6109
rect 21637 6100 21649 6103
rect 21324 6072 21649 6100
rect 21324 6060 21330 6072
rect 21637 6069 21649 6072
rect 21683 6069 21695 6103
rect 23474 6100 23480 6112
rect 23435 6072 23480 6100
rect 21637 6063 21695 6069
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 2774 5896 2780 5908
rect 2271 5868 2780 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 3329 5899 3387 5905
rect 3329 5896 3341 5899
rect 2924 5868 3341 5896
rect 2924 5856 2930 5868
rect 3329 5865 3341 5868
rect 3375 5896 3387 5899
rect 3786 5896 3792 5908
rect 3375 5868 3792 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 10318 5896 10324 5908
rect 10279 5868 10324 5896
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12492 5868 12817 5896
rect 12492 5856 12498 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 15841 5899 15899 5905
rect 15841 5896 15853 5899
rect 15804 5868 15853 5896
rect 15804 5856 15810 5868
rect 15841 5865 15853 5868
rect 15887 5865 15899 5899
rect 15841 5859 15899 5865
rect 16485 5899 16543 5905
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16850 5896 16856 5908
rect 16531 5868 16856 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 17000 5868 17049 5896
rect 17000 5856 17006 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17037 5859 17095 5865
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 19702 5896 19708 5908
rect 19615 5868 19708 5896
rect 19702 5856 19708 5868
rect 19760 5896 19766 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 19760 5868 20913 5896
rect 19760 5856 19766 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23532 5868 23857 5896
rect 23532 5856 23538 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 2590 5828 2596 5840
rect 2551 5800 2596 5828
rect 2590 5788 2596 5800
rect 2648 5788 2654 5840
rect 6270 5837 6276 5840
rect 6264 5828 6276 5837
rect 6231 5800 6276 5828
rect 6264 5791 6276 5800
rect 6270 5788 6276 5791
rect 6328 5788 6334 5840
rect 11882 5828 11888 5840
rect 11440 5800 11888 5828
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2464 5732 2820 5760
rect 2464 5720 2470 5732
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2498 5692 2504 5704
rect 2179 5664 2504 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2498 5652 2504 5664
rect 2556 5692 2562 5704
rect 2792 5701 2820 5732
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 11440 5769 11468 5800
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 17126 5828 17132 5840
rect 16448 5800 17132 5828
rect 16448 5788 16454 5800
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 19334 5788 19340 5840
rect 19392 5828 19398 5840
rect 19613 5831 19671 5837
rect 19613 5828 19625 5831
rect 19392 5800 19625 5828
rect 19392 5788 19398 5800
rect 19613 5797 19625 5800
rect 19659 5797 19671 5831
rect 22710 5831 22768 5837
rect 22710 5828 22722 5831
rect 19613 5791 19671 5797
rect 22112 5800 22722 5828
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5592 5732 6009 5760
rect 5592 5720 5598 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 11681 5763 11739 5769
rect 11681 5760 11693 5763
rect 11572 5732 11693 5760
rect 11572 5720 11578 5732
rect 11681 5729 11693 5732
rect 11727 5729 11739 5763
rect 11681 5723 11739 5729
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20772 5732 21281 5760
rect 20772 5720 20778 5732
rect 21269 5729 21281 5732
rect 21315 5760 21327 5763
rect 21910 5760 21916 5772
rect 21315 5732 21916 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 2685 5695 2743 5701
rect 2685 5692 2697 5695
rect 2556 5664 2697 5692
rect 2556 5652 2562 5664
rect 2685 5661 2697 5664
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16816 5664 17233 5692
rect 16816 5652 16822 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 19886 5692 19892 5704
rect 19847 5664 19892 5692
rect 17221 5655 17279 5661
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 21358 5692 21364 5704
rect 21319 5664 21364 5692
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21450 5652 21456 5704
rect 21508 5692 21514 5704
rect 22112 5692 22140 5800
rect 22710 5797 22722 5800
rect 22756 5797 22768 5831
rect 22710 5791 22768 5797
rect 22922 5788 22928 5840
rect 22980 5788 22986 5840
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 22940 5760 22968 5788
rect 22511 5732 22968 5760
rect 26513 5763 26571 5769
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 26786 5760 26792 5772
rect 26559 5732 26792 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 26786 5720 26792 5732
rect 26844 5720 26850 5772
rect 21508 5664 22140 5692
rect 21508 5652 21514 5664
rect 8846 5624 8852 5636
rect 8807 5596 8852 5624
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 26694 5624 26700 5636
rect 26655 5596 26700 5624
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 7374 5556 7380 5568
rect 7335 5528 7380 5556
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14645 5559 14703 5565
rect 14645 5556 14657 5559
rect 14608 5528 14657 5556
rect 14608 5516 14614 5528
rect 14645 5525 14657 5528
rect 14691 5525 14703 5559
rect 14645 5519 14703 5525
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 15286 5556 15292 5568
rect 14976 5528 15292 5556
rect 14976 5516 14982 5528
rect 15286 5516 15292 5528
rect 15344 5556 15350 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 15344 5528 15485 5556
rect 15344 5516 15350 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 16666 5556 16672 5568
rect 16627 5528 16672 5556
rect 15473 5519 15531 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 21266 5556 21272 5568
rect 20763 5528 21272 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 4706 5352 4712 5364
rect 4667 5324 4712 5352
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 6089 5355 6147 5361
rect 6089 5321 6101 5355
rect 6135 5352 6147 5355
rect 6270 5352 6276 5364
rect 6135 5324 6276 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 11882 5352 11888 5364
rect 11843 5324 11888 5352
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15160 5324 15577 5352
rect 15160 5312 15166 5324
rect 15565 5321 15577 5324
rect 15611 5352 15623 5355
rect 16758 5352 16764 5364
rect 15611 5324 16764 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17000 5324 17417 5352
rect 17000 5312 17006 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 17405 5315 17463 5321
rect 18969 5355 19027 5361
rect 18969 5321 18981 5355
rect 19015 5352 19027 5355
rect 19150 5352 19156 5364
rect 19015 5324 19156 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 20254 5312 20260 5364
rect 20312 5352 20318 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 20312 5324 20453 5352
rect 20312 5312 20318 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 20625 5355 20683 5361
rect 20625 5321 20637 5355
rect 20671 5352 20683 5355
rect 20714 5352 20720 5364
rect 20671 5324 20720 5352
rect 20671 5321 20683 5324
rect 20625 5315 20683 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21637 5355 21695 5361
rect 21637 5352 21649 5355
rect 21508 5324 21649 5352
rect 21508 5312 21514 5324
rect 21637 5321 21649 5324
rect 21683 5321 21695 5355
rect 21637 5315 21695 5321
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 2590 5284 2596 5296
rect 2363 5256 2596 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 5592 5256 6377 5284
rect 5592 5244 5598 5256
rect 6365 5253 6377 5256
rect 6411 5284 6423 5287
rect 6730 5284 6736 5296
rect 6411 5256 6736 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 8481 5287 8539 5293
rect 8481 5253 8493 5287
rect 8527 5284 8539 5287
rect 17126 5284 17132 5296
rect 8527 5256 9260 5284
rect 17087 5256 17132 5284
rect 8527 5253 8539 5256
rect 8481 5247 8539 5253
rect 9232 5228 9260 5256
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 19337 5287 19395 5293
rect 19337 5253 19349 5287
rect 19383 5284 19395 5287
rect 19886 5284 19892 5296
rect 19383 5256 19892 5284
rect 19383 5253 19395 5256
rect 19337 5247 19395 5253
rect 19886 5244 19892 5256
rect 19944 5244 19950 5296
rect 21652 5284 21680 5315
rect 21910 5312 21916 5364
rect 21968 5352 21974 5364
rect 22097 5355 22155 5361
rect 22097 5352 22109 5355
rect 21968 5324 22109 5352
rect 21968 5312 21974 5324
rect 22097 5321 22109 5324
rect 22143 5321 22155 5355
rect 22922 5352 22928 5364
rect 22883 5324 22928 5352
rect 22097 5315 22155 5321
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 26786 5312 26792 5364
rect 26844 5352 26850 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26844 5324 27353 5352
rect 26844 5312 26850 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 27341 5315 27399 5321
rect 22465 5287 22523 5293
rect 22465 5284 22477 5287
rect 21652 5256 22477 5284
rect 22465 5253 22477 5256
rect 22511 5253 22523 5287
rect 22465 5247 22523 5253
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3694 5216 3700 5228
rect 3191 5188 3700 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3694 5176 3700 5188
rect 3752 5216 3758 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3752 5188 3893 5216
rect 3752 5176 3758 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8754 5216 8760 5228
rect 8159 5188 8760 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8754 5176 8760 5188
rect 8812 5216 8818 5228
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8812 5188 9045 5216
rect 8812 5176 8818 5188
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 21266 5216 21272 5228
rect 21227 5188 21272 5216
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4706 5148 4712 5160
rect 4111 5120 4712 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8941 5151 8999 5157
rect 8941 5148 8953 5151
rect 7791 5120 8953 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8941 5117 8953 5120
rect 8987 5148 8999 5151
rect 9582 5148 9588 5160
rect 8987 5120 9588 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 14182 5148 14188 5160
rect 14143 5120 14188 5148
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21085 5151 21143 5157
rect 21085 5148 21097 5151
rect 20772 5120 21097 5148
rect 20772 5108 20778 5120
rect 21085 5117 21097 5120
rect 21131 5148 21143 5151
rect 21726 5148 21732 5160
rect 21131 5120 21732 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 14093 5083 14151 5089
rect 14093 5049 14105 5083
rect 14139 5080 14151 5083
rect 14430 5083 14488 5089
rect 14430 5080 14442 5083
rect 14139 5052 14442 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 14430 5049 14442 5052
rect 14476 5080 14488 5083
rect 14918 5080 14924 5092
rect 14476 5052 14924 5080
rect 14476 5049 14488 5052
rect 14430 5043 14488 5049
rect 14918 5040 14924 5052
rect 14976 5040 14982 5092
rect 20165 5083 20223 5089
rect 20165 5049 20177 5083
rect 20211 5080 20223 5083
rect 21358 5080 21364 5092
rect 20211 5052 21364 5080
rect 20211 5049 20223 5052
rect 20165 5043 20223 5049
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 3602 5012 3608 5024
rect 3007 4984 3608 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 4028 4984 4261 5012
rect 4028 4972 4034 4984
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 8570 5012 8576 5024
rect 8531 4984 8576 5012
rect 4249 4975 4307 4981
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 11422 5012 11428 5024
rect 11383 4984 11428 5012
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20312 4984 21005 5012
rect 20312 4972 20318 4984
rect 20993 4981 21005 4984
rect 21039 5012 21051 5015
rect 21726 5012 21732 5024
rect 21039 4984 21732 5012
rect 21039 4981 21051 4984
rect 20993 4975 21051 4981
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1452 4780 1593 4808
rect 1452 4768 1458 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2682 4808 2688 4820
rect 2455 4780 2688 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2866 4808 2872 4820
rect 2779 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4808 2930 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2924 4780 3433 4808
rect 2924 4768 2930 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4709 4811 4767 4817
rect 4709 4808 4721 4811
rect 4304 4780 4721 4808
rect 4304 4768 4310 4780
rect 4709 4777 4721 4780
rect 4755 4808 4767 4811
rect 5534 4808 5540 4820
rect 4755 4780 5540 4808
rect 4755 4777 4767 4780
rect 4709 4771 4767 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 7009 4811 7067 4817
rect 7009 4777 7021 4811
rect 7055 4808 7067 4811
rect 7374 4808 7380 4820
rect 7055 4780 7380 4808
rect 7055 4777 7067 4780
rect 7009 4771 7067 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 7607 4780 8401 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 8389 4777 8401 4780
rect 8435 4808 8447 4811
rect 8570 4808 8576 4820
rect 8435 4780 8576 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 10502 4808 10508 4820
rect 10463 4780 10508 4808
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 11480 4780 12817 4808
rect 11480 4768 11486 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 12805 4771 12863 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 20901 4811 20959 4817
rect 20901 4777 20913 4811
rect 20947 4808 20959 4811
rect 21358 4808 21364 4820
rect 20947 4780 21364 4808
rect 20947 4777 20959 4780
rect 20901 4771 20959 4777
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 11606 4700 11612 4752
rect 11664 4749 11670 4752
rect 11664 4743 11728 4749
rect 11664 4709 11682 4743
rect 11716 4709 11728 4743
rect 11664 4703 11728 4709
rect 11664 4700 11670 4703
rect 11882 4700 11888 4752
rect 11940 4700 11946 4752
rect 16758 4749 16764 4752
rect 16752 4740 16764 4749
rect 16719 4712 16764 4740
rect 16752 4703 16764 4712
rect 16758 4700 16764 4703
rect 16816 4700 16822 4752
rect 21174 4700 21180 4752
rect 21232 4740 21238 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 21232 4712 21281 4740
rect 21232 4700 21238 4712
rect 21269 4709 21281 4712
rect 21315 4740 21327 4743
rect 21542 4740 21548 4752
rect 21315 4712 21548 4740
rect 21315 4709 21327 4712
rect 21269 4703 21327 4709
rect 21542 4700 21548 4712
rect 21600 4700 21606 4752
rect 2317 4675 2375 4681
rect 2317 4641 2329 4675
rect 2363 4672 2375 4675
rect 2406 4672 2412 4684
rect 2363 4644 2412 4672
rect 2363 4641 2375 4644
rect 2317 4635 2375 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 2777 4675 2835 4681
rect 2777 4672 2789 4675
rect 2648 4644 2789 4672
rect 2648 4632 2654 4644
rect 2777 4641 2789 4644
rect 2823 4641 2835 4675
rect 2777 4635 2835 4641
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4614 4672 4620 4684
rect 4111 4644 4620 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11900 4672 11928 4700
rect 14182 4672 14188 4684
rect 11471 4644 14188 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 16482 4672 16488 4684
rect 16443 4644 16488 4672
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 26510 4672 26516 4684
rect 26471 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4632 26574 4684
rect 2424 4604 2452 4632
rect 3050 4604 3056 4616
rect 2424 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4604 7987 4607
rect 8478 4604 8484 4616
rect 7975 4576 8484 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 8628 4576 8673 4604
rect 20824 4576 21373 4604
rect 8628 4564 8634 4576
rect 20824 4548 20852 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 20806 4496 20812 4548
rect 20864 4496 20870 4548
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 21266 4536 21272 4548
rect 21048 4508 21272 4536
rect 21048 4496 21054 4508
rect 21266 4496 21272 4508
rect 21324 4536 21330 4548
rect 21468 4536 21496 4567
rect 21910 4536 21916 4548
rect 21324 4508 21916 4536
rect 21324 4496 21330 4508
rect 21910 4496 21916 4508
rect 21968 4496 21974 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4212 4440 4261 4468
rect 4212 4428 4218 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 6880 4440 8033 4468
rect 6880 4428 6886 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17862 4468 17868 4480
rect 16908 4440 17868 4468
rect 16908 4428 16914 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 26694 4468 26700 4480
rect 26655 4440 26700 4468
rect 26694 4428 26700 4440
rect 26752 4428 26758 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 2685 4267 2743 4273
rect 2685 4233 2697 4267
rect 2731 4264 2743 4267
rect 2866 4264 2872 4276
rect 2731 4236 2872 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3694 4264 3700 4276
rect 3655 4236 3700 4264
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 5316 4236 5641 4264
rect 5316 4224 5322 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8536 4236 8953 4264
rect 8536 4224 8542 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 8941 4227 8999 4233
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 21174 4264 21180 4276
rect 20947 4236 21180 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26568 4236 27353 4264
rect 26568 4224 26574 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 3142 4128 3148 4140
rect 2639 4100 3148 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3292 4100 3341 4128
rect 3292 4088 3298 4100
rect 3329 4097 3341 4100
rect 3375 4128 3387 4131
rect 3712 4128 3740 4224
rect 8570 4196 8576 4208
rect 8220 4168 8576 4196
rect 3375 4100 4384 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4020 1458 4072
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 4246 4060 4252 4072
rect 3752 4032 4252 4060
rect 3752 4020 3758 4032
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 4356 4060 4384 4100
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 5592 4100 6561 4128
rect 5592 4088 5598 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 4522 4069 4528 4072
rect 4505 4063 4528 4069
rect 4505 4060 4517 4063
rect 4356 4032 4517 4060
rect 4505 4029 4517 4032
rect 4580 4060 4586 4072
rect 4580 4032 4653 4060
rect 4505 4023 4528 4029
rect 4522 4020 4528 4023
rect 4580 4020 4586 4032
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 4614 3992 4620 4004
rect 4203 3964 4620 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 6564 3992 6592 4091
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8220 4128 8248 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 10502 4196 10508 4208
rect 9732 4168 10508 4196
rect 9732 4156 9738 4168
rect 10502 4156 10508 4168
rect 10560 4196 10566 4208
rect 14461 4199 14519 4205
rect 10560 4168 11008 4196
rect 10560 4156 10566 4168
rect 8159 4100 8248 4128
rect 8849 4131 8907 4137
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9214 4128 9220 4140
rect 8895 4100 9220 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9214 4088 9220 4100
rect 9272 4128 9278 4140
rect 9582 4128 9588 4140
rect 9272 4100 9588 4128
rect 9272 4088 9278 4100
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 10410 4088 10416 4100
rect 10468 4128 10474 4140
rect 10980 4128 11008 4168
rect 14461 4165 14473 4199
rect 14507 4196 14519 4199
rect 20990 4196 20996 4208
rect 14507 4168 15148 4196
rect 14507 4165 14519 4168
rect 14461 4159 14519 4165
rect 15120 4140 15148 4168
rect 20640 4168 20996 4196
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10468 4100 10916 4128
rect 10980 4100 11069 4128
rect 10468 4088 10474 4100
rect 7282 4060 7288 4072
rect 7243 4032 7288 4060
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8754 4060 8760 4072
rect 8527 4032 8760 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 8812 4032 9413 4060
rect 8812 4020 8818 4032
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 10888 4069 10916 4100
rect 11057 4097 11069 4100
rect 11103 4128 11115 4131
rect 11330 4128 11336 4140
rect 11103 4100 11336 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 15102 4128 15108 4140
rect 15063 4100 15108 4128
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16850 4128 16856 4140
rect 16347 4100 16856 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16850 4088 16856 4100
rect 16908 4128 16914 4140
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16908 4100 16957 4128
rect 16908 4088 16914 4100
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4128 20223 4131
rect 20640 4128 20668 4168
rect 20990 4156 20996 4168
rect 21048 4156 21054 4208
rect 22922 4196 22928 4208
rect 22020 4168 22928 4196
rect 20211 4100 20668 4128
rect 20916 4100 21128 4128
rect 20211 4097 20223 4100
rect 20165 4091 20223 4097
rect 10873 4063 10931 4069
rect 10376 4032 10640 4060
rect 10376 4020 10382 4032
rect 7377 3995 7435 4001
rect 7377 3992 7389 3995
rect 6564 3964 7389 3992
rect 7377 3961 7389 3964
rect 7423 3992 7435 3995
rect 7466 3992 7472 4004
rect 7423 3964 7472 3992
rect 7423 3961 7435 3964
rect 7377 3955 7435 3961
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 9180 3964 9321 3992
rect 9180 3952 9186 3964
rect 9309 3961 9321 3964
rect 9355 3992 9367 3995
rect 10612 3992 10640 4032
rect 10873 4029 10885 4063
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14700 4032 14933 4060
rect 14700 4020 14706 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15068 4032 15113 4060
rect 15068 4020 15074 4032
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16724 4032 16773 4060
rect 16724 4020 16730 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20916 4060 20944 4100
rect 20404 4032 20944 4060
rect 20993 4063 21051 4069
rect 20404 4020 20410 4032
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 21100 4060 21128 4100
rect 22020 4060 22048 4168
rect 22922 4156 22928 4168
rect 22980 4156 22986 4208
rect 26418 4060 26424 4072
rect 21039 4032 22048 4060
rect 26379 4032 26424 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 26418 4020 26424 4032
rect 26476 4060 26482 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26476 4032 26985 4060
rect 26476 4020 26482 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 21266 4001 21272 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 9355 3964 10548 3992
rect 10612 3964 10977 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 3053 3927 3111 3933
rect 3053 3924 3065 3927
rect 2271 3896 3065 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 3053 3893 3065 3896
rect 3099 3924 3111 3927
rect 5166 3924 5172 3936
rect 3099 3896 5172 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6917 3927 6975 3933
rect 6917 3893 6929 3927
rect 6963 3924 6975 3927
rect 7190 3924 7196 3936
rect 6963 3896 7196 3924
rect 6963 3893 6975 3896
rect 6917 3887 6975 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 10520 3933 10548 3964
rect 10965 3961 10977 3964
rect 11011 3961 11023 3995
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 10965 3955 11023 3961
rect 14568 3964 15853 3992
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3893 10563 3927
rect 11606 3924 11612 3936
rect 11567 3896 11612 3924
rect 10505 3887 10563 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 14568 3933 14596 3964
rect 15841 3961 15853 3964
rect 15887 3992 15899 3995
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 15887 3964 16865 3992
rect 15887 3961 15899 3964
rect 15841 3955 15899 3961
rect 16853 3961 16865 3964
rect 16899 3961 16911 3995
rect 16853 3955 16911 3961
rect 20533 3995 20591 4001
rect 20533 3961 20545 3995
rect 20579 3992 20591 3995
rect 21260 3992 21272 4001
rect 20579 3964 21272 3992
rect 20579 3961 20591 3964
rect 20533 3955 20591 3961
rect 21260 3955 21272 3964
rect 21266 3952 21272 3955
rect 21324 3952 21330 4004
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3893 14611 3927
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 14553 3887 14611 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 16632 3896 17417 3924
rect 16632 3884 16638 3896
rect 17405 3893 17417 3896
rect 17451 3924 17463 3927
rect 18138 3924 18144 3936
rect 17451 3896 18144 3924
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22373 3927 22431 3933
rect 22373 3924 22385 3927
rect 21968 3896 22385 3924
rect 21968 3884 21974 3896
rect 22373 3893 22385 3896
rect 22419 3893 22431 3927
rect 22373 3887 22431 3893
rect 26605 3927 26663 3933
rect 26605 3893 26617 3927
rect 26651 3924 26663 3927
rect 26786 3924 26792 3936
rect 26651 3896 26792 3924
rect 26651 3893 26663 3896
rect 26605 3887 26663 3893
rect 26786 3884 26792 3896
rect 26844 3884 26850 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1452 3692 1593 3720
rect 1452 3680 1458 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 1581 3683 1639 3689
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 2958 3720 2964 3732
rect 2915 3692 2964 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3108 3692 3433 3720
rect 3108 3680 3114 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4580 3692 4629 3720
rect 4580 3680 4586 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7282 3720 7288 3732
rect 7055 3692 7288 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 9122 3720 9128 3732
rect 9083 3692 9128 3720
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 10376 3692 10517 3720
rect 10376 3680 10382 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 11664 3692 12449 3720
rect 11664 3680 11670 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 15010 3720 15016 3732
rect 14691 3692 15016 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 16666 3680 16672 3732
rect 16724 3720 16730 3732
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 16724 3692 16865 3720
rect 16724 3680 16730 3692
rect 16853 3689 16865 3692
rect 16899 3689 16911 3723
rect 20346 3720 20352 3732
rect 20307 3692 20352 3720
rect 16853 3683 16911 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20717 3723 20775 3729
rect 20717 3689 20729 3723
rect 20763 3720 20775 3723
rect 20806 3720 20812 3732
rect 20763 3692 20812 3720
rect 20763 3689 20775 3692
rect 20717 3683 20775 3689
rect 20806 3680 20812 3692
rect 20864 3720 20870 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 20864 3692 20913 3720
rect 20864 3680 20870 3692
rect 20901 3689 20913 3692
rect 20947 3689 20959 3723
rect 21358 3720 21364 3732
rect 21319 3692 21364 3720
rect 20901 3683 20959 3689
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 7374 3661 7380 3664
rect 7368 3652 7380 3661
rect 7335 3624 7380 3652
rect 7368 3615 7380 3624
rect 7374 3612 7380 3615
rect 7432 3612 7438 3664
rect 11514 3652 11520 3664
rect 11072 3624 11520 3652
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 3602 3584 3608 3596
rect 2823 3556 3608 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 2884 3528 2912 3556
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3804 3556 4077 3584
rect 3804 3528 3832 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 4065 3547 4123 3553
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7006 3584 7012 3596
rect 6788 3556 7012 3584
rect 6788 3544 6794 3556
rect 7006 3544 7012 3556
rect 7064 3584 7070 3596
rect 11072 3593 11100 3624
rect 11514 3612 11520 3624
rect 11572 3652 11578 3664
rect 11882 3652 11888 3664
rect 11572 3624 11888 3652
rect 11572 3612 11578 3624
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 16577 3655 16635 3661
rect 16577 3621 16589 3655
rect 16623 3652 16635 3655
rect 16758 3652 16764 3664
rect 16623 3624 16764 3652
rect 16623 3621 16635 3624
rect 16577 3615 16635 3621
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 17954 3612 17960 3664
rect 18012 3652 18018 3664
rect 18386 3655 18444 3661
rect 18386 3652 18398 3655
rect 18012 3624 18398 3652
rect 18012 3612 18018 3624
rect 18386 3621 18398 3624
rect 18432 3621 18444 3655
rect 18386 3615 18444 3621
rect 21269 3655 21327 3661
rect 21269 3621 21281 3655
rect 21315 3652 21327 3655
rect 21634 3652 21640 3664
rect 21315 3624 21640 3652
rect 21315 3621 21327 3624
rect 21269 3615 21327 3621
rect 21634 3612 21640 3624
rect 21692 3612 21698 3664
rect 11330 3593 11336 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 7064 3556 7113 3584
rect 7064 3544 7070 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11324 3584 11336 3593
rect 11291 3556 11336 3584
rect 11057 3547 11115 3553
rect 11324 3547 11336 3556
rect 11330 3544 11336 3547
rect 11388 3544 11394 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 24854 3544 24860 3596
rect 24912 3584 24918 3596
rect 25314 3584 25320 3596
rect 24912 3556 25320 3584
rect 24912 3544 24918 3556
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2363 3488 2820 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2792 3448 2820 3488
rect 2866 3476 2872 3528
rect 2924 3476 2930 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2976 3488 3065 3516
rect 2976 3448 3004 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3234 3516 3240 3528
rect 3099 3488 3240 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3234 3476 3240 3488
rect 3292 3476 3298 3528
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 2792 3420 3004 3448
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 5353 3451 5411 3457
rect 5353 3448 5365 3451
rect 4028 3420 5365 3448
rect 4028 3408 4034 3420
rect 5353 3417 5365 3420
rect 5399 3417 5411 3451
rect 5353 3411 5411 3417
rect 8481 3451 8539 3457
rect 8481 3417 8493 3451
rect 8527 3448 8539 3451
rect 9582 3448 9588 3460
rect 8527 3420 9588 3448
rect 8527 3417 8539 3420
rect 8481 3411 8539 3417
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 19521 3451 19579 3457
rect 19521 3417 19533 3451
rect 19567 3448 19579 3451
rect 21266 3448 21272 3460
rect 19567 3420 21272 3448
rect 19567 3417 19579 3420
rect 19521 3411 19579 3417
rect 21266 3408 21272 3420
rect 21324 3448 21330 3460
rect 21468 3448 21496 3479
rect 25498 3448 25504 3460
rect 21324 3420 21496 3448
rect 25459 3420 25504 3448
rect 21324 3408 21330 3420
rect 25498 3408 25504 3420
rect 25556 3408 25562 3460
rect 2409 3383 2467 3389
rect 2409 3349 2421 3383
rect 2455 3380 2467 3383
rect 2590 3380 2596 3392
rect 2455 3352 2596 3380
rect 2455 3349 2467 3352
rect 2409 3343 2467 3349
rect 2590 3340 2596 3352
rect 2648 3380 2654 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 2648 3352 3801 3380
rect 2648 3340 2654 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 4246 3380 4252 3392
rect 4207 3352 4252 3380
rect 3789 3343 3847 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 26694 3380 26700 3392
rect 26655 3352 26700 3380
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2774 3176 2780 3188
rect 1995 3148 2780 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3384 3148 3801 3176
rect 3384 3136 3390 3148
rect 3789 3145 3801 3148
rect 3835 3145 3847 3179
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 3789 3139 3847 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5445 3179 5503 3185
rect 5445 3176 5457 3179
rect 5224 3148 5457 3176
rect 5224 3136 5230 3148
rect 5445 3145 5457 3148
rect 5491 3145 5503 3179
rect 5445 3139 5503 3145
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7653 3179 7711 3185
rect 7653 3176 7665 3179
rect 7432 3148 7665 3176
rect 7432 3136 7438 3148
rect 7653 3145 7665 3148
rect 7699 3145 7711 3179
rect 8754 3176 8760 3188
rect 8715 3148 8760 3176
rect 7653 3139 7711 3145
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11330 3176 11336 3188
rect 11195 3148 11336 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18012 3148 18245 3176
rect 18012 3136 18018 3148
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 18233 3139 18291 3145
rect 20349 3179 20407 3185
rect 20349 3145 20361 3179
rect 20395 3176 20407 3179
rect 20530 3176 20536 3188
rect 20395 3148 20536 3176
rect 20395 3145 20407 3148
rect 20349 3139 20407 3145
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7248 3080 8217 3108
rect 7248 3068 7254 3080
rect 8205 3077 8217 3080
rect 8251 3108 8263 3111
rect 8251 3080 9260 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 9232 3049 9260 3080
rect 18138 3068 18144 3120
rect 18196 3108 18202 3120
rect 18601 3111 18659 3117
rect 18601 3108 18613 3111
rect 18196 3080 18613 3108
rect 18196 3068 18202 3080
rect 18601 3077 18613 3080
rect 18647 3077 18659 3111
rect 18601 3071 18659 3077
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 3844 3012 4353 3040
rect 3844 3000 3850 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3040 9459 3043
rect 9582 3040 9588 3052
rect 9447 3012 9588 3040
rect 9447 3009 9459 3012
rect 9401 3003 9459 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2958 2972 2964 2984
rect 2455 2944 2964 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4856 2944 4905 2972
rect 4856 2932 4862 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 6641 2975 6699 2981
rect 6641 2941 6653 2975
rect 6687 2972 6699 2975
rect 6914 2972 6920 2984
rect 6687 2944 6920 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 9030 2972 9036 2984
rect 8711 2944 9036 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 9030 2932 9036 2944
rect 9088 2972 9094 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 9088 2944 9137 2972
rect 9088 2932 9094 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 10192 2944 10333 2972
rect 10192 2932 10198 2944
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 20456 2981 20484 3148
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 21358 3176 21364 3188
rect 21315 3148 21364 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 21634 3176 21640 3188
rect 21595 3148 21640 3176
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 24302 3136 24308 3188
rect 24360 3176 24366 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24360 3148 24409 3176
rect 24360 3136 24366 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 25314 3176 25320 3188
rect 25275 3148 25320 3176
rect 24397 3139 24455 3145
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 27341 3179 27399 3185
rect 27341 3176 27353 3179
rect 26568 3148 27353 3176
rect 26568 3136 26574 3148
rect 27341 3145 27353 3148
rect 27387 3145 27399 3179
rect 27341 3139 27399 3145
rect 27065 3111 27123 3117
rect 27065 3077 27077 3111
rect 27111 3108 27123 3111
rect 27246 3108 27252 3120
rect 27111 3080 27252 3108
rect 27111 3077 27123 3080
rect 27065 3071 27123 3077
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 13596 2944 13645 2972
rect 13596 2932 13602 2944
rect 13633 2941 13645 2944
rect 13679 2972 13691 2975
rect 14369 2975 14427 2981
rect 14369 2972 14381 2975
rect 13679 2944 14381 2972
rect 13679 2941 13691 2944
rect 13633 2935 13691 2941
rect 14369 2941 14381 2944
rect 14415 2941 14427 2975
rect 14369 2935 14427 2941
rect 20441 2975 20499 2981
rect 20441 2941 20453 2975
rect 20487 2941 20499 2975
rect 20441 2935 20499 2941
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2972 23719 2975
rect 24302 2972 24308 2984
rect 23707 2944 24308 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24302 2932 24308 2944
rect 24360 2932 24366 2984
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2972 26479 2975
rect 27080 2972 27108 3071
rect 27246 3068 27252 3080
rect 27304 3068 27310 3120
rect 27522 2972 27528 2984
rect 26467 2944 27108 2972
rect 27435 2944 27528 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27580 2944 28089 2972
rect 27580 2932 27586 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 2654 2907 2712 2913
rect 2654 2904 2666 2907
rect 2240 2876 2666 2904
rect 2038 2796 2044 2848
rect 2096 2836 2102 2848
rect 2240 2845 2268 2876
rect 2654 2873 2666 2876
rect 2700 2873 2712 2907
rect 2654 2867 2712 2873
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 7742 2904 7748 2916
rect 7239 2876 7748 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 10597 2907 10655 2913
rect 10597 2873 10609 2907
rect 10643 2904 10655 2907
rect 12066 2904 12072 2916
rect 10643 2876 12072 2904
rect 10643 2873 10655 2876
rect 10597 2867 10655 2873
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 13909 2907 13967 2913
rect 13909 2873 13921 2907
rect 13955 2904 13967 2907
rect 14918 2904 14924 2916
rect 13955 2876 14924 2904
rect 13955 2873 13967 2876
rect 13909 2867 13967 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 20717 2907 20775 2913
rect 20717 2904 20729 2907
rect 20680 2876 20729 2904
rect 20680 2864 20686 2876
rect 20717 2873 20729 2876
rect 20763 2873 20775 2907
rect 20717 2867 20775 2873
rect 23937 2907 23995 2913
rect 23937 2873 23949 2907
rect 23983 2904 23995 2907
rect 24854 2904 24860 2916
rect 23983 2876 24860 2904
rect 23983 2873 23995 2876
rect 23937 2867 23995 2873
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 2096 2808 2237 2836
rect 2096 2796 2102 2808
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 2225 2799 2283 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2836 27767 2839
rect 27798 2836 27804 2848
rect 27755 2808 27804 2836
rect 27755 2805 27767 2808
rect 27709 2799 27767 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 2682 2632 2688 2644
rect 2643 2604 2688 2632
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 2832 2604 3065 2632
rect 2832 2592 2838 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 3053 2595 3111 2601
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6822 2632 6828 2644
rect 6411 2604 6828 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 2792 2564 2820 2592
rect 2087 2536 2820 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 2056 2496 2084 2527
rect 2958 2524 2964 2576
rect 3016 2564 3022 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 3016 2536 3433 2564
rect 3016 2524 3022 2536
rect 3421 2533 3433 2536
rect 3467 2564 3479 2567
rect 3694 2564 3700 2576
rect 3467 2536 3700 2564
rect 3467 2533 3479 2536
rect 3421 2527 3479 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 1443 2468 2084 2496
rect 2409 2499 2467 2505
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2498 2496 2504 2508
rect 2455 2468 2504 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2496 4126 2508
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4120 2468 4813 2496
rect 4120 2456 4126 2468
rect 4801 2465 4813 2468
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 6380 2496 6408 2595
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 7064 2604 7113 2632
rect 7064 2592 7070 2604
rect 7101 2601 7113 2604
rect 7147 2601 7159 2635
rect 7101 2595 7159 2601
rect 8849 2635 8907 2641
rect 8849 2601 8861 2635
rect 8895 2632 8907 2635
rect 9582 2632 9588 2644
rect 8895 2604 9588 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 19242 2632 19248 2644
rect 19203 2604 19248 2632
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20625 2635 20683 2641
rect 20625 2601 20637 2635
rect 20671 2632 20683 2635
rect 20806 2632 20812 2644
rect 20671 2604 20812 2632
rect 20671 2601 20683 2604
rect 20625 2595 20683 2601
rect 7558 2496 7564 2508
rect 5583 2468 6408 2496
rect 7519 2468 7564 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 7558 2456 7564 2468
rect 7616 2496 7622 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 7616 2468 8309 2496
rect 7616 2456 7622 2468
rect 8297 2465 8309 2468
rect 8343 2465 8355 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8297 2459 8355 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 9824 2468 10517 2496
rect 9824 2456 9830 2468
rect 10505 2465 10517 2468
rect 10551 2465 10563 2499
rect 10505 2459 10563 2465
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10744 2468 11161 2496
rect 10744 2456 10750 2468
rect 11149 2465 11161 2468
rect 11195 2496 11207 2499
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11195 2468 11897 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 13872 2468 14105 2496
rect 13872 2456 13878 2468
rect 14093 2465 14105 2468
rect 14139 2496 14151 2499
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14139 2468 14841 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 16390 2496 16396 2508
rect 16351 2468 16396 2496
rect 14829 2459 14887 2465
rect 16390 2456 16396 2468
rect 16448 2496 16454 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16448 2468 17141 2496
rect 16448 2456 16454 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 19260 2496 19288 2592
rect 18555 2468 19288 2496
rect 19797 2499 19855 2505
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 19797 2465 19809 2499
rect 19843 2496 19855 2499
rect 20640 2496 20668 2595
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 20993 2635 21051 2641
rect 20993 2601 21005 2635
rect 21039 2632 21051 2635
rect 21266 2632 21272 2644
rect 21039 2604 21272 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 19843 2468 20668 2496
rect 19843 2465 19855 2468
rect 19797 2459 19855 2465
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 22152 2468 22293 2496
rect 22152 2456 22158 2468
rect 22281 2465 22293 2468
rect 22327 2496 22339 2499
rect 23017 2499 23075 2505
rect 23017 2496 23029 2499
rect 22327 2468 23029 2496
rect 22327 2465 22339 2468
rect 22281 2459 22339 2465
rect 23017 2465 23029 2468
rect 23063 2465 23075 2499
rect 24302 2496 24308 2508
rect 24263 2468 24308 2496
rect 23017 2459 23075 2465
rect 24302 2456 24308 2468
rect 24360 2496 24366 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24360 2468 25053 2496
rect 24360 2456 24366 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 25130 2456 25136 2508
rect 25188 2496 25194 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25188 2468 25697 2496
rect 25188 2456 25194 2468
rect 25685 2465 25697 2468
rect 25731 2496 25743 2499
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25731 2468 26249 2496
rect 25731 2465 25743 2468
rect 25685 2459 25743 2465
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4890 2428 4896 2440
rect 4387 2400 4896 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6362 2428 6368 2440
rect 5859 2400 6368 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 9214 2428 9220 2440
rect 7883 2400 9220 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10594 2428 10600 2440
rect 10091 2400 10600 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 13446 2428 13452 2440
rect 11471 2400 13452 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 16298 2428 16304 2440
rect 14415 2400 16304 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2428 16727 2431
rect 17770 2428 17776 2440
rect 16715 2400 17776 2428
rect 16715 2397 16727 2400
rect 16669 2391 16727 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18785 2431 18843 2437
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 19150 2428 19156 2440
rect 18831 2400 19156 2428
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 22002 2428 22008 2440
rect 20119 2400 22008 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 23474 2428 23480 2440
rect 22603 2400 23480 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2428 24639 2431
rect 26326 2428 26332 2440
rect 24627 2400 26332 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 27065 2295 27123 2301
rect 27065 2261 27077 2295
rect 27111 2292 27123 2295
rect 29178 2292 29184 2304
rect 27111 2264 29184 2292
rect 27111 2261 27123 2264
rect 27065 2255 27123 2261
rect 29178 2252 29184 2264
rect 29236 2252 29242 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3424 22108 3476 22160
rect 10416 22108 10468 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 22376 20952 22428 21004
rect 22284 20927 22336 20936
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 2872 20748 2924 20800
rect 18052 20748 18104 20800
rect 23572 20748 23624 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 21548 20544 21600 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 20444 20340 20496 20392
rect 14096 20272 14148 20324
rect 19708 20272 19760 20324
rect 22284 20340 22336 20392
rect 23480 20272 23532 20324
rect 14832 20204 14884 20256
rect 26240 20247 26292 20256
rect 26240 20213 26249 20247
rect 26249 20213 26283 20247
rect 26283 20213 26292 20247
rect 26240 20204 26292 20213
rect 27528 20204 27580 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 19708 20043 19760 20052
rect 19708 20009 19717 20043
rect 19717 20009 19751 20043
rect 19751 20009 19760 20043
rect 19708 20000 19760 20009
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 22468 20000 22520 20052
rect 18328 19932 18380 19984
rect 23572 19864 23624 19916
rect 17960 19796 18012 19848
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 24952 19660 25004 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 13636 19320 13688 19372
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 18328 19320 18380 19372
rect 15844 19252 15896 19304
rect 17960 19252 18012 19304
rect 23480 19252 23532 19304
rect 8484 19227 8536 19236
rect 8484 19193 8493 19227
rect 8493 19193 8527 19227
rect 8527 19193 8536 19227
rect 8484 19184 8536 19193
rect 10324 19116 10376 19168
rect 14832 19116 14884 19168
rect 18604 19227 18656 19236
rect 18604 19193 18613 19227
rect 18613 19193 18647 19227
rect 18647 19193 18656 19227
rect 18604 19184 18656 19193
rect 24952 19184 25004 19236
rect 16488 19159 16540 19168
rect 16488 19125 16497 19159
rect 16497 19125 16531 19159
rect 16531 19125 16540 19159
rect 16488 19116 16540 19125
rect 18328 19116 18380 19168
rect 18696 19159 18748 19168
rect 18696 19125 18705 19159
rect 18705 19125 18739 19159
rect 18739 19125 18748 19159
rect 18696 19116 18748 19125
rect 18788 19116 18840 19168
rect 23572 19116 23624 19168
rect 24400 19116 24452 19168
rect 25688 19116 25740 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 14096 18955 14148 18964
rect 14096 18921 14105 18955
rect 14105 18921 14139 18955
rect 14139 18921 14148 18955
rect 14096 18912 14148 18921
rect 14464 18912 14516 18964
rect 18788 18955 18840 18964
rect 18788 18921 18797 18955
rect 18797 18921 18831 18955
rect 18831 18921 18840 18955
rect 18788 18912 18840 18921
rect 21824 18912 21876 18964
rect 24216 18912 24268 18964
rect 24952 18912 25004 18964
rect 4160 18776 4212 18828
rect 8576 18776 8628 18828
rect 9220 18776 9272 18828
rect 10692 18844 10744 18896
rect 18328 18887 18380 18896
rect 18328 18853 18337 18887
rect 18337 18853 18371 18887
rect 18371 18853 18380 18887
rect 18328 18844 18380 18853
rect 10324 18776 10376 18828
rect 12808 18776 12860 18828
rect 18696 18776 18748 18828
rect 23204 18819 23256 18828
rect 23204 18785 23213 18819
rect 23213 18785 23247 18819
rect 23247 18785 23256 18819
rect 23204 18776 23256 18785
rect 23296 18819 23348 18828
rect 23296 18785 23305 18819
rect 23305 18785 23339 18819
rect 23339 18785 23348 18819
rect 23296 18776 23348 18785
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 4068 18751 4120 18760
rect 1492 18572 1544 18624
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 18880 18708 18932 18760
rect 19708 18708 19760 18760
rect 21548 18751 21600 18760
rect 21272 18640 21324 18692
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 22744 18708 22796 18760
rect 24308 18708 24360 18760
rect 25688 18708 25740 18760
rect 5448 18615 5500 18624
rect 5448 18581 5457 18615
rect 5457 18581 5491 18615
rect 5491 18581 5500 18615
rect 5448 18572 5500 18581
rect 7380 18572 7432 18624
rect 10876 18572 10928 18624
rect 12716 18572 12768 18624
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 21364 18572 21416 18624
rect 22836 18615 22888 18624
rect 22836 18581 22845 18615
rect 22845 18581 22879 18615
rect 22879 18581 22888 18615
rect 22836 18572 22888 18581
rect 24400 18572 24452 18624
rect 25780 18572 25832 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 4068 18368 4120 18420
rect 5632 18368 5684 18420
rect 8484 18411 8536 18420
rect 3792 18300 3844 18352
rect 4160 18343 4212 18352
rect 4160 18309 4169 18343
rect 4169 18309 4203 18343
rect 4203 18309 4212 18343
rect 4160 18300 4212 18309
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 9588 18368 9640 18420
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 12808 18411 12860 18420
rect 12808 18377 12817 18411
rect 12817 18377 12851 18411
rect 12851 18377 12860 18411
rect 12808 18368 12860 18377
rect 18696 18368 18748 18420
rect 18880 18411 18932 18420
rect 18880 18377 18889 18411
rect 18889 18377 18923 18411
rect 18923 18377 18932 18411
rect 18880 18368 18932 18377
rect 19708 18368 19760 18420
rect 21548 18411 21600 18420
rect 12624 18300 12676 18352
rect 14004 18300 14056 18352
rect 18328 18343 18380 18352
rect 18328 18309 18337 18343
rect 18337 18309 18371 18343
rect 18371 18309 18380 18343
rect 18328 18300 18380 18309
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 21824 18411 21876 18420
rect 21824 18377 21833 18411
rect 21833 18377 21867 18411
rect 21867 18377 21876 18411
rect 21824 18368 21876 18377
rect 23204 18368 23256 18420
rect 25228 18368 25280 18420
rect 25504 18368 25556 18420
rect 21272 18300 21324 18352
rect 22744 18343 22796 18352
rect 22744 18309 22753 18343
rect 22753 18309 22787 18343
rect 22787 18309 22796 18343
rect 22744 18300 22796 18309
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 25688 18275 25740 18284
rect 25688 18241 25697 18275
rect 25697 18241 25731 18275
rect 25731 18241 25740 18275
rect 25688 18232 25740 18241
rect 1492 18164 1544 18216
rect 2504 18096 2556 18148
rect 7380 18139 7432 18148
rect 7380 18105 7414 18139
rect 7414 18105 7432 18139
rect 7380 18096 7432 18105
rect 19340 18164 19392 18216
rect 20444 18164 20496 18216
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 24768 18164 24820 18216
rect 14740 18139 14792 18148
rect 14740 18105 14749 18139
rect 14749 18105 14783 18139
rect 14783 18105 14792 18139
rect 14740 18096 14792 18105
rect 19156 18096 19208 18148
rect 9772 18028 9824 18080
rect 10324 18028 10376 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 13912 18028 13964 18080
rect 18604 18028 18656 18080
rect 22192 18096 22244 18148
rect 20720 18028 20772 18080
rect 25688 18096 25740 18148
rect 25780 18028 25832 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 1768 17824 1820 17876
rect 2964 17824 3016 17876
rect 13728 17824 13780 17876
rect 18880 17824 18932 17876
rect 19248 17867 19300 17876
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 20628 17824 20680 17876
rect 21272 17824 21324 17876
rect 22376 17824 22428 17876
rect 22836 17824 22888 17876
rect 23296 17824 23348 17876
rect 5448 17756 5500 17808
rect 13452 17756 13504 17808
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 5632 17731 5684 17740
rect 5632 17697 5641 17731
rect 5641 17697 5675 17731
rect 5675 17697 5684 17731
rect 5632 17688 5684 17697
rect 10416 17688 10468 17740
rect 11060 17688 11112 17740
rect 14004 17731 14056 17740
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 9956 17620 10008 17672
rect 14096 17663 14148 17672
rect 9680 17552 9732 17604
rect 10232 17552 10284 17604
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 16488 17756 16540 17808
rect 19156 17756 19208 17808
rect 22192 17799 22244 17808
rect 22192 17765 22201 17799
rect 22201 17765 22235 17799
rect 22235 17765 22244 17799
rect 22192 17756 22244 17765
rect 15844 17688 15896 17740
rect 19340 17688 19392 17740
rect 23204 17688 23256 17740
rect 23664 17731 23716 17740
rect 23664 17697 23673 17731
rect 23673 17697 23707 17731
rect 23707 17697 23716 17731
rect 23664 17688 23716 17697
rect 24768 17688 24820 17740
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 23848 17663 23900 17672
rect 18328 17552 18380 17604
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 24216 17620 24268 17672
rect 19984 17552 20036 17604
rect 1768 17527 1820 17536
rect 1768 17493 1777 17527
rect 1777 17493 1811 17527
rect 1811 17493 1820 17527
rect 1768 17484 1820 17493
rect 2320 17484 2372 17536
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 4712 17527 4764 17536
rect 4712 17493 4721 17527
rect 4721 17493 4755 17527
rect 4755 17493 4764 17527
rect 4712 17484 4764 17493
rect 7380 17484 7432 17536
rect 9772 17484 9824 17536
rect 10140 17527 10192 17536
rect 10140 17493 10149 17527
rect 10149 17493 10183 17527
rect 10183 17493 10192 17527
rect 10140 17484 10192 17493
rect 13636 17527 13688 17536
rect 13636 17493 13645 17527
rect 13645 17493 13679 17527
rect 13679 17493 13688 17527
rect 13636 17484 13688 17493
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 24124 17484 24176 17536
rect 25688 17484 25740 17536
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 1676 17280 1728 17332
rect 2228 17280 2280 17332
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 5448 17280 5500 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 14004 17280 14056 17332
rect 16488 17280 16540 17332
rect 18328 17280 18380 17332
rect 19340 17323 19392 17332
rect 19340 17289 19349 17323
rect 19349 17289 19383 17323
rect 19383 17289 19392 17323
rect 19340 17280 19392 17289
rect 20628 17280 20680 17332
rect 24768 17323 24820 17332
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 1768 17144 1820 17196
rect 4160 17144 4212 17196
rect 4436 17144 4488 17196
rect 9772 17212 9824 17264
rect 5632 17144 5684 17196
rect 10140 17144 10192 17196
rect 14096 17212 14148 17264
rect 14740 17144 14792 17196
rect 15844 17144 15896 17196
rect 16672 17144 16724 17196
rect 18144 17144 18196 17196
rect 19984 17187 20036 17196
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 22100 17144 22152 17196
rect 24124 17187 24176 17196
rect 2320 17119 2372 17128
rect 2320 17085 2329 17119
rect 2329 17085 2363 17119
rect 2363 17085 2372 17119
rect 2320 17076 2372 17085
rect 9956 17076 10008 17128
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 12992 17076 13044 17128
rect 22376 17119 22428 17128
rect 22376 17085 22385 17119
rect 22385 17085 22419 17119
rect 22419 17085 22428 17119
rect 22376 17076 22428 17085
rect 24124 17153 24133 17187
rect 24133 17153 24167 17187
rect 24167 17153 24176 17187
rect 24124 17144 24176 17153
rect 24308 17187 24360 17196
rect 24308 17153 24317 17187
rect 24317 17153 24351 17187
rect 24351 17153 24360 17187
rect 24308 17144 24360 17153
rect 4712 17051 4764 17060
rect 4712 17017 4721 17051
rect 4721 17017 4755 17051
rect 4755 17017 4764 17051
rect 4712 17008 4764 17017
rect 10416 17008 10468 17060
rect 3700 16940 3752 16992
rect 4344 16983 4396 16992
rect 4344 16949 4353 16983
rect 4353 16949 4387 16983
rect 4387 16949 4396 16983
rect 4344 16940 4396 16949
rect 10784 16940 10836 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14648 16983 14700 16992
rect 14188 16940 14240 16949
rect 14648 16949 14657 16983
rect 14657 16949 14691 16983
rect 14691 16949 14700 16983
rect 14648 16940 14700 16949
rect 19708 17008 19760 17060
rect 23204 17051 23256 17060
rect 23204 17017 23213 17051
rect 23213 17017 23247 17051
rect 23247 17017 23256 17051
rect 23204 17008 23256 17017
rect 24032 17051 24084 17060
rect 24032 17017 24041 17051
rect 24041 17017 24075 17051
rect 24075 17017 24084 17051
rect 24032 17008 24084 17017
rect 25688 17008 25740 17060
rect 27160 17076 27212 17128
rect 14832 16940 14884 16992
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 19892 16983 19944 16992
rect 19892 16949 19901 16983
rect 19901 16949 19935 16983
rect 19935 16949 19944 16983
rect 19892 16940 19944 16949
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 27344 16983 27396 16992
rect 27344 16949 27353 16983
rect 27353 16949 27387 16983
rect 27387 16949 27396 16983
rect 27344 16940 27396 16949
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 1768 16736 1820 16788
rect 2688 16736 2740 16788
rect 4436 16736 4488 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 10692 16736 10744 16788
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 13636 16736 13688 16788
rect 19984 16736 20036 16788
rect 22100 16779 22152 16788
rect 22100 16745 22109 16779
rect 22109 16745 22143 16779
rect 22143 16745 22152 16779
rect 22100 16736 22152 16745
rect 24032 16736 24084 16788
rect 24308 16779 24360 16788
rect 24308 16745 24317 16779
rect 24317 16745 24351 16779
rect 24351 16745 24360 16779
rect 24308 16736 24360 16745
rect 2412 16600 2464 16652
rect 4896 16600 4948 16652
rect 2504 16532 2556 16584
rect 4528 16575 4580 16584
rect 4528 16541 4537 16575
rect 4537 16541 4571 16575
rect 4571 16541 4580 16575
rect 4528 16532 4580 16541
rect 3700 16464 3752 16516
rect 4160 16464 4212 16516
rect 6644 16532 6696 16584
rect 9680 16600 9732 16652
rect 10968 16668 11020 16720
rect 23848 16668 23900 16720
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 7380 16575 7432 16584
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 11060 16600 11112 16652
rect 13728 16600 13780 16652
rect 10876 16575 10928 16584
rect 7380 16532 7432 16541
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 18420 16643 18472 16652
rect 18420 16609 18454 16643
rect 18454 16609 18472 16643
rect 18420 16600 18472 16609
rect 19800 16600 19852 16652
rect 10784 16464 10836 16516
rect 14372 16532 14424 16584
rect 23480 16600 23532 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 21456 16532 21508 16584
rect 23848 16575 23900 16584
rect 13544 16464 13596 16516
rect 22744 16464 22796 16516
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 26424 16464 26476 16516
rect 3608 16396 3660 16448
rect 7748 16396 7800 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 20444 16396 20496 16448
rect 25688 16396 25740 16448
rect 26700 16439 26752 16448
rect 26700 16405 26709 16439
rect 26709 16405 26743 16439
rect 26743 16405 26752 16439
rect 26700 16396 26752 16405
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 2412 16192 2464 16244
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 6920 16192 6972 16244
rect 7288 16192 7340 16244
rect 9680 16192 9732 16244
rect 10416 16235 10468 16244
rect 10416 16201 10425 16235
rect 10425 16201 10459 16235
rect 10459 16201 10468 16235
rect 10416 16192 10468 16201
rect 11060 16192 11112 16244
rect 13544 16192 13596 16244
rect 18144 16192 18196 16244
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 21456 16235 21508 16244
rect 21456 16201 21465 16235
rect 21465 16201 21499 16235
rect 21499 16201 21508 16235
rect 21456 16192 21508 16201
rect 22744 16235 22796 16244
rect 22744 16201 22753 16235
rect 22753 16201 22787 16235
rect 22787 16201 22796 16235
rect 22744 16192 22796 16201
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 24124 16192 24176 16244
rect 24952 16192 25004 16244
rect 25412 16192 25464 16244
rect 26516 16235 26568 16244
rect 26516 16201 26525 16235
rect 26525 16201 26559 16235
rect 26559 16201 26568 16235
rect 26516 16192 26568 16201
rect 4528 16167 4580 16176
rect 4528 16133 4537 16167
rect 4537 16133 4571 16167
rect 4571 16133 4580 16167
rect 4528 16124 4580 16133
rect 14372 16124 14424 16176
rect 3700 16099 3752 16108
rect 3700 16065 3709 16099
rect 3709 16065 3743 16099
rect 3743 16065 3752 16099
rect 3700 16056 3752 16065
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 8484 16056 8536 16108
rect 9772 16056 9824 16108
rect 10232 16056 10284 16108
rect 13452 16056 13504 16108
rect 1676 15988 1728 16040
rect 2780 15988 2832 16040
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 8944 15988 8996 16040
rect 13820 15988 13872 16040
rect 23848 16124 23900 16176
rect 8760 15920 8812 15972
rect 10968 15920 11020 15972
rect 13452 15920 13504 15972
rect 18420 16056 18472 16108
rect 19984 16056 20036 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 18972 16031 19024 16040
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 1400 15852 1452 15904
rect 1768 15852 1820 15904
rect 2596 15852 2648 15904
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 4896 15895 4948 15904
rect 4896 15861 4905 15895
rect 4905 15861 4939 15895
rect 4939 15861 4948 15895
rect 4896 15852 4948 15861
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 7564 15852 7616 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 14740 15895 14792 15904
rect 14740 15861 14749 15895
rect 14749 15861 14783 15895
rect 14783 15861 14792 15895
rect 14740 15852 14792 15861
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15660 15895 15712 15904
rect 15200 15852 15252 15861
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 19432 15895 19484 15904
rect 15752 15852 15804 15861
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 19616 15852 19668 15904
rect 20812 15852 20864 15904
rect 23940 15920 23992 15972
rect 21732 15852 21784 15904
rect 24124 15895 24176 15904
rect 24124 15861 24133 15895
rect 24133 15861 24167 15895
rect 24167 15861 24176 15895
rect 24124 15852 24176 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 4896 15648 4948 15700
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 7288 15648 7340 15700
rect 8760 15648 8812 15700
rect 8944 15648 8996 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 10876 15648 10928 15700
rect 13544 15648 13596 15700
rect 15200 15648 15252 15700
rect 15752 15648 15804 15700
rect 19524 15648 19576 15700
rect 24124 15648 24176 15700
rect 4160 15580 4212 15632
rect 4436 15623 4488 15632
rect 4436 15589 4445 15623
rect 4445 15589 4479 15623
rect 4479 15589 4488 15623
rect 4436 15580 4488 15589
rect 7380 15580 7432 15632
rect 7932 15580 7984 15632
rect 16764 15580 16816 15632
rect 17500 15580 17552 15632
rect 23848 15580 23900 15632
rect 1492 15512 1544 15564
rect 1676 15555 1728 15564
rect 1676 15521 1710 15555
rect 1710 15521 1728 15555
rect 1676 15512 1728 15521
rect 9772 15512 9824 15564
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 20720 15555 20772 15564
rect 20720 15521 20729 15555
rect 20729 15521 20763 15555
rect 20763 15521 20772 15555
rect 20720 15512 20772 15521
rect 23204 15512 23256 15564
rect 26792 15512 26844 15564
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 3700 15376 3752 15428
rect 4804 15444 4856 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 13268 15444 13320 15496
rect 14464 15444 14516 15496
rect 23296 15376 23348 15428
rect 5816 15351 5868 15360
rect 5816 15317 5825 15351
rect 5825 15317 5859 15351
rect 5859 15317 5868 15351
rect 5816 15308 5868 15317
rect 7564 15308 7616 15360
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 13728 15308 13780 15360
rect 18236 15308 18288 15360
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 20168 15308 20220 15360
rect 21732 15308 21784 15360
rect 22652 15308 22704 15360
rect 23572 15444 23624 15496
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 27344 15444 27396 15496
rect 25688 15308 25740 15360
rect 26332 15308 26384 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 1676 15104 1728 15156
rect 2688 15147 2740 15156
rect 2688 15113 2697 15147
rect 2697 15113 2731 15147
rect 2731 15113 2740 15147
rect 2688 15104 2740 15113
rect 4436 15104 4488 15156
rect 4528 15147 4580 15156
rect 4528 15113 4537 15147
rect 4537 15113 4571 15147
rect 4571 15113 4580 15147
rect 4804 15147 4856 15156
rect 4528 15104 4580 15113
rect 4804 15113 4813 15147
rect 4813 15113 4847 15147
rect 4847 15113 4856 15147
rect 4804 15104 4856 15113
rect 5724 15104 5776 15156
rect 6368 15104 6420 15156
rect 10232 15104 10284 15156
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 13452 15104 13504 15156
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 16764 15147 16816 15156
rect 16764 15113 16773 15147
rect 16773 15113 16807 15147
rect 16807 15113 16816 15147
rect 16764 15104 16816 15113
rect 18972 15104 19024 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 6828 15011 6880 15020
rect 6828 14977 6837 15011
rect 6837 14977 6871 15011
rect 6871 14977 6880 15011
rect 6828 14968 6880 14977
rect 13544 14968 13596 15020
rect 14740 15036 14792 15088
rect 16672 15036 16724 15088
rect 17960 15036 18012 15088
rect 19708 15036 19760 15088
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 19984 14968 20036 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 4068 14900 4120 14952
rect 14556 14900 14608 14952
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 15476 14900 15528 14909
rect 19064 14900 19116 14952
rect 19524 14900 19576 14952
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 23296 14900 23348 14952
rect 25228 14968 25280 15020
rect 25780 14900 25832 14952
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 2780 14764 2832 14816
rect 6460 14832 6512 14884
rect 7104 14875 7156 14884
rect 7104 14841 7138 14875
rect 7138 14841 7156 14875
rect 7104 14832 7156 14841
rect 13176 14832 13228 14884
rect 13728 14832 13780 14884
rect 14924 14875 14976 14884
rect 14924 14841 14933 14875
rect 14933 14841 14967 14875
rect 14967 14841 14976 14875
rect 14924 14832 14976 14841
rect 15384 14832 15436 14884
rect 19892 14832 19944 14884
rect 20260 14832 20312 14884
rect 26148 14832 26200 14884
rect 26332 14875 26384 14884
rect 26332 14841 26366 14875
rect 26366 14841 26384 14875
rect 26332 14832 26384 14841
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10140 14807 10192 14816
rect 10140 14773 10149 14807
rect 10149 14773 10183 14807
rect 10183 14773 10192 14807
rect 10140 14764 10192 14773
rect 13268 14764 13320 14816
rect 23204 14764 23256 14816
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 27436 14807 27488 14816
rect 27436 14773 27445 14807
rect 27445 14773 27479 14807
rect 27479 14773 27488 14807
rect 27436 14764 27488 14773
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 1492 14560 1544 14612
rect 1676 14560 1728 14612
rect 3240 14560 3292 14612
rect 5816 14560 5868 14612
rect 9220 14603 9272 14612
rect 3700 14492 3752 14544
rect 5632 14492 5684 14544
rect 9220 14569 9229 14603
rect 9229 14569 9263 14603
rect 9263 14569 9272 14603
rect 9220 14560 9272 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 13544 14560 13596 14612
rect 26332 14560 26384 14612
rect 27344 14560 27396 14612
rect 1492 14424 1544 14476
rect 3240 14424 3292 14476
rect 7104 14424 7156 14476
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 7196 14356 7248 14408
rect 10232 14492 10284 14544
rect 8116 14424 8168 14476
rect 10876 14492 10928 14544
rect 14096 14492 14148 14544
rect 11704 14424 11756 14476
rect 9036 14356 9088 14408
rect 14464 14424 14516 14476
rect 15660 14424 15712 14476
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 17960 14467 18012 14476
rect 17960 14433 17969 14467
rect 17969 14433 18003 14467
rect 18003 14433 18012 14467
rect 17960 14424 18012 14433
rect 18236 14467 18288 14476
rect 18236 14433 18270 14467
rect 18270 14433 18288 14467
rect 18236 14424 18288 14433
rect 22652 14424 22704 14476
rect 6276 14288 6328 14340
rect 8208 14288 8260 14340
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 7932 14220 7984 14272
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 15844 14356 15896 14408
rect 22560 14399 22612 14408
rect 15568 14288 15620 14340
rect 22560 14365 22569 14399
rect 22569 14365 22603 14399
rect 22603 14365 22612 14399
rect 22560 14356 22612 14365
rect 14188 14220 14240 14272
rect 16396 14220 16448 14272
rect 16488 14220 16540 14272
rect 19340 14263 19392 14272
rect 19340 14229 19349 14263
rect 19349 14229 19383 14263
rect 19383 14229 19392 14263
rect 19340 14220 19392 14229
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 24032 14220 24084 14272
rect 25228 14220 25280 14272
rect 26792 14263 26844 14272
rect 26792 14229 26801 14263
rect 26801 14229 26835 14263
rect 26835 14229 26844 14263
rect 26792 14220 26844 14229
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 1492 14016 1544 14068
rect 1676 14016 1728 14068
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 5816 14016 5868 14068
rect 7104 14016 7156 14068
rect 10508 14059 10560 14068
rect 10508 14025 10517 14059
rect 10517 14025 10551 14059
rect 10551 14025 10560 14059
rect 10508 14016 10560 14025
rect 11704 14059 11756 14068
rect 11704 14025 11713 14059
rect 11713 14025 11747 14059
rect 11747 14025 11756 14059
rect 11704 14016 11756 14025
rect 12440 14016 12492 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 17960 14016 18012 14068
rect 19984 14016 20036 14068
rect 22652 14059 22704 14068
rect 22652 14025 22661 14059
rect 22661 14025 22695 14059
rect 22695 14025 22704 14059
rect 22652 14016 22704 14025
rect 25228 14016 25280 14068
rect 6276 13948 6328 14000
rect 6828 13948 6880 14000
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 8208 13880 8260 13932
rect 9220 13880 9272 13932
rect 11888 13948 11940 14000
rect 15200 13948 15252 14000
rect 23480 13948 23532 14000
rect 24032 13948 24084 14000
rect 7196 13855 7248 13864
rect 3240 13744 3292 13796
rect 7196 13821 7205 13855
rect 7205 13821 7239 13855
rect 7239 13821 7248 13855
rect 7196 13812 7248 13821
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 10876 13880 10928 13932
rect 14188 13880 14240 13932
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16212 13880 16264 13932
rect 9036 13812 9088 13821
rect 10232 13812 10284 13864
rect 10508 13812 10560 13864
rect 10600 13812 10652 13864
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 8024 13744 8076 13796
rect 9772 13744 9824 13796
rect 10416 13744 10468 13796
rect 11704 13744 11756 13796
rect 16764 13744 16816 13796
rect 7472 13676 7524 13728
rect 10232 13719 10284 13728
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 17868 13812 17920 13864
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 24492 13880 24544 13932
rect 25228 13923 25280 13932
rect 20444 13855 20496 13864
rect 20444 13821 20478 13855
rect 20478 13821 20496 13855
rect 20444 13812 20496 13821
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 26056 13880 26108 13889
rect 26332 13880 26384 13932
rect 27436 13880 27488 13932
rect 26240 13812 26292 13864
rect 17316 13676 17368 13728
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 22192 13676 22244 13728
rect 22560 13676 22612 13728
rect 24676 13719 24728 13728
rect 24676 13685 24685 13719
rect 24685 13685 24719 13719
rect 24719 13685 24728 13719
rect 24676 13676 24728 13685
rect 26332 13744 26384 13796
rect 27160 13744 27212 13796
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 6828 13472 6880 13524
rect 7472 13472 7524 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 10416 13472 10468 13524
rect 12440 13472 12492 13524
rect 5540 13404 5592 13456
rect 6552 13404 6604 13456
rect 8208 13404 8260 13456
rect 8760 13404 8812 13456
rect 8116 13336 8168 13388
rect 8852 13336 8904 13388
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 16304 13472 16356 13524
rect 16764 13515 16816 13524
rect 16764 13481 16773 13515
rect 16773 13481 16807 13515
rect 16807 13481 16816 13515
rect 16764 13472 16816 13481
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 17868 13472 17920 13524
rect 20168 13515 20220 13524
rect 20168 13481 20177 13515
rect 20177 13481 20211 13515
rect 20211 13481 20220 13515
rect 20168 13472 20220 13481
rect 24492 13472 24544 13524
rect 25136 13472 25188 13524
rect 26240 13515 26292 13524
rect 26240 13481 26249 13515
rect 26249 13481 26283 13515
rect 26283 13481 26292 13515
rect 26240 13472 26292 13481
rect 16212 13404 16264 13456
rect 17132 13447 17184 13456
rect 17132 13413 17141 13447
rect 17141 13413 17175 13447
rect 17175 13413 17184 13447
rect 17132 13404 17184 13413
rect 22560 13404 22612 13456
rect 23388 13404 23440 13456
rect 13360 13336 13412 13388
rect 18696 13379 18748 13388
rect 18696 13345 18705 13379
rect 18705 13345 18739 13379
rect 18739 13345 18748 13379
rect 18696 13336 18748 13345
rect 1860 13268 1912 13320
rect 3240 13268 3292 13320
rect 5724 13268 5776 13320
rect 8208 13200 8260 13252
rect 9036 13268 9088 13320
rect 10232 13268 10284 13320
rect 16580 13268 16632 13320
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 18328 13268 18380 13320
rect 18236 13200 18288 13252
rect 22192 13268 22244 13320
rect 26884 13379 26936 13388
rect 26884 13345 26893 13379
rect 26893 13345 26927 13379
rect 26927 13345 26936 13379
rect 26884 13336 26936 13345
rect 25228 13268 25280 13320
rect 26700 13268 26752 13320
rect 27436 13268 27488 13320
rect 18972 13200 19024 13252
rect 24860 13200 24912 13252
rect 25688 13243 25740 13252
rect 25688 13209 25697 13243
rect 25697 13209 25731 13243
rect 25731 13209 25740 13243
rect 25688 13200 25740 13209
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 10876 13132 10928 13184
rect 13912 13132 13964 13184
rect 14740 13175 14792 13184
rect 14740 13141 14749 13175
rect 14749 13141 14783 13175
rect 14783 13141 14792 13175
rect 14740 13132 14792 13141
rect 23480 13132 23532 13184
rect 24308 13132 24360 13184
rect 26332 13132 26384 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 5724 12928 5776 12980
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 8116 12928 8168 12980
rect 8760 12928 8812 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 15108 12928 15160 12980
rect 16488 12928 16540 12980
rect 17224 12928 17276 12980
rect 18972 12928 19024 12980
rect 22192 12971 22244 12980
rect 22192 12937 22201 12971
rect 22201 12937 22235 12971
rect 22235 12937 22244 12971
rect 22192 12928 22244 12937
rect 22560 12971 22612 12980
rect 22560 12937 22569 12971
rect 22569 12937 22603 12971
rect 22603 12937 22612 12971
rect 22560 12928 22612 12937
rect 26884 12928 26936 12980
rect 9036 12860 9088 12912
rect 14740 12860 14792 12912
rect 16212 12860 16264 12912
rect 16304 12860 16356 12912
rect 17132 12860 17184 12912
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 8300 12792 8352 12844
rect 9864 12792 9916 12844
rect 10876 12792 10928 12844
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 4712 12724 4764 12776
rect 5540 12724 5592 12776
rect 8484 12724 8536 12776
rect 12072 12724 12124 12776
rect 12900 12724 12952 12776
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 5356 12656 5408 12708
rect 10140 12699 10192 12708
rect 10140 12665 10149 12699
rect 10149 12665 10183 12699
rect 10183 12665 10192 12699
rect 10140 12656 10192 12665
rect 1768 12588 1820 12640
rect 4896 12588 4948 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 12900 12588 12952 12640
rect 13452 12724 13504 12776
rect 13912 12588 13964 12640
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 23848 12792 23900 12844
rect 24676 12860 24728 12912
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 25504 12835 25556 12844
rect 24308 12792 24360 12801
rect 25504 12801 25513 12835
rect 25513 12801 25547 12835
rect 25547 12801 25556 12835
rect 25504 12792 25556 12801
rect 14740 12767 14792 12776
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 15108 12724 15160 12776
rect 16212 12724 16264 12776
rect 16948 12724 17000 12776
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 24860 12724 24912 12776
rect 25688 12724 25740 12776
rect 26424 12724 26476 12776
rect 26700 12767 26752 12776
rect 26700 12733 26709 12767
rect 26709 12733 26743 12767
rect 26743 12733 26752 12767
rect 26700 12724 26752 12733
rect 27436 12724 27488 12776
rect 23480 12699 23532 12708
rect 23480 12665 23489 12699
rect 23489 12665 23523 12699
rect 23523 12665 23532 12699
rect 23480 12656 23532 12665
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 18328 12631 18380 12640
rect 18328 12597 18337 12631
rect 18337 12597 18371 12631
rect 18371 12597 18380 12631
rect 18328 12588 18380 12597
rect 24308 12656 24360 12708
rect 25688 12631 25740 12640
rect 25688 12597 25697 12631
rect 25697 12597 25731 12631
rect 25731 12597 25740 12631
rect 25688 12588 25740 12597
rect 25872 12656 25924 12708
rect 27528 12656 27580 12708
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 5540 12384 5592 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8208 12384 8260 12436
rect 13084 12384 13136 12436
rect 13360 12384 13412 12436
rect 17316 12384 17368 12436
rect 23848 12427 23900 12436
rect 23848 12393 23857 12427
rect 23857 12393 23891 12427
rect 23891 12393 23900 12427
rect 23848 12384 23900 12393
rect 24860 12427 24912 12436
rect 24860 12393 24869 12427
rect 24869 12393 24903 12427
rect 24903 12393 24912 12427
rect 24860 12384 24912 12393
rect 25320 12427 25372 12436
rect 25320 12393 25329 12427
rect 25329 12393 25363 12427
rect 25363 12393 25372 12427
rect 25320 12384 25372 12393
rect 25688 12384 25740 12436
rect 27436 12384 27488 12436
rect 16488 12316 16540 12368
rect 21272 12316 21324 12368
rect 25596 12316 25648 12368
rect 26148 12316 26200 12368
rect 4988 12291 5040 12300
rect 4988 12257 4997 12291
rect 4997 12257 5031 12291
rect 5031 12257 5040 12291
rect 4988 12248 5040 12257
rect 5448 12248 5500 12300
rect 13452 12248 13504 12300
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 21916 12248 21968 12300
rect 22744 12248 22796 12300
rect 23848 12248 23900 12300
rect 26516 12291 26568 12300
rect 26516 12257 26525 12291
rect 26525 12257 26559 12291
rect 26559 12257 26568 12291
rect 26516 12248 26568 12257
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 17132 12180 17184 12232
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 24952 12180 25004 12232
rect 25136 12180 25188 12232
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9680 12044 9732 12096
rect 10140 12044 10192 12096
rect 10876 12044 10928 12096
rect 11152 12044 11204 12096
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 17224 12044 17276 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 21824 12044 21876 12096
rect 26332 12044 26384 12096
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 5080 11840 5132 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 12716 11840 12768 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 21272 11883 21324 11892
rect 17500 11840 17552 11849
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 5172 11704 5224 11756
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13360 11704 13412 11756
rect 4252 11636 4304 11688
rect 4528 11636 4580 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 7380 11636 7432 11688
rect 10508 11636 10560 11688
rect 2688 11568 2740 11620
rect 3976 11568 4028 11620
rect 5264 11568 5316 11620
rect 7196 11611 7248 11620
rect 7196 11577 7205 11611
rect 7205 11577 7239 11611
rect 7239 11577 7248 11611
rect 7196 11568 7248 11577
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 7840 11500 7892 11552
rect 12348 11568 12400 11620
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 24952 11883 25004 11892
rect 24952 11849 24961 11883
rect 24961 11849 24995 11883
rect 24995 11849 25004 11883
rect 24952 11840 25004 11849
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 25596 11883 25648 11892
rect 25596 11849 25605 11883
rect 25605 11849 25639 11883
rect 25639 11849 25648 11883
rect 25596 11840 25648 11849
rect 26516 11840 26568 11892
rect 13912 11704 13964 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 17960 11636 18012 11688
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 17776 11568 17828 11620
rect 19156 11611 19208 11620
rect 19156 11577 19165 11611
rect 19165 11577 19199 11611
rect 19199 11577 19208 11611
rect 19156 11568 19208 11577
rect 11336 11500 11388 11552
rect 12992 11500 13044 11552
rect 13636 11500 13688 11552
rect 17132 11543 17184 11552
rect 17132 11509 17141 11543
rect 17141 11509 17175 11543
rect 17175 11509 17184 11543
rect 17132 11500 17184 11509
rect 19064 11500 19116 11552
rect 21916 11500 21968 11552
rect 26608 11543 26660 11552
rect 26608 11509 26617 11543
rect 26617 11509 26651 11543
rect 26651 11509 26660 11543
rect 26608 11500 26660 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 12348 11296 12400 11348
rect 13360 11296 13412 11348
rect 13636 11296 13688 11348
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 14372 11296 14424 11348
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 17224 11271 17276 11280
rect 17224 11237 17233 11271
rect 17233 11237 17267 11271
rect 17267 11237 17276 11271
rect 17224 11228 17276 11237
rect 2044 11160 2096 11212
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 21916 11160 21968 11212
rect 22836 11160 22888 11212
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 4160 11092 4212 11144
rect 5264 11092 5316 11144
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 14280 11135 14332 11144
rect 7840 11092 7892 11101
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 16948 11092 17000 11144
rect 18512 11092 18564 11144
rect 19064 11135 19116 11144
rect 19064 11101 19073 11135
rect 19073 11101 19107 11135
rect 19107 11101 19116 11135
rect 19064 11092 19116 11101
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 7564 11024 7616 11076
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 13728 11024 13780 11076
rect 16856 11067 16908 11076
rect 16856 11033 16865 11067
rect 16865 11033 16899 11067
rect 16899 11033 16908 11067
rect 16856 11024 16908 11033
rect 17776 11024 17828 11076
rect 22192 10956 22244 11008
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1492 10752 1544 10804
rect 2044 10795 2096 10804
rect 2044 10761 2053 10795
rect 2053 10761 2087 10795
rect 2087 10761 2096 10795
rect 2044 10752 2096 10761
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 3424 10752 3476 10804
rect 4068 10752 4120 10804
rect 7840 10752 7892 10804
rect 14280 10752 14332 10804
rect 17316 10795 17368 10804
rect 17316 10761 17325 10795
rect 17325 10761 17359 10795
rect 17359 10761 17368 10795
rect 17316 10752 17368 10761
rect 17776 10795 17828 10804
rect 17776 10761 17785 10795
rect 17785 10761 17819 10795
rect 17819 10761 17828 10795
rect 17776 10752 17828 10761
rect 18788 10752 18840 10804
rect 20720 10752 20772 10804
rect 22836 10795 22888 10804
rect 4436 10727 4488 10736
rect 4436 10693 4445 10727
rect 4445 10693 4479 10727
rect 4479 10693 4488 10727
rect 4436 10684 4488 10693
rect 7748 10727 7800 10736
rect 7748 10693 7757 10727
rect 7757 10693 7791 10727
rect 7791 10693 7800 10727
rect 7748 10684 7800 10693
rect 17224 10684 17276 10736
rect 17868 10684 17920 10736
rect 20628 10684 20680 10736
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 5172 10616 5224 10668
rect 7656 10616 7708 10668
rect 22836 10761 22845 10795
rect 22845 10761 22879 10795
rect 22879 10761 22888 10795
rect 22836 10752 22888 10761
rect 26516 10795 26568 10804
rect 26516 10761 26525 10795
rect 26525 10761 26559 10795
rect 26559 10761 26568 10795
rect 26516 10752 26568 10761
rect 2412 10548 2464 10600
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 23388 10616 23440 10668
rect 13636 10548 13688 10600
rect 18880 10548 18932 10600
rect 24216 10591 24268 10600
rect 24216 10557 24225 10591
rect 24225 10557 24259 10591
rect 24259 10557 24268 10591
rect 24216 10548 24268 10557
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 16948 10455 17000 10464
rect 4896 10412 4948 10421
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 20720 10412 20772 10464
rect 22192 10455 22244 10464
rect 22192 10421 22201 10455
rect 22201 10421 22235 10455
rect 22235 10421 22244 10455
rect 22192 10412 22244 10421
rect 22284 10455 22336 10464
rect 22284 10421 22293 10455
rect 22293 10421 22327 10455
rect 22327 10421 22336 10455
rect 22284 10412 22336 10421
rect 23572 10412 23624 10464
rect 25596 10455 25648 10464
rect 25596 10421 25605 10455
rect 25605 10421 25639 10455
rect 25639 10421 25648 10455
rect 25596 10412 25648 10421
rect 26608 10412 26660 10464
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2688 10208 2740 10260
rect 2780 10208 2832 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 14372 10208 14424 10260
rect 18972 10208 19024 10260
rect 21824 10208 21876 10260
rect 22284 10208 22336 10260
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 24860 10251 24912 10260
rect 24860 10217 24869 10251
rect 24869 10217 24903 10251
rect 24903 10217 24912 10251
rect 24860 10208 24912 10217
rect 25320 10251 25372 10260
rect 25320 10217 25329 10251
rect 25329 10217 25363 10251
rect 25363 10217 25372 10251
rect 25320 10208 25372 10217
rect 26976 10251 27028 10260
rect 26976 10217 26985 10251
rect 26985 10217 27019 10251
rect 27019 10217 27028 10251
rect 26976 10208 27028 10217
rect 4988 10140 5040 10192
rect 12992 10140 13044 10192
rect 2228 10072 2280 10124
rect 4068 10072 4120 10124
rect 5172 10072 5224 10124
rect 10232 10115 10284 10124
rect 10232 10081 10241 10115
rect 10241 10081 10275 10115
rect 10275 10081 10284 10115
rect 10232 10072 10284 10081
rect 10876 10072 10928 10124
rect 5448 10004 5500 10056
rect 2136 9868 2188 9920
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 3516 9911 3568 9920
rect 2780 9868 2832 9877
rect 3516 9877 3525 9911
rect 3525 9877 3559 9911
rect 3559 9877 3568 9911
rect 3516 9868 3568 9877
rect 6920 9868 6972 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 11612 9911 11664 9920
rect 11612 9877 11621 9911
rect 11621 9877 11655 9911
rect 11655 9877 11664 9911
rect 11612 9868 11664 9877
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 13912 10140 13964 10192
rect 14280 10140 14332 10192
rect 18420 10140 18472 10192
rect 18788 10140 18840 10192
rect 14004 10072 14056 10124
rect 15844 10115 15896 10124
rect 15844 10081 15878 10115
rect 15878 10081 15896 10115
rect 15844 10072 15896 10081
rect 20628 10115 20680 10124
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 22744 10115 22796 10124
rect 22744 10081 22753 10115
rect 22753 10081 22787 10115
rect 22787 10081 22796 10115
rect 22744 10072 22796 10081
rect 25688 10072 25740 10124
rect 26884 10115 26936 10124
rect 26884 10081 26893 10115
rect 26893 10081 26927 10115
rect 26927 10081 26936 10115
rect 26884 10072 26936 10081
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 19156 10004 19208 10056
rect 22836 10047 22888 10056
rect 22836 10013 22845 10047
rect 22845 10013 22879 10047
rect 22879 10013 22888 10047
rect 22836 10004 22888 10013
rect 22928 10047 22980 10056
rect 22928 10013 22937 10047
rect 22937 10013 22971 10047
rect 22971 10013 22980 10047
rect 22928 10004 22980 10013
rect 24860 10004 24912 10056
rect 25596 10004 25648 10056
rect 18144 9979 18196 9988
rect 18144 9945 18153 9979
rect 18153 9945 18187 9979
rect 18187 9945 18196 9979
rect 18144 9936 18196 9945
rect 12440 9868 12492 9877
rect 13636 9868 13688 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17408 9868 17460 9920
rect 17868 9868 17920 9920
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 18512 9868 18564 9920
rect 19800 9868 19852 9920
rect 20168 9868 20220 9920
rect 20444 9911 20496 9920
rect 20444 9877 20453 9911
rect 20453 9877 20487 9911
rect 20487 9877 20496 9911
rect 20444 9868 20496 9877
rect 21916 9868 21968 9920
rect 24216 9936 24268 9988
rect 23572 9868 23624 9920
rect 26424 9868 26476 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2228 9664 2280 9716
rect 3424 9707 3476 9716
rect 3424 9673 3433 9707
rect 3433 9673 3467 9707
rect 3467 9673 3476 9707
rect 3424 9664 3476 9673
rect 4712 9664 4764 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 15844 9664 15896 9716
rect 17776 9664 17828 9716
rect 18972 9664 19024 9716
rect 20628 9664 20680 9716
rect 22928 9664 22980 9716
rect 24860 9707 24912 9716
rect 24860 9673 24869 9707
rect 24869 9673 24903 9707
rect 24903 9673 24912 9707
rect 24860 9664 24912 9673
rect 25320 9707 25372 9716
rect 25320 9673 25329 9707
rect 25329 9673 25363 9707
rect 25363 9673 25372 9707
rect 25320 9664 25372 9673
rect 26884 9707 26936 9716
rect 26884 9673 26893 9707
rect 26893 9673 26927 9707
rect 26927 9673 26936 9707
rect 26884 9664 26936 9673
rect 26976 9664 27028 9716
rect 2780 9528 2832 9580
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 3516 9460 3568 9512
rect 4620 9460 4672 9512
rect 2044 9435 2096 9444
rect 2044 9401 2053 9435
rect 2053 9401 2087 9435
rect 2087 9401 2096 9435
rect 2044 9392 2096 9401
rect 3608 9392 3660 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4068 9324 4120 9376
rect 4804 9596 4856 9648
rect 12164 9639 12216 9648
rect 5448 9528 5500 9580
rect 5908 9528 5960 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 12164 9605 12173 9639
rect 12173 9605 12207 9639
rect 12207 9605 12216 9639
rect 12164 9596 12216 9605
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 12440 9528 12492 9580
rect 10416 9460 10468 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 22744 9596 22796 9648
rect 25780 9639 25832 9648
rect 25780 9605 25789 9639
rect 25789 9605 25823 9639
rect 25823 9605 25832 9639
rect 25780 9596 25832 9605
rect 19064 9528 19116 9580
rect 19156 9528 19208 9580
rect 20352 9528 20404 9580
rect 21824 9528 21876 9580
rect 23572 9528 23624 9580
rect 26424 9571 26476 9580
rect 26424 9537 26433 9571
rect 26433 9537 26467 9571
rect 26467 9537 26476 9571
rect 26424 9528 26476 9537
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 18144 9460 18196 9512
rect 19800 9460 19852 9512
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 5724 9324 5776 9376
rect 12164 9392 12216 9444
rect 12900 9435 12952 9444
rect 12900 9401 12909 9435
rect 12909 9401 12943 9435
rect 12943 9401 12952 9435
rect 12900 9392 12952 9401
rect 15016 9392 15068 9444
rect 20536 9392 20588 9444
rect 21548 9392 21600 9444
rect 23848 9460 23900 9512
rect 25964 9460 26016 9512
rect 26608 9460 26660 9512
rect 26884 9460 26936 9512
rect 23664 9392 23716 9444
rect 25780 9392 25832 9444
rect 8392 9324 8444 9376
rect 12256 9324 12308 9376
rect 12532 9324 12584 9376
rect 15108 9324 15160 9376
rect 15568 9324 15620 9376
rect 16672 9324 16724 9376
rect 17868 9324 17920 9376
rect 18236 9324 18288 9376
rect 19708 9367 19760 9376
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21456 9367 21508 9376
rect 21456 9333 21465 9367
rect 21465 9333 21499 9367
rect 21499 9333 21508 9367
rect 21456 9324 21508 9333
rect 23756 9324 23808 9376
rect 24216 9324 24268 9376
rect 25688 9324 25740 9376
rect 27620 9367 27672 9376
rect 27620 9333 27629 9367
rect 27629 9333 27663 9367
rect 27663 9333 27672 9367
rect 27620 9324 27672 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 2136 9120 2188 9172
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 4436 9120 4488 9172
rect 4988 9120 5040 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 6920 9163 6972 9172
rect 6920 9129 6929 9163
rect 6929 9129 6963 9163
rect 6963 9129 6972 9163
rect 6920 9120 6972 9129
rect 10784 9120 10836 9172
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 16856 9120 16908 9172
rect 17868 9163 17920 9172
rect 17868 9129 17877 9163
rect 17877 9129 17911 9163
rect 17911 9129 17920 9163
rect 17868 9120 17920 9129
rect 19892 9120 19944 9172
rect 20352 9163 20404 9172
rect 20352 9129 20361 9163
rect 20361 9129 20395 9163
rect 20395 9129 20404 9163
rect 20352 9120 20404 9129
rect 21548 9163 21600 9172
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 22836 9120 22888 9172
rect 25688 9120 25740 9172
rect 25964 9163 26016 9172
rect 25964 9129 25973 9163
rect 25973 9129 26007 9163
rect 26007 9129 26016 9163
rect 25964 9120 26016 9129
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 2412 9052 2464 9104
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 4620 8984 4672 9036
rect 6644 8984 6696 9036
rect 8116 8984 8168 9036
rect 18788 9095 18840 9104
rect 18788 9061 18797 9095
rect 18797 9061 18831 9095
rect 18831 9061 18840 9095
rect 18788 9052 18840 9061
rect 20076 9052 20128 9104
rect 21456 9052 21508 9104
rect 22744 9095 22796 9104
rect 22744 9061 22753 9095
rect 22753 9061 22787 9095
rect 22787 9061 22796 9095
rect 22744 9052 22796 9061
rect 23204 9052 23256 9104
rect 26424 9052 26476 9104
rect 26976 9052 27028 9104
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 18236 8984 18288 9036
rect 19156 8984 19208 9036
rect 23388 9027 23440 9036
rect 23388 8993 23397 9027
rect 23397 8993 23431 9027
rect 23431 8993 23440 9027
rect 23388 8984 23440 8993
rect 23848 8984 23900 9036
rect 24032 8984 24084 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 3424 8916 3476 8968
rect 5448 8916 5500 8968
rect 6920 8916 6972 8968
rect 11980 8916 12032 8968
rect 12440 8916 12492 8968
rect 17408 8916 17460 8968
rect 19064 8916 19116 8968
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 9404 8780 9456 8832
rect 9680 8780 9732 8832
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 11152 8780 11204 8832
rect 13636 8780 13688 8832
rect 14004 8823 14056 8832
rect 14004 8789 14013 8823
rect 14013 8789 14047 8823
rect 14047 8789 14056 8823
rect 14004 8780 14056 8789
rect 16948 8780 17000 8832
rect 24124 8823 24176 8832
rect 24124 8789 24133 8823
rect 24133 8789 24167 8823
rect 24167 8789 24176 8823
rect 24124 8780 24176 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 9128 8576 9180 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 19064 8576 19116 8628
rect 19892 8576 19944 8628
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 26516 8576 26568 8628
rect 1400 8508 1452 8560
rect 2228 8508 2280 8560
rect 3424 8551 3476 8560
rect 3424 8517 3433 8551
rect 3433 8517 3467 8551
rect 3467 8517 3476 8551
rect 3424 8508 3476 8517
rect 4436 8508 4488 8560
rect 5448 8508 5500 8560
rect 6920 8508 6972 8560
rect 9496 8508 9548 8560
rect 2504 8440 2556 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 8392 8440 8444 8492
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 11152 8483 11204 8492
rect 11152 8449 11161 8483
rect 11161 8449 11195 8483
rect 11195 8449 11204 8483
rect 11152 8440 11204 8449
rect 16304 8508 16356 8560
rect 23572 8508 23624 8560
rect 26976 8551 27028 8560
rect 26976 8517 26985 8551
rect 26985 8517 27019 8551
rect 27019 8517 27028 8551
rect 26976 8508 27028 8517
rect 11612 8440 11664 8492
rect 12532 8440 12584 8492
rect 2044 8372 2096 8424
rect 9128 8372 9180 8424
rect 9404 8415 9456 8424
rect 9404 8381 9413 8415
rect 9413 8381 9447 8415
rect 9447 8381 9456 8415
rect 9404 8372 9456 8381
rect 12256 8372 12308 8424
rect 17868 8440 17920 8492
rect 22652 8440 22704 8492
rect 23940 8440 23992 8492
rect 24124 8440 24176 8492
rect 16856 8372 16908 8424
rect 6092 8304 6144 8356
rect 7104 8304 7156 8356
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 7840 8279 7892 8288
rect 7840 8245 7849 8279
rect 7849 8245 7883 8279
rect 7883 8245 7892 8279
rect 8944 8279 8996 8288
rect 7840 8236 7892 8245
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 11980 8304 12032 8356
rect 16212 8347 16264 8356
rect 16212 8313 16221 8347
rect 16221 8313 16255 8347
rect 16255 8313 16264 8347
rect 16212 8304 16264 8313
rect 16488 8304 16540 8356
rect 16948 8304 17000 8356
rect 23940 8304 23992 8356
rect 25596 8415 25648 8424
rect 25596 8381 25605 8415
rect 25605 8381 25639 8415
rect 25639 8381 25648 8415
rect 25596 8372 25648 8381
rect 24584 8304 24636 8356
rect 24676 8304 24728 8356
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 23480 8236 23532 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 2136 8032 2188 8084
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 7840 8032 7892 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9864 8032 9916 8084
rect 10876 8032 10928 8084
rect 4896 8007 4948 8016
rect 4896 7973 4905 8007
rect 4905 7973 4939 8007
rect 4939 7973 4948 8007
rect 4896 7964 4948 7973
rect 8944 7964 8996 8016
rect 1676 7896 1728 7948
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 7288 7896 7340 7948
rect 10600 7896 10652 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 8116 7828 8168 7880
rect 9496 7828 9548 7880
rect 9588 7828 9640 7880
rect 12440 8032 12492 8084
rect 14740 8032 14792 8084
rect 15016 8032 15068 8084
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 17960 8032 18012 8084
rect 20076 8032 20128 8084
rect 23204 8032 23256 8084
rect 24768 8032 24820 8084
rect 25596 8075 25648 8084
rect 25596 8041 25605 8075
rect 25605 8041 25639 8075
rect 25639 8041 25648 8075
rect 25596 8032 25648 8041
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 11888 7896 11940 7948
rect 12624 7964 12676 8016
rect 13636 7964 13688 8016
rect 12348 7939 12400 7948
rect 12348 7905 12382 7939
rect 12382 7905 12400 7939
rect 12348 7896 12400 7905
rect 16672 7939 16724 7948
rect 16672 7905 16681 7939
rect 16681 7905 16715 7939
rect 16715 7905 16724 7939
rect 16672 7896 16724 7905
rect 16764 7896 16816 7948
rect 17408 7896 17460 7948
rect 20444 7896 20496 7948
rect 21272 7939 21324 7948
rect 21272 7905 21281 7939
rect 21281 7905 21315 7939
rect 21315 7905 21324 7939
rect 21272 7896 21324 7905
rect 23112 7896 23164 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 23296 7828 23348 7880
rect 23848 7828 23900 7880
rect 24676 7828 24728 7880
rect 4620 7760 4672 7812
rect 7012 7760 7064 7812
rect 19524 7760 19576 7812
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 5172 7692 5224 7744
rect 19156 7735 19208 7744
rect 19156 7701 19165 7735
rect 19165 7701 19199 7735
rect 19199 7701 19208 7735
rect 19156 7692 19208 7701
rect 20352 7692 20404 7744
rect 20812 7692 20864 7744
rect 21548 7692 21600 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2504 7488 2556 7540
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 4988 7488 5040 7540
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8484 7531 8536 7540
rect 8484 7497 8493 7531
rect 8493 7497 8527 7531
rect 8527 7497 8536 7531
rect 8484 7488 8536 7497
rect 8944 7488 8996 7540
rect 9588 7488 9640 7540
rect 9864 7488 9916 7540
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 4896 7420 4948 7472
rect 16672 7420 16724 7472
rect 2136 7352 2188 7404
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 12348 7352 12400 7404
rect 12440 7352 12492 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 4528 7284 4580 7336
rect 10508 7284 10560 7336
rect 20352 7284 20404 7336
rect 2504 7259 2556 7268
rect 2504 7225 2538 7259
rect 2538 7225 2556 7259
rect 2504 7216 2556 7225
rect 10324 7216 10376 7268
rect 14280 7216 14332 7268
rect 15108 7216 15160 7268
rect 19156 7216 19208 7268
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 19248 7148 19300 7200
rect 20444 7191 20496 7200
rect 20444 7157 20453 7191
rect 20453 7157 20487 7191
rect 20487 7157 20496 7191
rect 20444 7148 20496 7157
rect 20628 7148 20680 7200
rect 23112 7531 23164 7540
rect 23112 7497 23121 7531
rect 23121 7497 23155 7531
rect 23155 7497 23164 7531
rect 23112 7488 23164 7497
rect 23480 7488 23532 7540
rect 26608 7531 26660 7540
rect 26608 7497 26617 7531
rect 26617 7497 26651 7531
rect 26651 7497 26660 7531
rect 26608 7488 26660 7497
rect 26516 7420 26568 7472
rect 27712 7463 27764 7472
rect 27712 7429 27721 7463
rect 27721 7429 27755 7463
rect 27755 7429 27764 7463
rect 27712 7420 27764 7429
rect 24676 7352 24728 7404
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24032 7284 24084 7293
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 27528 7327 27580 7336
rect 27528 7293 27537 7327
rect 27537 7293 27571 7327
rect 27571 7293 27580 7327
rect 27528 7284 27580 7293
rect 21364 7216 21416 7268
rect 23848 7216 23900 7268
rect 25136 7216 25188 7268
rect 21456 7148 21508 7200
rect 23756 7148 23808 7200
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 2504 6944 2556 6996
rect 5080 6944 5132 6996
rect 10600 6944 10652 6996
rect 15660 6987 15712 6996
rect 15660 6953 15669 6987
rect 15669 6953 15703 6987
rect 15703 6953 15712 6987
rect 15660 6944 15712 6953
rect 19800 6944 19852 6996
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 24032 6987 24084 6996
rect 24032 6953 24041 6987
rect 24041 6953 24075 6987
rect 24075 6953 24084 6987
rect 24032 6944 24084 6953
rect 1860 6808 1912 6860
rect 5172 6851 5224 6860
rect 5172 6817 5206 6851
rect 5206 6817 5224 6851
rect 5172 6808 5224 6817
rect 5540 6808 5592 6860
rect 7012 6876 7064 6928
rect 10324 6808 10376 6860
rect 13636 6808 13688 6860
rect 14004 6851 14056 6860
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 14188 6808 14240 6860
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 15292 6740 15344 6792
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16120 6808 16172 6860
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 19524 6876 19576 6928
rect 21364 6876 21416 6928
rect 21180 6808 21232 6860
rect 17224 6740 17276 6792
rect 26332 6808 26384 6860
rect 27344 6808 27396 6860
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 5080 6604 5132 6656
rect 5264 6604 5316 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 9312 6604 9364 6656
rect 15016 6604 15068 6656
rect 17684 6672 17736 6724
rect 20720 6672 20772 6724
rect 20996 6672 21048 6724
rect 21824 6672 21876 6724
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 15752 6604 15804 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 23756 6647 23808 6656
rect 23756 6613 23765 6647
rect 23765 6613 23799 6647
rect 23799 6613 23808 6647
rect 23756 6604 23808 6613
rect 24676 6604 24728 6656
rect 25320 6604 25372 6656
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1860 6400 1912 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 14280 6400 14332 6452
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 17316 6400 17368 6452
rect 20996 6443 21048 6452
rect 5172 6332 5224 6384
rect 9680 6332 9732 6384
rect 17224 6332 17276 6384
rect 3608 6264 3660 6316
rect 6276 6264 6328 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 10508 6264 10560 6316
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 4712 6196 4764 6248
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 9128 6239 9180 6248
rect 8668 6196 8720 6205
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10324 6196 10376 6248
rect 15108 6264 15160 6316
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 21272 6443 21324 6452
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 26608 6375 26660 6384
rect 26608 6341 26617 6375
rect 26617 6341 26651 6375
rect 26651 6341 26660 6375
rect 26608 6332 26660 6341
rect 15292 6264 15344 6273
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 22928 6196 22980 6248
rect 24768 6196 24820 6248
rect 27160 6400 27212 6452
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 8852 6128 8904 6180
rect 10140 6128 10192 6180
rect 14556 6128 14608 6180
rect 16764 6171 16816 6180
rect 16764 6137 16773 6171
rect 16773 6137 16807 6171
rect 16807 6137 16816 6171
rect 16764 6128 16816 6137
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 2688 6060 2740 6112
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 4252 6060 4304 6112
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 21272 6060 21324 6112
rect 23480 6103 23532 6112
rect 23480 6069 23489 6103
rect 23489 6069 23523 6103
rect 23523 6069 23532 6103
rect 23480 6060 23532 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2780 5856 2832 5908
rect 2872 5856 2924 5908
rect 3792 5856 3844 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 12440 5856 12492 5908
rect 15752 5856 15804 5908
rect 16856 5856 16908 5908
rect 16948 5856 17000 5908
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 19708 5899 19760 5908
rect 19708 5865 19717 5899
rect 19717 5865 19751 5899
rect 19751 5865 19760 5899
rect 19708 5856 19760 5865
rect 23480 5856 23532 5908
rect 2596 5831 2648 5840
rect 2596 5797 2605 5831
rect 2605 5797 2639 5831
rect 2639 5797 2648 5831
rect 2596 5788 2648 5797
rect 6276 5831 6328 5840
rect 6276 5797 6310 5831
rect 6310 5797 6328 5831
rect 6276 5788 6328 5797
rect 2412 5720 2464 5772
rect 2504 5652 2556 5704
rect 5540 5720 5592 5772
rect 11888 5788 11940 5840
rect 16396 5788 16448 5840
rect 17132 5831 17184 5840
rect 17132 5797 17141 5831
rect 17141 5797 17175 5831
rect 17175 5797 17184 5831
rect 17132 5788 17184 5797
rect 19340 5788 19392 5840
rect 11520 5720 11572 5772
rect 20720 5720 20772 5772
rect 21916 5720 21968 5772
rect 16764 5652 16816 5704
rect 19892 5695 19944 5704
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 22928 5788 22980 5840
rect 26792 5720 26844 5772
rect 21456 5652 21508 5661
rect 8852 5627 8904 5636
rect 8852 5593 8861 5627
rect 8861 5593 8895 5627
rect 8895 5593 8904 5627
rect 8852 5584 8904 5593
rect 26700 5627 26752 5636
rect 26700 5593 26709 5627
rect 26709 5593 26743 5627
rect 26743 5593 26752 5627
rect 26700 5584 26752 5593
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 14556 5516 14608 5568
rect 14924 5516 14976 5568
rect 15292 5516 15344 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 21272 5516 21324 5568
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 6276 5312 6328 5364
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 15108 5312 15160 5364
rect 16764 5355 16816 5364
rect 16764 5321 16773 5355
rect 16773 5321 16807 5355
rect 16807 5321 16816 5355
rect 16764 5312 16816 5321
rect 16948 5312 17000 5364
rect 19156 5312 19208 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 20260 5312 20312 5364
rect 20720 5312 20772 5364
rect 21456 5312 21508 5364
rect 2596 5244 2648 5296
rect 5540 5244 5592 5296
rect 6736 5244 6788 5296
rect 17132 5287 17184 5296
rect 17132 5253 17141 5287
rect 17141 5253 17175 5287
rect 17175 5253 17184 5287
rect 17132 5244 17184 5253
rect 19892 5244 19944 5296
rect 21916 5312 21968 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 26792 5312 26844 5364
rect 3700 5176 3752 5228
rect 8760 5176 8812 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 4712 5108 4764 5160
rect 9588 5108 9640 5160
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 20720 5108 20772 5160
rect 21732 5108 21784 5160
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 14924 5040 14976 5092
rect 21364 5040 21416 5092
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 3608 4972 3660 4981
rect 3976 4972 4028 5024
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 11428 5015 11480 5024
rect 11428 4981 11437 5015
rect 11437 4981 11471 5015
rect 11471 4981 11480 5015
rect 11428 4972 11480 4981
rect 20260 4972 20312 5024
rect 21732 4972 21784 5024
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 1400 4768 1452 4820
rect 2688 4768 2740 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4252 4768 4304 4820
rect 5540 4768 5592 4820
rect 7380 4768 7432 4820
rect 8576 4768 8628 4820
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 11428 4768 11480 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 21364 4768 21416 4820
rect 11612 4700 11664 4752
rect 11888 4700 11940 4752
rect 16764 4743 16816 4752
rect 16764 4709 16798 4743
rect 16798 4709 16816 4743
rect 16764 4700 16816 4709
rect 21180 4700 21232 4752
rect 21548 4700 21600 4752
rect 2412 4632 2464 4684
rect 2596 4632 2648 4684
rect 4620 4632 4672 4684
rect 14188 4675 14240 4684
rect 14188 4641 14197 4675
rect 14197 4641 14231 4675
rect 14231 4641 14240 4675
rect 14188 4632 14240 4641
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 20812 4496 20864 4548
rect 20996 4496 21048 4548
rect 21272 4496 21324 4548
rect 21916 4496 21968 4548
rect 4160 4428 4212 4480
rect 6828 4428 6880 4480
rect 16856 4428 16908 4480
rect 17868 4471 17920 4480
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 2872 4224 2924 4276
rect 3700 4267 3752 4276
rect 3700 4233 3709 4267
rect 3709 4233 3743 4267
rect 3743 4233 3752 4267
rect 3700 4224 3752 4233
rect 5264 4224 5316 4276
rect 8484 4224 8536 4276
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 21180 4224 21232 4276
rect 26516 4224 26568 4276
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3240 4088 3292 4140
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 3700 4020 3752 4072
rect 4252 4063 4304 4072
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 5540 4088 5592 4140
rect 4528 4063 4580 4072
rect 4528 4029 4551 4063
rect 4551 4029 4580 4063
rect 4528 4020 4580 4029
rect 4620 3952 4672 4004
rect 7380 4088 7432 4140
rect 8576 4156 8628 4208
rect 9680 4156 9732 4208
rect 10508 4156 10560 4208
rect 9220 4088 9272 4140
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 8760 4020 8812 4072
rect 10324 4020 10376 4072
rect 11336 4088 11388 4140
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 16856 4088 16908 4140
rect 20996 4156 21048 4208
rect 7472 3952 7524 4004
rect 9128 3952 9180 4004
rect 14648 4020 14700 4072
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15016 4020 15068 4029
rect 16672 4020 16724 4072
rect 20352 4020 20404 4072
rect 22928 4156 22980 4208
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 5172 3884 5224 3936
rect 7196 3884 7248 3936
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 21272 3995 21324 4004
rect 21272 3961 21306 3995
rect 21306 3961 21324 3995
rect 21272 3952 21324 3961
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 16580 3884 16632 3936
rect 18144 3884 18196 3936
rect 21916 3884 21968 3936
rect 26792 3884 26844 3936
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1400 3680 1452 3732
rect 2964 3680 3016 3732
rect 3056 3680 3108 3732
rect 4528 3680 4580 3732
rect 7288 3680 7340 3732
rect 9128 3723 9180 3732
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 10324 3680 10376 3732
rect 11612 3680 11664 3732
rect 15016 3680 15068 3732
rect 16672 3680 16724 3732
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 20812 3680 20864 3732
rect 21364 3723 21416 3732
rect 21364 3689 21373 3723
rect 21373 3689 21407 3723
rect 21407 3689 21416 3723
rect 21364 3680 21416 3689
rect 7380 3655 7432 3664
rect 7380 3621 7414 3655
rect 7414 3621 7432 3655
rect 7380 3612 7432 3621
rect 3608 3544 3660 3596
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 6736 3544 6788 3596
rect 7012 3544 7064 3596
rect 11520 3612 11572 3664
rect 11888 3612 11940 3664
rect 16764 3612 16816 3664
rect 17960 3612 18012 3664
rect 21640 3612 21692 3664
rect 11336 3587 11388 3596
rect 11336 3553 11370 3587
rect 11370 3553 11388 3587
rect 11336 3544 11388 3553
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 24860 3544 24912 3596
rect 25320 3587 25372 3596
rect 25320 3553 25329 3587
rect 25329 3553 25363 3587
rect 25363 3553 25372 3587
rect 25320 3544 25372 3553
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 2872 3476 2924 3528
rect 3240 3476 3292 3528
rect 3792 3476 3844 3528
rect 3976 3408 4028 3460
rect 9588 3408 9640 3460
rect 21272 3408 21324 3460
rect 25504 3451 25556 3460
rect 25504 3417 25513 3451
rect 25513 3417 25547 3451
rect 25547 3417 25556 3451
rect 25504 3408 25556 3417
rect 2596 3340 2648 3392
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2780 3136 2832 3188
rect 3332 3136 3384 3188
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5172 3136 5224 3188
rect 7380 3136 7432 3188
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 11336 3136 11388 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 17960 3136 18012 3188
rect 7196 3068 7248 3120
rect 3792 3000 3844 3052
rect 18144 3068 18196 3120
rect 9588 3000 9640 3052
rect 2964 2932 3016 2984
rect 4804 2932 4856 2984
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 9036 2932 9088 2984
rect 10140 2932 10192 2984
rect 13544 2932 13596 2984
rect 20536 3136 20588 3188
rect 21364 3136 21416 3188
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 24308 3136 24360 3188
rect 25320 3179 25372 3188
rect 25320 3145 25329 3179
rect 25329 3145 25363 3179
rect 25363 3145 25372 3179
rect 25320 3136 25372 3145
rect 26516 3136 26568 3188
rect 24308 2932 24360 2984
rect 27252 3068 27304 3120
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 2044 2796 2096 2848
rect 7748 2864 7800 2916
rect 12072 2864 12124 2916
rect 14924 2864 14976 2916
rect 20628 2864 20680 2916
rect 24860 2864 24912 2916
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 27804 2796 27856 2848
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 2688 2635 2740 2644
rect 2688 2601 2697 2635
rect 2697 2601 2731 2635
rect 2731 2601 2740 2635
rect 2688 2592 2740 2601
rect 2780 2592 2832 2644
rect 2964 2524 3016 2576
rect 3700 2524 3752 2576
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 6828 2592 6880 2644
rect 7012 2592 7064 2644
rect 9588 2592 9640 2644
rect 19248 2635 19300 2644
rect 19248 2601 19257 2635
rect 19257 2601 19291 2635
rect 19291 2601 19300 2635
rect 19248 2592 19300 2601
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 10692 2456 10744 2508
rect 13820 2456 13872 2508
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 20812 2592 20864 2644
rect 21272 2592 21324 2644
rect 22100 2456 22152 2508
rect 24308 2499 24360 2508
rect 24308 2465 24317 2499
rect 24317 2465 24351 2499
rect 24351 2465 24360 2499
rect 24308 2456 24360 2465
rect 25136 2456 25188 2508
rect 4896 2388 4948 2440
rect 6368 2388 6420 2440
rect 9220 2388 9272 2440
rect 10600 2388 10652 2440
rect 13452 2388 13504 2440
rect 16304 2388 16356 2440
rect 17776 2388 17828 2440
rect 19156 2388 19208 2440
rect 22008 2388 22060 2440
rect 23480 2388 23532 2440
rect 26332 2388 26384 2440
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 29184 2252 29236 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 3330 23624 3386 23633
rect 3330 23559 3386 23568
rect 2410 22400 2466 22409
rect 2410 22335 2466 22344
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18222 1532 18566
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 10441 1440 15846
rect 1504 15570 1532 18158
rect 1780 17882 1808 18702
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 2318 17776 2374 17785
rect 2318 17711 2320 17720
rect 2372 17711 2374 17720
rect 2320 17682 2372 17688
rect 2332 17626 2360 17682
rect 2240 17598 2360 17626
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1688 16794 1716 17274
rect 1780 17202 1808 17478
rect 2240 17338 2268 17598
rect 2320 17536 2372 17542
rect 2424 17513 2452 22335
rect 3054 21856 3110 21865
rect 3054 21791 3110 21800
rect 2870 21312 2926 21321
rect 2870 21247 2926 21256
rect 2884 20806 2912 21247
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2870 20088 2926 20097
rect 2870 20023 2926 20032
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 17678 2544 18090
rect 2686 17912 2742 17921
rect 2686 17847 2742 17856
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2320 17478 2372 17484
rect 2410 17504 2466 17513
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16794 1808 17138
rect 2332 17134 2360 17478
rect 2410 17439 2466 17448
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1688 16046 1716 16730
rect 2424 16658 2452 17439
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2424 16250 2452 16594
rect 2516 16590 2544 17614
rect 2700 16794 2728 17847
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2700 16130 2728 16730
rect 2608 16102 2728 16130
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 2608 15910 2636 16102
rect 2780 16040 2832 16046
rect 2700 15988 2780 15994
rect 2700 15982 2832 15988
rect 2700 15966 2820 15982
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1504 14618 1532 15506
rect 1688 15162 1716 15506
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1688 14618 1716 15098
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 14113 1532 14418
rect 1490 14104 1546 14113
rect 1688 14074 1716 14554
rect 1490 14039 1492 14048
rect 1544 14039 1546 14048
rect 1676 14068 1728 14074
rect 1492 14010 1544 14016
rect 1676 14010 1728 14016
rect 1504 13979 1532 14010
rect 1780 13954 1808 15846
rect 2700 15162 2728 15966
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2780 14816 2832 14822
rect 1950 14784 2006 14793
rect 2780 14758 2832 14764
rect 1950 14719 2006 14728
rect 1688 13926 1808 13954
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 10810 1532 11591
rect 1582 11112 1638 11121
rect 1582 11047 1584 11056
rect 1636 11047 1638 11056
rect 1584 11018 1636 11024
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1688 10554 1716 13926
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1504 10526 1716 10554
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1412 7449 1440 8502
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1504 7290 1532 10526
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8673 1624 8774
rect 1582 8664 1638 8673
rect 1582 8599 1638 8608
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1412 7262 1532 7290
rect 1412 5166 1440 7262
rect 1596 6905 1624 7686
rect 1688 7342 1716 7890
rect 1676 7336 1728 7342
rect 1674 7304 1676 7313
rect 1728 7304 1730 7313
rect 1674 7239 1730 7248
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6361 1624 6598
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1596 5370 1624 5607
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1400 5160 1452 5166
rect 1780 5137 1808 12582
rect 1872 12442 1900 13262
rect 1964 12782 1992 14719
rect 2792 12889 2820 14758
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1872 11762 1900 12378
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2042 11248 2098 11257
rect 2042 11183 2044 11192
rect 2096 11183 2098 11192
rect 2044 11154 2096 11160
rect 2056 10810 2084 11154
rect 2410 10840 2466 10849
rect 2044 10804 2096 10810
rect 2410 10775 2412 10784
rect 2044 10746 2096 10752
rect 2464 10775 2466 10784
rect 2412 10746 2464 10752
rect 2424 10606 2452 10746
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2700 10266 2728 11562
rect 2792 10577 2820 12815
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2884 10441 2912 20023
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2976 17338 3004 17818
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 3068 17082 3096 21791
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 3160 17241 3188 19343
rect 3146 17232 3202 17241
rect 3344 17218 3372 23559
rect 7470 23520 7526 24000
rect 22466 23520 22522 24000
rect 25594 23624 25650 23633
rect 25594 23559 25650 23568
rect 3422 23080 3478 23089
rect 3422 23015 3478 23024
rect 3436 22166 3464 23015
rect 3424 22160 3476 22166
rect 3424 22102 3476 22108
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 3882 20632 3938 20641
rect 5956 20624 6252 20644
rect 3882 20567 3938 20576
rect 3792 18352 3844 18358
rect 3514 18320 3570 18329
rect 3792 18294 3844 18300
rect 3514 18255 3570 18264
rect 3344 17190 3464 17218
rect 3146 17167 3202 17176
rect 3068 17054 3188 17082
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 14249 3096 15846
rect 3054 14240 3110 14249
rect 3054 14175 3110 14184
rect 3054 13968 3110 13977
rect 3054 13903 3110 13912
rect 2962 13424 3018 13433
rect 2962 13359 3018 13368
rect 2976 12889 3004 13359
rect 2962 12880 3018 12889
rect 2962 12815 3018 12824
rect 2870 10432 2926 10441
rect 2870 10367 2926 10376
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2228 10124 2280 10130
rect 2228 10066 2280 10072
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2042 9480 2098 9489
rect 2042 9415 2044 9424
rect 2096 9415 2098 9424
rect 2044 9386 2096 9392
rect 2148 9178 2176 9862
rect 2240 9722 2268 10066
rect 2792 9926 2820 10202
rect 2780 9920 2832 9926
rect 2686 9888 2742 9897
rect 2780 9862 2832 9868
rect 2686 9823 2742 9832
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2042 9072 2098 9081
rect 2042 9007 2098 9016
rect 2056 8634 2084 9007
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2056 8430 2084 8570
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2148 8090 2176 9114
rect 2240 8566 2268 9658
rect 2410 9616 2466 9625
rect 2410 9551 2466 9560
rect 2424 9110 2452 9551
rect 2700 9178 2728 9823
rect 2792 9586 2820 9862
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2424 8634 2452 9046
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2516 8498 2544 8978
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2686 8120 2742 8129
rect 2136 8084 2188 8090
rect 2686 8055 2688 8064
rect 2136 8026 2188 8032
rect 2740 8055 2742 8064
rect 2688 8026 2740 8032
rect 2148 7410 2176 8026
rect 2502 7984 2558 7993
rect 2502 7919 2504 7928
rect 2556 7919 2558 7928
rect 2504 7890 2556 7896
rect 2516 7546 2544 7890
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2516 7002 2544 7210
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 1858 6896 1914 6905
rect 1858 6831 1860 6840
rect 1912 6831 1914 6840
rect 1860 6802 1912 6808
rect 1872 6458 1900 6802
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5953 2452 6054
rect 2410 5944 2466 5953
rect 2410 5879 2466 5888
rect 2516 5794 2544 6938
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6118 2728 6598
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2688 6112 2740 6118
rect 2594 6080 2650 6089
rect 2688 6054 2740 6060
rect 2594 6015 2650 6024
rect 2608 5846 2636 6015
rect 2424 5778 2544 5794
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2412 5772 2544 5778
rect 2464 5766 2544 5772
rect 2412 5714 2464 5720
rect 1400 5102 1452 5108
rect 1766 5128 1822 5137
rect 1412 4826 1440 5102
rect 1766 5063 1822 5072
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 2424 4690 2452 5714
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5370 2544 5646
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2608 5302 2636 5782
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2700 4826 2728 6054
rect 2792 5914 2820 6190
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2884 5166 2912 5850
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 1582 4448 1638 4457
rect 1582 4383 1638 4392
rect 1400 4072 1452 4078
rect 1398 4040 1400 4049
rect 1452 4040 1454 4049
rect 1398 3975 1454 3984
rect 662 3768 718 3777
rect 1412 3738 1440 3975
rect 1596 3942 1624 4383
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 662 3703 718 3712
rect 1400 3732 1452 3738
rect 676 480 704 3703
rect 1400 3674 1452 3680
rect 2608 3398 2636 4626
rect 2884 4282 2912 4762
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2686 3904 2742 3913
rect 2686 3839 2742 3848
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 1465 1624 2246
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 2056 480 2084 2790
rect 2700 2650 2728 3839
rect 2976 3738 3004 12815
rect 3068 6089 3096 13903
rect 3160 13138 3188 17054
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3252 14618 3280 14962
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3252 13802 3280 14418
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3252 13326 3280 13738
rect 3240 13320 3292 13326
rect 3238 13288 3240 13297
rect 3292 13288 3294 13297
rect 3238 13223 3294 13232
rect 3160 13110 3280 13138
rect 3252 10169 3280 13110
rect 3436 11665 3464 17190
rect 3528 13977 3556 18255
rect 3804 17338 3832 18294
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3790 17096 3846 17105
rect 3790 17031 3846 17040
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16522 3740 16934
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3620 16046 3648 16390
rect 3712 16114 3740 16458
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3712 15434 3740 16050
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 14550 3740 14758
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3606 14240 3662 14249
rect 3606 14175 3662 14184
rect 3514 13968 3570 13977
rect 3514 13903 3570 13912
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3238 10160 3294 10169
rect 3238 10095 3294 10104
rect 3436 9722 3464 10746
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3528 9518 3556 9862
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3620 9450 3648 14175
rect 3804 13569 3832 17031
rect 3896 15745 3924 20567
rect 7484 20369 7512 23520
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 7470 20360 7526 20369
rect 7470 20295 7526 20304
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 4160 18828 4212 18834
rect 3988 16017 4016 18799
rect 4160 18770 4212 18776
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4080 18426 4108 18702
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4172 18358 4200 18770
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 5460 17814 5488 18566
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 4066 17640 4122 17649
rect 4066 17575 4122 17584
rect 4080 16130 4108 17575
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4448 17202 4476 17478
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4172 16522 4200 17138
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4172 16250 4200 16458
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4080 16102 4200 16130
rect 3974 16008 4030 16017
rect 3974 15943 4030 15952
rect 3882 15736 3938 15745
rect 3882 15671 3938 15680
rect 4172 15638 4200 16102
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3882 15328 3938 15337
rect 3882 15263 3938 15272
rect 3790 13560 3846 13569
rect 3790 13495 3846 13504
rect 3790 12608 3846 12617
rect 3790 12543 3846 12552
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8566 3464 8910
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3514 7848 3570 7857
rect 3514 7783 3570 7792
rect 3146 7032 3202 7041
rect 3146 6967 3202 6976
rect 3054 6080 3110 6089
rect 3054 6015 3110 6024
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3068 3738 3096 4558
rect 3160 4146 3188 6967
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2976 3618 3004 3674
rect 2792 3590 3004 3618
rect 2792 3194 2820 3590
rect 3252 3534 3280 4082
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 3074 2912 3470
rect 3252 3210 3280 3470
rect 3252 3194 3372 3210
rect 3252 3188 3384 3194
rect 3252 3182 3332 3188
rect 3332 3130 3384 3136
rect 2792 3046 2912 3074
rect 2792 2650 2820 3046
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2976 2582 3004 2926
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2516 2417 2544 2450
rect 2502 2408 2558 2417
rect 2502 2343 2558 2352
rect 3528 480 3556 7783
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6322 3648 7142
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3804 5914 3832 12543
rect 3896 6361 3924 15263
rect 4068 14952 4120 14958
rect 4120 14900 4292 14906
rect 4068 14894 4292 14900
rect 4080 14878 4292 14894
rect 4066 14648 4122 14657
rect 4066 14583 4122 14592
rect 4080 13433 4108 14583
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 4264 11694 4292 14878
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3988 10674 4016 11562
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11144 4212 11150
rect 4066 11112 4122 11121
rect 4160 11086 4212 11092
rect 4066 11047 4068 11056
rect 4120 11047 4122 11056
rect 4068 11018 4120 11024
rect 4068 10804 4120 10810
rect 4172 10792 4200 11086
rect 4120 10764 4200 10792
rect 4068 10746 4120 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4080 9586 4108 10066
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9178 4108 9318
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4264 8265 4292 11494
rect 4250 8256 4306 8265
rect 4250 8191 4306 8200
rect 4264 7993 4292 8191
rect 4250 7984 4306 7993
rect 4250 7919 4306 7928
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4264 6905 4292 7482
rect 4250 6896 4306 6905
rect 4250 6831 4306 6840
rect 3882 6352 3938 6361
rect 3882 6287 3938 6296
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3608 5024 3660 5030
rect 3606 4992 3608 5001
rect 3660 4992 3662 5001
rect 3606 4927 3662 4936
rect 3712 4282 3740 5170
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3606 3904 3662 3913
rect 3606 3839 3662 3848
rect 3620 3602 3648 3839
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3712 2582 3740 4014
rect 3804 3534 3832 5850
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 3618 4016 4966
rect 3896 3590 4016 3618
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3804 3058 3832 3470
rect 3896 3369 3924 3590
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3882 3360 3938 3369
rect 3882 3295 3938 3304
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 662 0 718 480
rect 2042 0 2098 480
rect 3514 0 3570 480
rect 3988 377 4016 3402
rect 4080 2514 4108 6054
rect 4264 5953 4292 6054
rect 4250 5944 4306 5953
rect 4250 5879 4252 5888
rect 4304 5879 4306 5888
rect 4252 5850 4304 5856
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4172 2394 4200 4422
rect 4264 4078 4292 4762
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4356 3505 4384 16934
rect 4448 16794 4476 17138
rect 4724 17066 4752 17478
rect 5460 17338 5488 17750
rect 5644 17746 5672 18362
rect 7392 18154 7420 18566
rect 8496 18426 8524 19178
rect 8588 18834 8616 19246
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10336 18834 10364 19110
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5644 17202 5672 17682
rect 7392 17542 7420 18090
rect 7470 17776 7526 17785
rect 7470 17711 7526 17720
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4540 16182 4568 16526
rect 4710 16416 4766 16425
rect 4710 16351 4766 16360
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4436 15632 4488 15638
rect 4434 15600 4436 15609
rect 4488 15600 4490 15609
rect 4434 15535 4490 15544
rect 4448 15162 4476 15535
rect 4540 15502 4568 15533
rect 4528 15496 4580 15502
rect 4526 15464 4528 15473
rect 4580 15464 4582 15473
rect 4526 15399 4582 15408
rect 4540 15162 4568 15399
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4434 14104 4490 14113
rect 4434 14039 4436 14048
rect 4488 14039 4490 14048
rect 4436 14010 4488 14016
rect 4540 12186 4568 15098
rect 4724 14906 4752 16351
rect 4908 15910 4936 16594
rect 7392 16590 7420 17478
rect 7484 17377 7512 17711
rect 7470 17368 7526 17377
rect 7470 17303 7526 17312
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 8298 16552 8354 16561
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6656 16250 6684 16526
rect 7300 16250 7328 16526
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4908 15706 4936 15846
rect 5722 15736 5778 15745
rect 4896 15700 4948 15706
rect 5722 15671 5778 15680
rect 6182 15736 6238 15745
rect 6182 15671 6184 15680
rect 4896 15642 4948 15648
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4816 15162 4844 15438
rect 5736 15162 5764 15671
rect 6236 15671 6238 15680
rect 6184 15642 6236 15648
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 4802 14920 4858 14929
rect 4724 14878 4802 14906
rect 4802 14855 4858 14864
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12782 4752 13126
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4816 12458 4844 14855
rect 5828 14618 5856 15302
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 6288 14822 6316 15438
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 14816 6328 14822
rect 6274 14784 6276 14793
rect 6328 14784 6330 14793
rect 6274 14719 6330 14728
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13462 5580 14214
rect 5644 13530 5672 14486
rect 5722 14104 5778 14113
rect 5828 14074 5856 14554
rect 6288 14521 6316 14719
rect 6274 14512 6330 14521
rect 6274 14447 6330 14456
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5722 14039 5778 14048
rect 5816 14068 5868 14074
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5736 13326 5764 14039
rect 5816 14010 5868 14016
rect 6288 14006 6316 14282
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5736 12986 5764 13262
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 4896 12640 4948 12646
rect 4948 12600 5028 12628
rect 4896 12582 4948 12588
rect 4816 12430 4936 12458
rect 4540 12158 4752 12186
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4448 10742 4476 11154
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4434 10568 4490 10577
rect 4434 10503 4490 10512
rect 4448 9178 4476 10503
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4448 8566 4476 9114
rect 4540 9024 4568 11630
rect 4632 11393 4660 12038
rect 4618 11384 4674 11393
rect 4618 11319 4674 11328
rect 4724 9722 4752 12158
rect 4908 10554 4936 12430
rect 5000 12306 5028 12600
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11898 5120 12174
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5184 11762 5212 12786
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5264 12232 5316 12238
rect 5262 12200 5264 12209
rect 5316 12200 5318 12209
rect 5262 12135 5318 12144
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5080 11688 5132 11694
rect 5078 11656 5080 11665
rect 5132 11656 5134 11665
rect 5078 11591 5134 11600
rect 5184 11354 5212 11698
rect 5276 11626 5304 12135
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5184 10674 5212 11290
rect 5276 11150 5304 11562
rect 5368 11529 5396 12650
rect 5552 12442 5580 12718
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5368 10849 5396 11455
rect 5460 11354 5488 12242
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5354 10840 5410 10849
rect 5354 10775 5410 10784
rect 5446 10704 5502 10713
rect 5172 10668 5224 10674
rect 5446 10639 5502 10648
rect 5172 10610 5224 10616
rect 4908 10526 5028 10554
rect 4804 10464 4856 10470
rect 4802 10432 4804 10441
rect 4896 10464 4948 10470
rect 4856 10432 4858 10441
rect 4896 10406 4948 10412
rect 4802 10367 4858 10376
rect 4908 10266 4936 10406
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5000 10198 5028 10526
rect 4988 10192 5040 10198
rect 4894 10160 4950 10169
rect 4988 10134 5040 10140
rect 4894 10095 4950 10104
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4804 9648 4856 9654
rect 4632 9596 4804 9602
rect 4632 9590 4856 9596
rect 4632 9574 4844 9590
rect 4632 9518 4660 9574
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4620 9036 4672 9042
rect 4540 8996 4620 9024
rect 4620 8978 4672 8984
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4540 7342 4568 8230
rect 4632 7818 4660 8978
rect 4908 8022 4936 10095
rect 5000 9178 5028 10134
rect 5184 10130 5212 10610
rect 5460 10266 5488 10639
rect 5448 10260 5500 10266
rect 5500 10220 5580 10248
rect 5448 10202 5500 10208
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5460 9586 5488 9998
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4986 8528 5042 8537
rect 4986 8463 4988 8472
rect 5040 8463 5042 8472
rect 5080 8492 5132 8498
rect 4988 8434 5040 8440
rect 5080 8434 5132 8440
rect 4986 8120 5042 8129
rect 4986 8055 4988 8064
rect 5040 8055 5042 8064
rect 4988 8026 5040 8032
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4632 4690 4660 7754
rect 4908 7478 4936 7958
rect 5000 7546 5028 8026
rect 5092 7886 5120 8434
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6254 4752 7142
rect 5092 7002 5120 7822
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7410 5212 7686
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5092 6662 5120 6938
rect 5276 6882 5304 7346
rect 5184 6866 5304 6882
rect 5172 6860 5304 6866
rect 5224 6854 5304 6860
rect 5172 6802 5224 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5184 6390 5212 6802
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5914 4752 6190
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4710 5672 4766 5681
rect 4710 5607 4766 5616
rect 4724 5370 4752 5607
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4724 5166 4752 5306
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4632 4185 4660 4626
rect 4802 4584 4858 4593
rect 4802 4519 4858 4528
rect 4618 4176 4674 4185
rect 4618 4111 4674 4120
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4540 3738 4568 4014
rect 4632 4010 4660 4111
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4342 3496 4398 3505
rect 4342 3431 4398 3440
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 2689 4292 3334
rect 4816 3194 4844 4519
rect 5276 4282 5304 6598
rect 5368 4593 5396 9386
rect 5460 8974 5488 9522
rect 5552 9178 5580 10220
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5540 9172 5592 9178
rect 5592 9132 5672 9160
rect 5540 9114 5592 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5354 4584 5410 4593
rect 5354 4519 5410 4528
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5460 4162 5488 8502
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6458 5580 6802
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5552 5778 5580 6394
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 5302 5580 5714
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 4826 5580 5238
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5460 4146 5580 4162
rect 5460 4140 5592 4146
rect 5460 4134 5540 4140
rect 5540 4082 5592 4088
rect 5644 4049 5672 9132
rect 5736 8401 5764 9318
rect 5722 8392 5778 8401
rect 5722 8327 5778 8336
rect 5630 4040 5686 4049
rect 5630 3975 5686 3984
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3777 5212 3878
rect 5170 3768 5226 3777
rect 5170 3703 5226 3712
rect 5184 3602 5212 3703
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3194 5212 3538
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4816 2990 4844 3130
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4250 2680 4306 2689
rect 4250 2615 4306 2624
rect 4080 2366 4200 2394
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4080 921 4108 2366
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 4908 480 4936 2382
rect 5092 2145 5120 2790
rect 5828 2553 5856 13126
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6288 12986 6316 13466
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5920 9178 5948 9522
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6104 8090 6132 8298
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6380 7993 6408 15098
rect 6472 14890 6500 15438
rect 6656 15337 6684 16186
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6826 15056 6882 15065
rect 6826 14991 6828 15000
rect 6880 14991 6882 15000
rect 6828 14962 6880 14968
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6932 14113 6960 16186
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15706 7328 15846
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7392 15638 7420 16526
rect 8298 16487 8354 16496
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16114 7788 16390
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7576 15366 7604 15846
rect 7944 15638 7972 16050
rect 8312 15881 8340 16487
rect 8496 16114 8524 18362
rect 9126 16552 9182 16561
rect 9126 16487 9182 16496
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8956 16046 8984 16390
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8298 15872 8354 15881
rect 8298 15807 8354 15816
rect 8772 15706 8800 15914
rect 8956 15706 8984 15982
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7116 14482 7144 14826
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 6918 14104 6974 14113
rect 7116 14074 7144 14418
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 6918 14039 6974 14048
rect 7104 14068 7156 14074
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6840 13530 6868 13942
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6564 12986 6592 13398
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6932 12345 6960 14039
rect 7104 14010 7156 14016
rect 7208 13870 7236 14350
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6918 12336 6974 12345
rect 7208 12322 7236 13806
rect 7484 13734 7512 14418
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 13530 7512 13670
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7378 13288 7434 13297
rect 7378 13223 7434 13232
rect 7392 13190 7420 13223
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12442 7420 13126
rect 7576 13025 7604 15302
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 13938 7972 14214
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8036 13530 8064 13738
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8128 13394 8156 14418
rect 8220 14346 8248 14758
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8220 13938 8248 14282
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8220 13462 8248 13874
rect 9048 13870 9076 14350
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8390 13560 8446 13569
rect 8312 13504 8390 13512
rect 8312 13484 8392 13504
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7562 13016 7618 13025
rect 8128 12986 8156 13330
rect 8312 13297 8340 13484
rect 8444 13495 8446 13504
rect 8392 13466 8444 13472
rect 8772 13462 8800 13493
rect 8760 13456 8812 13462
rect 8758 13424 8760 13433
rect 8812 13424 8814 13433
rect 8758 13359 8814 13368
rect 8852 13388 8904 13394
rect 8298 13288 8354 13297
rect 8208 13252 8260 13258
rect 8298 13223 8354 13232
rect 8208 13194 8260 13200
rect 7562 12951 7618 12960
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8220 12442 8248 13194
rect 8312 12850 8340 13223
rect 8772 12986 8800 13359
rect 8852 13330 8904 13336
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 6918 12271 6974 12280
rect 7116 12294 7236 12322
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9178 6960 9862
rect 7116 9625 7144 12294
rect 7194 12200 7250 12209
rect 7194 12135 7250 12144
rect 7208 11626 7236 12135
rect 7392 11694 7420 12378
rect 8496 12102 8524 12718
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11801 8524 12038
rect 8482 11792 8538 11801
rect 8482 11727 8538 11736
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7930 11520 7986 11529
rect 7654 11384 7710 11393
rect 7654 11319 7656 11328
rect 7708 11319 7710 11328
rect 7656 11290 7708 11296
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7102 9616 7158 9625
rect 7102 9551 7158 9560
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 8634 6684 8978
rect 6932 8974 6960 9114
rect 6920 8968 6972 8974
rect 6972 8928 7052 8956
rect 6920 8910 6972 8916
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6366 7984 6422 7993
rect 6366 7919 6422 7928
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6322 6316 6598
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5846 6316 6258
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 6288 5370 6316 5782
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 6748 3602 6776 5238
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6840 2650 6868 4422
rect 6932 2990 6960 8502
rect 7024 7818 7052 8928
rect 7286 8800 7342 8809
rect 7286 8735 7342 8744
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7116 8090 7144 8298
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7300 7954 7328 8735
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 7024 6934 7052 7754
rect 7300 7546 7328 7890
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 4826 7420 5510
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7286 4176 7342 4185
rect 7392 4146 7420 4762
rect 7286 4111 7342 4120
rect 7380 4140 7432 4146
rect 7300 4078 7328 4111
rect 7380 4082 7432 4088
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7024 2650 7052 3538
rect 7208 3126 7236 3878
rect 7300 3738 7328 4014
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7392 3670 7420 4082
rect 7484 4010 7512 5743
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7392 3194 7420 3606
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5814 2544 5870 2553
rect 7576 2514 7604 11018
rect 7668 10674 7696 11290
rect 7852 11150 7880 11494
rect 7930 11455 7986 11464
rect 7748 11144 7800 11150
rect 7746 11112 7748 11121
rect 7840 11144 7892 11150
rect 7800 11112 7802 11121
rect 7944 11121 7972 11455
rect 7840 11086 7892 11092
rect 7930 11112 7986 11121
rect 7746 11047 7802 11056
rect 7760 10742 7788 11047
rect 7852 10810 7880 11086
rect 7930 11047 7986 11056
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8772 10554 8800 12922
rect 8864 12646 8892 13330
rect 9048 13326 9076 13806
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9048 12918 9076 13262
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 8852 12640 8904 12646
rect 8850 12608 8852 12617
rect 8904 12608 8906 12617
rect 8850 12543 8906 12552
rect 8312 10526 8800 10554
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8090 7880 8230
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 8128 7886 8156 8978
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5953 7788 6054
rect 7746 5944 7802 5953
rect 7746 5879 7802 5888
rect 8312 5001 8340 10526
rect 8666 10432 8722 10441
rect 8666 10367 8722 10376
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8838 8432 9318
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8498 8432 8774
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8496 7546 8524 8026
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8680 6254 8708 10367
rect 9140 8634 9168 16487
rect 9232 15065 9260 18770
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9600 17626 9628 18362
rect 10336 18086 10364 18770
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 9600 17610 9720 17626
rect 9600 17604 9732 17610
rect 9600 17598 9680 17604
rect 9680 17546 9732 17552
rect 9784 17542 9812 18022
rect 10428 17746 10456 22102
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 13648 20058 13676 20334
rect 14096 20324 14148 20330
rect 14096 20266 14148 20272
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13648 19378 13676 19994
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 14108 18970 14136 20266
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14844 19174 14872 20198
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 17972 19310 18000 19790
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10704 18737 10732 18838
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12716 18760 12768 18766
rect 10690 18728 10746 18737
rect 12714 18728 12716 18737
rect 12768 18728 12770 18737
rect 10690 18663 10746 18672
rect 12636 18686 12714 18714
rect 10704 18426 10732 18663
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9784 17270 9812 17478
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 16250 9720 16594
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16114 9812 17206
rect 9968 17134 9996 17614
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10152 17202 10180 17478
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 9956 17128 10008 17134
rect 9954 17096 9956 17105
rect 10008 17096 10010 17105
rect 9954 17031 10010 17040
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9218 15056 9274 15065
rect 9218 14991 9274 15000
rect 9232 14618 9260 14991
rect 9784 14822 9812 15506
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9784 13977 9812 14758
rect 9770 13968 9826 13977
rect 9220 13932 9272 13938
rect 9770 13903 9826 13912
rect 9220 13874 9272 13880
rect 9232 13530 9260 13874
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9784 12986 9812 13738
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9862 12880 9918 12889
rect 9862 12815 9864 12824
rect 9916 12815 9918 12824
rect 9864 12786 9916 12792
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 8838 9720 12038
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9140 8430 9168 8570
rect 9416 8430 9444 8774
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9128 8424 9180 8430
rect 9034 8392 9090 8401
rect 9128 8366 9180 8372
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9034 8327 9090 8336
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 8022 8984 8230
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8956 7546 8984 7958
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5234 8800 6054
rect 8864 5681 8892 6122
rect 8850 5672 8906 5681
rect 8850 5607 8852 5616
rect 8904 5607 8906 5616
rect 8852 5578 8904 5584
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8576 5024 8628 5030
rect 8298 4992 8354 5001
rect 8576 4966 8628 4972
rect 8298 4927 8354 4936
rect 8312 3641 8340 4927
rect 8588 4826 8616 4966
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8574 4720 8630 4729
rect 8574 4655 8630 4664
rect 8588 4622 8616 4655
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8496 4282 8524 4558
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8588 4214 8616 4558
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 8772 3194 8800 4014
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9048 2990 9076 8327
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6322 9352 6598
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9128 6248 9180 6254
rect 9126 6216 9128 6225
rect 9180 6216 9182 6225
rect 9126 6151 9182 6160
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 4146 9260 5170
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9140 3738 9168 3946
rect 9416 3913 9444 8366
rect 9508 7886 9536 8502
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9600 7886 9628 8434
rect 9876 8090 9904 12786
rect 9968 8129 9996 17031
rect 10244 16794 10272 17546
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10244 16114 10272 16730
rect 10428 16250 10456 17002
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16794 10824 16934
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10244 15502 10272 16050
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10152 14822 10180 15438
rect 10244 15162 10272 15438
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10046 13424 10102 13433
rect 10046 13359 10048 13368
rect 10100 13359 10102 13368
rect 10048 13330 10100 13336
rect 10152 12753 10180 14758
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10244 13870 10272 14486
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13326 10272 13670
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10138 12744 10194 12753
rect 10138 12679 10140 12688
rect 10192 12679 10194 12688
rect 10140 12650 10192 12656
rect 10152 12102 10180 12650
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10336 11257 10364 15846
rect 10414 15328 10470 15337
rect 10414 15263 10470 15272
rect 10428 13802 10456 15263
rect 10506 14104 10562 14113
rect 10562 14048 10640 14056
rect 10506 14039 10508 14048
rect 10560 14028 10640 14048
rect 10508 14010 10560 14016
rect 10612 13870 10640 14028
rect 10508 13864 10560 13870
rect 10600 13864 10652 13870
rect 10508 13806 10560 13812
rect 10598 13832 10600 13841
rect 10652 13832 10654 13841
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10428 13530 10456 13738
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10322 11248 10378 11257
rect 10322 11183 10378 11192
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9722 10272 10066
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10428 9602 10456 13466
rect 10520 11694 10548 13806
rect 10598 13767 10654 13776
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10336 9574 10456 9602
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 9954 8120 10010 8129
rect 9864 8084 9916 8090
rect 9954 8055 10010 8064
rect 9864 8026 9916 8032
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7546 9628 7822
rect 9876 7546 9904 8026
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 10152 6769 10180 8191
rect 10336 7274 10364 9574
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 8838 10456 9454
rect 10416 8832 10468 8838
rect 10414 8800 10416 8809
rect 10468 8800 10470 8809
rect 10414 8735 10470 8744
rect 10612 8072 10640 13767
rect 10520 8044 10640 8072
rect 10520 7546 10548 8044
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10520 7342 10548 7482
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10336 6866 10364 7210
rect 10520 7041 10548 7278
rect 10612 7206 10640 7890
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10506 7032 10562 7041
rect 10612 7002 10640 7142
rect 10506 6967 10562 6976
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10138 6760 10194 6769
rect 10138 6695 10194 6704
rect 10152 6458 10180 6695
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 5250 9720 6326
rect 10152 6186 10180 6394
rect 10336 6338 10364 6802
rect 10244 6310 10364 6338
rect 10414 6352 10470 6361
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9600 5222 9720 5250
rect 9600 5166 9628 5222
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 4049 9628 4082
rect 9586 4040 9642 4049
rect 9586 3975 9642 3984
rect 9402 3904 9458 3913
rect 9402 3839 9458 3848
rect 9692 3754 9720 4150
rect 10244 3777 10272 6310
rect 10414 6287 10470 6296
rect 10508 6316 10560 6322
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10336 5953 10364 6190
rect 10322 5944 10378 5953
rect 10322 5879 10324 5888
rect 10376 5879 10378 5888
rect 10324 5850 10376 5856
rect 10322 4584 10378 4593
rect 10322 4519 10378 4528
rect 10336 4078 10364 4519
rect 10428 4146 10456 6287
rect 10508 6258 10560 6264
rect 10520 4826 10548 6258
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10520 4214 10548 4762
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9600 3726 9720 3754
rect 10230 3768 10286 3777
rect 9600 3466 9628 3726
rect 10336 3738 10364 4014
rect 10230 3703 10286 3712
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10138 3496 10194 3505
rect 9588 3460 9640 3466
rect 10138 3431 10194 3440
rect 9588 3402 9640 3408
rect 9600 3058 9628 3402
rect 10152 3194 10180 3431
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 5814 2479 5870 2488
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5078 2136 5134 2145
rect 5956 2128 6252 2148
rect 5078 2071 5134 2080
rect 6380 480 6408 2382
rect 7760 480 7788 2858
rect 9600 2650 9628 2994
rect 10152 2990 10180 3130
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9770 2544 9826 2553
rect 10704 2514 10732 16730
rect 10888 16674 10916 18566
rect 12636 18358 12664 18686
rect 12714 18663 12770 18672
rect 12716 18624 12768 18630
rect 12820 18612 12848 18770
rect 12768 18584 12848 18612
rect 12716 18566 12768 18572
rect 12820 18426 12848 18584
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 13820 18080 13872 18086
rect 13740 18028 13820 18034
rect 13740 18022 13872 18028
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13740 18006 13860 18022
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 13740 17882 13768 18006
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11072 17134 11100 17682
rect 13464 17338 13492 17750
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10796 16646 10916 16674
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10796 16522 10824 16646
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 15706 10824 16458
rect 10888 15706 10916 16526
rect 10980 15978 11008 16662
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 16250 11100 16594
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10888 13938 10916 14486
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11716 14074 11744 14418
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11900 14006 11928 14214
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10888 13190 10916 13874
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11716 13569 11744 13738
rect 11702 13560 11758 13569
rect 12452 13530 12480 14010
rect 11702 13495 11758 13504
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12850 10916 13126
rect 13004 12866 13032 17070
rect 13464 16114 13492 17274
rect 13648 16794 13676 17478
rect 13924 17377 13952 18022
rect 14016 17746 14044 18294
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13910 17368 13966 17377
rect 14016 17338 14044 17682
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14186 17640 14242 17649
rect 13910 17303 13966 17312
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14108 17270 14136 17614
rect 14186 17575 14242 17584
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 14200 16998 14228 17575
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13556 16250 13584 16458
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13082 15600 13138 15609
rect 13082 15535 13138 15544
rect 13096 15337 13124 15535
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13082 15328 13138 15337
rect 13082 15263 13138 15272
rect 13096 15162 13124 15263
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13188 14618 13216 14826
rect 13280 14822 13308 15438
rect 13464 15162 13492 15914
rect 13556 15706 13584 16186
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13556 15026 13584 15302
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13082 12880 13138 12889
rect 10876 12844 10928 12850
rect 13004 12838 13082 12866
rect 13082 12815 13138 12824
rect 10876 12786 10928 12792
rect 10888 12646 10916 12786
rect 13096 12782 13124 12815
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13174 12744 13230 12753
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10888 12102 10916 12582
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11898 11192 12038
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10782 11792 10838 11801
rect 10782 11727 10838 11736
rect 10796 9178 10824 11727
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11348 11257 11376 11494
rect 11334 11248 11390 11257
rect 11334 11183 11390 11192
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9586 10916 10066
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8498 11192 8774
rect 11624 8498 11652 9862
rect 12084 9081 12112 12718
rect 12912 12646 12940 12718
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12728 11898 12756 12582
rect 13096 12442 13124 12718
rect 13174 12679 13230 12688
rect 13188 12481 13216 12679
rect 13174 12472 13230 12481
rect 13084 12436 13136 12442
rect 13174 12407 13230 12416
rect 13084 12378 13136 12384
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12990 11792 13046 11801
rect 12990 11727 12992 11736
rect 13044 11727 13046 11736
rect 12992 11698 13044 11704
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12360 11354 12388 11562
rect 13004 11558 13032 11698
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 10198 13032 10542
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12164 9648 12216 9654
rect 12162 9616 12164 9625
rect 12216 9616 12218 9625
rect 12452 9586 12480 9862
rect 12162 9551 12218 9560
rect 12440 9580 12492 9586
rect 12176 9450 12204 9551
rect 12440 9522 12492 9528
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12070 9072 12126 9081
rect 11796 9036 11848 9042
rect 12070 9007 12126 9016
rect 11796 8978 11848 8984
rect 11808 8634 11836 8978
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11152 8492 11204 8498
rect 11072 8452 11152 8480
rect 11072 8378 11100 8452
rect 11152 8434 11204 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 10888 8350 11100 8378
rect 10888 8090 10916 8350
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11808 7993 11836 8570
rect 11992 8362 12020 8910
rect 12268 8430 12296 9318
rect 12452 8974 12480 9522
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 9178 12572 9318
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11992 8129 12020 8298
rect 11978 8120 12034 8129
rect 12452 8090 12480 8910
rect 12544 8498 12572 9114
rect 12912 8945 12940 9386
rect 12898 8936 12954 8945
rect 12898 8871 12954 8880
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 13280 8401 13308 14758
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13450 13696 13506 13705
rect 13450 13631 13506 13640
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12850 13400 13330
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13372 12481 13400 12786
rect 13464 12782 13492 13631
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13358 12472 13414 12481
rect 13358 12407 13360 12416
rect 13412 12407 13414 12416
rect 13360 12378 13412 12384
rect 13372 11762 13400 12378
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13372 11354 13400 11698
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13358 11112 13414 11121
rect 13464 11098 13492 12242
rect 13648 11642 13676 16390
rect 13740 16130 13768 16594
rect 14372 16584 14424 16590
rect 14370 16552 14372 16561
rect 14424 16552 14426 16561
rect 14370 16487 14426 16496
rect 14384 16182 14412 16487
rect 14372 16176 14424 16182
rect 13740 16102 13860 16130
rect 14372 16118 14424 16124
rect 13832 16046 13860 16102
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 14002 15600 14058 15609
rect 14002 15535 14004 15544
rect 14056 15535 14058 15544
rect 14004 15506 14056 15512
rect 14476 15502 14504 18906
rect 14844 18290 14872 19110
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14738 18184 14794 18193
rect 14738 18119 14740 18128
rect 14792 18119 14794 18128
rect 14740 18090 14792 18096
rect 14844 17626 14872 18226
rect 15856 17746 15884 19246
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16500 17814 16528 19110
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 14752 17598 14872 17626
rect 14752 17542 14780 17598
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17202 14780 17478
rect 15856 17202 15884 17682
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 16500 17338 16528 17750
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16578 17232 16634 17241
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 15844 17196 15896 17202
rect 16578 17167 16634 17176
rect 16672 17196 16724 17202
rect 15844 17138 15896 17144
rect 14648 16992 14700 16998
rect 14646 16960 14648 16969
rect 14700 16960 14702 16969
rect 14646 16895 14702 16904
rect 14752 16454 14780 17138
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 15910 14780 16390
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13740 14890 13768 15302
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14108 13870 14136 14486
rect 14476 14482 14504 15438
rect 14752 15094 14780 15846
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 13938 14228 14214
rect 14476 14074 14504 14418
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12646 13952 13126
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 11762 13952 12582
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13414 11070 13492 11098
rect 13556 11614 13676 11642
rect 13358 11047 13360 11056
rect 13412 11047 13414 11056
rect 13360 11018 13412 11024
rect 13266 8392 13322 8401
rect 13266 8327 13322 8336
rect 11978 8055 12034 8064
rect 12440 8084 12492 8090
rect 11794 7984 11850 7993
rect 11794 7919 11850 7928
rect 11888 7948 11940 7954
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 11808 7041 11836 7919
rect 11888 7890 11940 7896
rect 11794 7032 11850 7041
rect 11794 6967 11850 6976
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 11900 5846 11928 7890
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11520 5772 11572 5778
rect 11440 5732 11520 5760
rect 11440 5030 11468 5732
rect 11520 5714 11572 5720
rect 11900 5370 11928 5782
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 11440 4826 11468 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11440 4729 11468 4762
rect 11900 4758 11928 5306
rect 11612 4752 11664 4758
rect 11426 4720 11482 4729
rect 11612 4694 11664 4700
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11426 4655 11482 4664
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 11348 3602 11376 4082
rect 11624 4049 11652 4694
rect 11900 4282 11928 4694
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11610 4040 11666 4049
rect 11610 3975 11666 3984
rect 11624 3942 11652 3975
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3738 11652 3878
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11900 3670 11928 4218
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11348 3194 11376 3538
rect 11532 3194 11560 3606
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 9770 2479 9772 2488
rect 9824 2479 9826 2488
rect 10692 2508 10744 2514
rect 9772 2450 9824 2456
rect 10692 2450 10744 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 10600 2440 10652 2446
rect 11992 2417 12020 8055
rect 12440 8026 12492 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7410 12388 7890
rect 12636 7546 12664 7958
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 5914 12480 7346
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 13556 2990 13584 11614
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11354 13676 11494
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13924 11234 13952 11698
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13648 11206 13952 11234
rect 13648 10606 13676 11206
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 8838 13676 9862
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 8022 13676 8774
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13648 6118 13676 6802
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5817 13676 6054
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 10600 2382 10652 2388
rect 11978 2408 12034 2417
rect 9232 480 9260 2382
rect 10612 480 10640 2382
rect 11978 2343 12034 2352
rect 12084 480 12112 2858
rect 13740 2530 13768 11018
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13924 9722 13952 10134
rect 14016 10130 14044 11290
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 8838 14044 9454
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14108 8650 14136 13806
rect 14200 9353 14228 13874
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 11354 14412 12582
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10810 14320 11086
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14292 10198 14320 10746
rect 14384 10266 14412 11290
rect 14568 10713 14596 14894
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14752 12918 14780 13126
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14752 12782 14780 12854
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14646 12200 14702 12209
rect 14646 12135 14702 12144
rect 14660 12102 14688 12135
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11937 14688 12038
rect 14646 11928 14702 11937
rect 14646 11863 14702 11872
rect 14844 10713 14872 16934
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15198 16008 15254 16017
rect 15198 15943 15254 15952
rect 15474 16008 15530 16017
rect 15474 15943 15530 15952
rect 15212 15910 15240 15943
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15212 15178 15240 15642
rect 15120 15162 15240 15178
rect 15108 15156 15240 15162
rect 15160 15150 15240 15156
rect 15108 15098 15160 15104
rect 15488 14958 15516 15943
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15672 15178 15700 15846
rect 15764 15706 15792 15846
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 15672 15150 15792 15178
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14952 15528 14958
rect 14922 14920 14978 14929
rect 15476 14894 15528 14900
rect 14922 14855 14924 14864
rect 14976 14855 14978 14864
rect 15384 14884 15436 14890
rect 14924 14826 14976 14832
rect 15384 14826 15436 14832
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15120 12866 15148 12922
rect 15212 12866 15240 13942
rect 15120 12838 15240 12866
rect 15120 12782 15148 12838
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 14554 10704 14610 10713
rect 14554 10639 14610 10648
rect 14830 10704 14886 10713
rect 14830 10639 14886 10648
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14186 9344 14242 9353
rect 14186 9279 14242 9288
rect 14016 8622 14136 8650
rect 14016 8265 14044 8622
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 14016 6866 14044 8191
rect 14200 6866 14228 9279
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14752 7410 14780 8026
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14844 7313 14872 10639
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15028 8090 15056 9386
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14830 7304 14886 7313
rect 14280 7268 14332 7274
rect 15120 7274 15148 9318
rect 14830 7239 14886 7248
rect 15108 7268 15160 7274
rect 14280 7210 14332 7216
rect 15108 7210 15160 7216
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14016 6118 14044 6802
rect 14292 6798 14320 7210
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 14292 6458 14320 6734
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 4185 14044 6054
rect 14568 5574 14596 6122
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4690 14228 5102
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14568 4593 14596 5510
rect 14660 4826 14688 6054
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5098 14964 5510
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14554 4584 14610 4593
rect 14554 4519 14610 4528
rect 14002 4176 14058 4185
rect 14002 4111 14058 4120
rect 14660 4078 14688 4762
rect 15028 4078 15056 6598
rect 15106 6352 15162 6361
rect 15304 6322 15332 6734
rect 15106 6287 15108 6296
rect 15160 6287 15162 6296
rect 15292 6316 15344 6322
rect 15108 6258 15160 6264
rect 15292 6258 15344 6264
rect 15304 5574 15332 6258
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15120 4146 15148 5306
rect 15396 5137 15424 14826
rect 15672 14482 15700 14962
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14074 15608 14282
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15580 9382 15608 9998
rect 15764 9625 15792 15150
rect 16394 14512 16450 14521
rect 16394 14447 16396 14456
rect 16448 14447 16450 14456
rect 16396 14418 16448 14424
rect 15844 14408 15896 14414
rect 16408 14362 16436 14418
rect 15844 14350 15896 14356
rect 15856 13938 15884 14350
rect 16316 14334 16436 14362
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16210 13968 16266 13977
rect 15844 13932 15896 13938
rect 16210 13903 16212 13912
rect 15844 13874 15896 13880
rect 16264 13903 16266 13912
rect 16212 13874 16264 13880
rect 15856 13297 15884 13874
rect 16224 13462 16252 13874
rect 16316 13530 16344 14334
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 15842 13288 15898 13297
rect 16224 13274 16252 13398
rect 16224 13246 16344 13274
rect 15842 13223 15898 13232
rect 15856 12345 15884 13223
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 16316 12918 16344 13246
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16224 12782 16252 12854
rect 16408 12850 16436 14214
rect 16500 13274 16528 14214
rect 16592 13546 16620 17167
rect 16672 17138 16724 17144
rect 16684 15570 16712 17138
rect 17512 16561 17540 17478
rect 17498 16552 17554 16561
rect 17498 16487 17554 16496
rect 17512 15638 17540 16487
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 15094 16712 15506
rect 16776 15162 16804 15574
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 14482 18000 15030
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 14074 18000 14418
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17868 13864 17920 13870
rect 17222 13832 17278 13841
rect 16764 13796 16816 13802
rect 17868 13806 17920 13812
rect 17222 13767 17278 13776
rect 16764 13738 16816 13744
rect 16592 13518 16712 13546
rect 16776 13530 16804 13738
rect 17130 13560 17186 13569
rect 16580 13320 16632 13326
rect 16500 13268 16580 13274
rect 16500 13262 16632 13268
rect 16500 13246 16620 13262
rect 16684 13002 16712 13518
rect 16764 13524 16816 13530
rect 17236 13530 17264 13767
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17130 13495 17186 13504
rect 17224 13524 17276 13530
rect 16764 13466 16816 13472
rect 17144 13462 17172 13495
rect 17224 13466 17276 13472
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 16500 12986 16712 13002
rect 16488 12980 16712 12986
rect 16540 12974 16712 12980
rect 16488 12922 16540 12928
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16500 12481 16528 12786
rect 16486 12472 16542 12481
rect 16486 12407 16542 12416
rect 16500 12374 16528 12407
rect 16488 12368 16540 12374
rect 15842 12336 15898 12345
rect 16488 12310 16540 12316
rect 15842 12271 15898 12280
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9722 15884 10066
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15750 9616 15806 9625
rect 15750 9551 15806 9560
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 15658 8392 15714 8401
rect 15658 8327 15714 8336
rect 16212 8356 16264 8362
rect 15672 7002 15700 8327
rect 16212 8298 16264 8304
rect 16224 7993 16252 8298
rect 16210 7984 16266 7993
rect 16210 7919 16266 7928
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15672 6458 15700 6938
rect 16132 6866 16160 7142
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15764 6662 15792 6734
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15764 5914 15792 6598
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15382 5128 15438 5137
rect 15382 5063 15438 5072
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15028 3738 15056 4014
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 13740 2514 13860 2530
rect 13740 2508 13872 2514
rect 13740 2502 13820 2508
rect 13820 2450 13872 2456
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13464 480 13492 2382
rect 14936 480 14964 2858
rect 16316 2553 16344 8502
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8090 16528 8298
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16592 7449 16620 12974
rect 17144 12918 17172 13398
rect 17236 12986 17264 13466
rect 17328 13326 17356 13670
rect 17880 13530 17908 13806
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 16948 12776 17000 12782
rect 16946 12744 16948 12753
rect 17144 12753 17172 12854
rect 17000 12744 17002 12753
rect 16946 12679 17002 12688
rect 17130 12744 17186 12753
rect 17130 12679 17186 12688
rect 17328 12442 17356 13262
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11558 17172 12174
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11257 17172 11494
rect 17236 11286 17264 12038
rect 17512 11898 17540 12242
rect 17592 12232 17644 12238
rect 17590 12200 17592 12209
rect 17776 12232 17828 12238
rect 17644 12200 17646 12209
rect 17776 12174 17828 12180
rect 17590 12135 17646 12144
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17788 11626 17816 12174
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17224 11280 17276 11286
rect 17130 11248 17186 11257
rect 17224 11222 17276 11228
rect 17130 11183 17186 11192
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 7954 16712 9318
rect 16868 9178 16896 11018
rect 16960 10470 16988 11086
rect 17236 10742 17264 11222
rect 17328 10810 17356 11290
rect 17788 11082 17816 11562
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17788 10810 17816 11018
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 9926 16988 10406
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16868 8430 16896 9114
rect 17420 8974 17448 9862
rect 17788 9722 17816 10746
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17880 9926 17908 10678
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9518 17908 9862
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17868 9376 17920 9382
rect 17972 9364 18000 11630
rect 18064 10010 18092 20742
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 19720 20058 19748 20266
rect 20456 20058 20484 20334
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18340 19378 18368 19926
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18340 19174 18368 19314
rect 19154 19272 19210 19281
rect 18604 19236 18656 19242
rect 19154 19207 19210 19216
rect 18604 19178 18656 19184
rect 18328 19168 18380 19174
rect 18616 19145 18644 19178
rect 18696 19168 18748 19174
rect 18328 19110 18380 19116
rect 18602 19136 18658 19145
rect 18340 18902 18368 19110
rect 18696 19110 18748 19116
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18602 19071 18658 19080
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18340 18358 18368 18838
rect 18708 18834 18736 19110
rect 18800 18970 18828 19110
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18708 18426 18736 18770
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18892 18426 18920 18702
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18340 17610 18368 18294
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18510 17776 18566 17785
rect 18510 17711 18566 17720
rect 18328 17604 18380 17610
rect 18328 17546 18380 17552
rect 18340 17338 18368 17546
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16658 18184 17138
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18156 16250 18184 16594
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18432 16114 18460 16594
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18524 15994 18552 17711
rect 18432 15966 18552 15994
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18248 14482 18276 15302
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18248 13734 18276 14418
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13258 18276 13670
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18340 12646 18368 13262
rect 18328 12640 18380 12646
rect 18326 12608 18328 12617
rect 18380 12608 18382 12617
rect 18326 12543 18382 12552
rect 18432 10198 18460 15966
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18524 10985 18552 11086
rect 18510 10976 18566 10985
rect 18510 10911 18566 10920
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18142 10024 18198 10033
rect 18064 9982 18142 10010
rect 18524 10010 18552 10911
rect 18616 10169 18644 18022
rect 18892 17882 18920 18362
rect 19168 18154 19196 19207
rect 19720 18766 19748 19994
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 21560 18766 21588 20538
rect 22296 20398 22324 20878
rect 22388 20602 22416 20946
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22480 20058 22508 23520
rect 25502 23080 25558 23089
rect 25502 23015 25558 23024
rect 24858 22400 24914 22409
rect 24858 22335 24914 22344
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 23492 19854 23520 20266
rect 23584 19922 23612 20742
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 19310 23520 19790
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23584 19174 23612 19858
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 19720 18426 19748 18702
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 20456 18222 20484 18566
rect 21284 18358 21312 18634
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 19340 18216 19392 18222
rect 19260 18164 19340 18170
rect 19260 18158 19392 18164
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19260 18142 19380 18158
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 19168 17814 19196 18090
rect 19260 17882 19288 18142
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 20628 17876 20680 17882
rect 20732 17864 20760 18022
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21284 17882 21312 18294
rect 20680 17836 20760 17864
rect 21272 17876 21324 17882
rect 20628 17818 20680 17824
rect 21272 17818 21324 17824
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19062 16280 19118 16289
rect 19062 16215 19118 16224
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18878 15872 18934 15881
rect 18878 15807 18934 15816
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18708 13161 18736 13330
rect 18694 13152 18750 13161
rect 18694 13087 18750 13096
rect 18708 12782 18736 13087
rect 18892 12866 18920 15807
rect 18984 15162 19012 15982
rect 19076 15881 19104 16215
rect 19062 15872 19118 15881
rect 19062 15807 19118 15816
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 19076 14958 19104 15302
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18984 12986 19012 13194
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18892 12838 19012 12866
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18878 12064 18934 12073
rect 18878 11999 18934 12008
rect 18786 11656 18842 11665
rect 18786 11591 18842 11600
rect 18800 11354 18828 11591
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18800 11257 18828 11290
rect 18786 11248 18842 11257
rect 18786 11183 18842 11192
rect 18800 10810 18828 11183
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18892 10606 18920 11999
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18984 10266 19012 12838
rect 19076 12073 19104 14894
rect 19168 13705 19196 17750
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19352 17377 19380 17682
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19338 17368 19394 17377
rect 19338 17303 19340 17312
rect 19392 17303 19394 17312
rect 19340 17274 19392 17280
rect 19720 17066 19748 17614
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19996 17202 20024 17546
rect 20640 17338 20668 17818
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19522 16144 19578 16153
rect 19522 16079 19578 16088
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 13977 19380 14214
rect 19338 13968 19394 13977
rect 19338 13903 19394 13912
rect 19154 13696 19210 13705
rect 19154 13631 19210 13640
rect 19444 12753 19472 15846
rect 19536 15706 19564 16079
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19536 14958 19564 15642
rect 19524 14952 19576 14958
rect 19628 14929 19656 15846
rect 19720 15094 19748 17002
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19812 16658 19840 16934
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19904 16250 19932 16934
rect 19996 16794 20024 17138
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 20456 16114 20484 16390
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 19996 15366 20024 16050
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20258 15464 20314 15473
rect 20258 15399 20314 15408
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 19708 15088 19760 15094
rect 19708 15030 19760 15036
rect 19996 15026 20024 15302
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19524 14894 19576 14900
rect 19614 14920 19670 14929
rect 19614 14855 19670 14864
rect 19892 14884 19944 14890
rect 19628 13841 19656 14855
rect 19892 14826 19944 14832
rect 19904 13954 19932 14826
rect 19996 14278 20024 14962
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19996 14074 20024 14214
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19904 13926 20024 13954
rect 19614 13832 19670 13841
rect 19614 13767 19670 13776
rect 19430 12744 19486 12753
rect 19430 12679 19486 12688
rect 19248 12096 19300 12102
rect 19062 12064 19118 12073
rect 19248 12038 19300 12044
rect 19062 11999 19118 12008
rect 19260 11762 19288 12038
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11150 19104 11494
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18788 10192 18840 10198
rect 18602 10160 18658 10169
rect 18788 10134 18840 10140
rect 18602 10095 18658 10104
rect 18142 9959 18144 9968
rect 18196 9959 18198 9968
rect 18432 9982 18552 10010
rect 18144 9930 18196 9936
rect 18156 9518 18184 9930
rect 18432 9926 18460 9982
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18144 9512 18196 9518
rect 18432 9489 18460 9862
rect 18524 9586 18552 9862
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18144 9454 18196 9460
rect 18418 9480 18474 9489
rect 18418 9415 18474 9424
rect 17920 9336 18000 9364
rect 18236 9376 18288 9382
rect 17868 9318 17920 9324
rect 18236 9318 18288 9324
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16960 8362 16988 8774
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 17420 8294 17448 8910
rect 17880 8634 17908 9114
rect 18248 9042 18276 9318
rect 18616 9081 18644 10095
rect 18800 9110 18828 10134
rect 18984 9722 19012 10202
rect 19168 10062 19196 11562
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 19168 9586 19196 9998
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 18788 9104 18840 9110
rect 18602 9072 18658 9081
rect 18236 9036 18288 9042
rect 18788 9046 18840 9052
rect 18602 9007 18658 9016
rect 18236 8978 18288 8984
rect 18248 8634 18276 8978
rect 19076 8974 19104 9522
rect 19168 9042 19196 9522
rect 19812 9518 19840 9862
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19708 9376 19760 9382
rect 19706 9344 19708 9353
rect 19760 9344 19762 9353
rect 19706 9279 19762 9288
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19076 8634 19104 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7954 17448 8230
rect 17880 8106 17908 8434
rect 19812 8265 19840 9454
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 9178 19932 9318
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 19904 8634 19932 9114
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19798 8256 19854 8265
rect 19854 8214 19932 8242
rect 19798 8191 19854 8200
rect 17880 8090 18000 8106
rect 17880 8084 18012 8090
rect 17880 8078 17960 8084
rect 17960 8026 18012 8032
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 16684 7478 16712 7890
rect 16776 7546 16804 7890
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16672 7472 16724 7478
rect 16578 7440 16634 7449
rect 16672 7414 16724 7420
rect 16578 7375 16634 7384
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5846 16436 6054
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16684 5658 16712 7414
rect 19168 7274 19196 7686
rect 19536 7410 19564 7754
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17224 6792 17276 6798
rect 17222 6760 17224 6769
rect 17276 6760 17278 6769
rect 17222 6695 17278 6704
rect 16948 6656 17000 6662
rect 16854 6624 16910 6633
rect 16948 6598 17000 6604
rect 16854 6559 16910 6568
rect 16868 6254 16896 6559
rect 16856 6248 16908 6254
rect 16762 6216 16818 6225
rect 16856 6190 16908 6196
rect 16762 6151 16764 6160
rect 16816 6151 16818 6160
rect 16764 6122 16816 6128
rect 16868 5914 16896 6190
rect 16960 5914 16988 6598
rect 17236 6390 17264 6695
rect 17328 6458 17356 6802
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17696 5914 17724 6666
rect 19260 5930 19288 7142
rect 19536 6934 19564 7346
rect 19812 7002 19840 7822
rect 19904 7585 19932 8214
rect 19996 8106 20024 13926
rect 20088 13410 20116 14894
rect 20180 14113 20208 15302
rect 20272 14890 20300 15399
rect 20732 15162 20760 15506
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20824 15065 20852 15846
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20810 15056 20866 15065
rect 20810 14991 20866 15000
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20166 14104 20222 14113
rect 20166 14039 20222 14048
rect 20180 13870 20208 14039
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20444 13864 20496 13870
rect 20496 13812 20576 13818
rect 20444 13806 20576 13812
rect 20180 13530 20208 13806
rect 20456 13790 20576 13806
rect 20548 13682 20576 13790
rect 20548 13654 20668 13682
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20088 13382 20300 13410
rect 20166 13016 20222 13025
rect 20166 12951 20222 12960
rect 20180 9926 20208 12951
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20088 8634 20116 9046
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20074 8120 20130 8129
rect 19996 8078 20074 8106
rect 20074 8055 20076 8064
rect 20128 8055 20130 8064
rect 20076 8026 20128 8032
rect 19890 7576 19946 7585
rect 20088 7546 20116 8026
rect 19890 7511 19946 7520
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 19168 5902 19380 5930
rect 16592 5630 16712 5658
rect 16764 5704 16816 5710
rect 16868 5681 16896 5850
rect 16764 5646 16816 5652
rect 16854 5672 16910 5681
rect 16488 4684 16540 4690
rect 16592 4672 16620 5630
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16540 4644 16620 4672
rect 16488 4626 16540 4632
rect 16592 3942 16620 4644
rect 16684 4078 16712 5510
rect 16776 5370 16804 5646
rect 16854 5607 16910 5616
rect 16960 5370 16988 5850
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16776 4758 16804 5306
rect 17144 5302 17172 5782
rect 19168 5370 19196 5902
rect 19352 5846 19380 5902
rect 19708 5908 19760 5914
rect 19708 5850 19760 5856
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16302 2544 16358 2553
rect 16408 2514 16436 3878
rect 16684 3738 16712 4014
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16776 3670 16804 4694
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 16868 4146 16896 4422
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16764 3664 16816 3670
rect 17880 3652 17908 4422
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 17960 3664 18012 3670
rect 17880 3624 17960 3652
rect 16764 3606 16816 3612
rect 17960 3606 18012 3612
rect 17972 3194 18000 3606
rect 18156 3602 18184 3878
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18156 3126 18184 3538
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 19260 2650 19288 5510
rect 19720 5370 19748 5850
rect 19890 5808 19946 5817
rect 19890 5743 19946 5752
rect 19904 5710 19932 5743
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19904 5302 19932 5646
rect 20272 5370 20300 13382
rect 20640 10826 20668 13654
rect 20718 12744 20774 12753
rect 20718 12679 20774 12688
rect 20732 12073 20760 12679
rect 20824 12617 20852 14991
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 21270 12744 21326 12753
rect 21270 12679 21326 12688
rect 20810 12608 20866 12617
rect 20810 12543 20866 12552
rect 20718 12064 20774 12073
rect 20718 11999 20774 12008
rect 20640 10810 20760 10826
rect 20640 10804 20772 10810
rect 20640 10798 20720 10804
rect 20720 10746 20772 10752
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20640 10130 20668 10678
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20364 9178 20392 9522
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20456 8106 20484 9862
rect 20640 9722 20668 10066
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20548 8537 20576 9386
rect 20534 8528 20590 8537
rect 20534 8463 20590 8472
rect 20364 8078 20484 8106
rect 20364 7750 20392 8078
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20364 7342 20392 7686
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 20272 5030 20300 5306
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20364 4078 20392 7278
rect 20456 7206 20484 7890
rect 20732 7290 20760 10406
rect 20824 7750 20852 12543
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 21284 12374 21312 12679
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21284 11898 21312 12310
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21284 8945 21312 9318
rect 21270 8936 21326 8945
rect 21270 8871 21326 8880
rect 21284 8401 21312 8871
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 21270 7984 21326 7993
rect 21270 7919 21272 7928
rect 21324 7919 21326 7928
rect 21272 7890 21324 7896
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 21376 7562 21404 18566
rect 21560 18426 21588 18702
rect 21836 18426 21864 18906
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 22756 18358 22784 18702
rect 22836 18624 22888 18630
rect 22836 18566 22888 18572
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22204 17814 22232 18090
rect 22848 17882 22876 18566
rect 23216 18426 23244 18770
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23308 17882 23336 18770
rect 23480 18216 23532 18222
rect 23478 18184 23480 18193
rect 23532 18184 23534 18193
rect 23478 18119 23534 18128
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 16250 21496 16526
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15366 21772 15846
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21744 13705 21772 15302
rect 21730 13696 21786 13705
rect 21730 13631 21786 13640
rect 21744 13161 21772 13631
rect 21730 13152 21786 13161
rect 21730 13087 21786 13096
rect 21638 12064 21694 12073
rect 21638 11999 21694 12008
rect 21548 9444 21600 9450
rect 21548 9386 21600 9392
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21468 9110 21496 9318
rect 21560 9178 21588 9386
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21456 9104 21508 9110
rect 21456 9046 21508 9052
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 20548 7262 20760 7290
rect 20824 7534 21404 7562
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20456 7041 20484 7142
rect 20442 7032 20498 7041
rect 20442 6967 20498 6976
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20364 3738 20392 4014
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20548 3194 20576 7262
rect 20628 7200 20680 7206
rect 20680 7148 20760 7154
rect 20628 7142 20760 7148
rect 20640 7126 20760 7142
rect 20732 6730 20760 7126
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20732 5370 20760 5714
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20732 4826 20760 5102
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20824 4672 20852 7534
rect 21468 7290 21496 7822
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21376 7274 21496 7290
rect 21364 7268 21496 7274
rect 21416 7262 21496 7268
rect 21364 7210 21416 7216
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 21008 6458 21036 6666
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21192 6338 21220 6802
rect 21284 6458 21312 6938
rect 21376 6934 21404 7210
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21192 6310 21312 6338
rect 21284 6118 21312 6310
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 21284 5574 21312 6054
rect 21468 5710 21496 7142
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21284 5234 21312 5510
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 20732 4644 20852 4672
rect 20732 3618 20760 4644
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20824 3738 20852 4490
rect 21008 4214 21036 4490
rect 21192 4282 21220 4694
rect 21284 4554 21312 5170
rect 21376 5098 21404 5646
rect 21468 5370 21496 5646
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21376 4826 21404 5034
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 21560 4758 21588 7686
rect 21548 4752 21600 4758
rect 21548 4694 21600 4700
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 21192 4049 21220 4218
rect 21178 4040 21234 4049
rect 21178 3975 21234 3984
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20732 3590 20852 3618
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 16302 2479 16358 2488
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 480 16344 2382
rect 17788 480 17816 2382
rect 19168 480 19196 2382
rect 20640 480 20668 2858
rect 20824 2650 20852 3590
rect 21284 3466 21312 3946
rect 21362 3768 21418 3777
rect 21362 3703 21364 3712
rect 21416 3703 21418 3712
rect 21364 3674 21416 3680
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 21284 2650 21312 3402
rect 21376 3194 21404 3674
rect 21652 3670 21680 11999
rect 21744 5166 21772 13087
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 10266 21864 12038
rect 21928 11558 21956 12242
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21928 11218 21956 11494
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 9586 21864 10202
rect 21928 9926 21956 11154
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21822 8800 21878 8809
rect 21822 8735 21878 8744
rect 21836 6730 21864 8735
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21928 5370 21956 5714
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21744 4729 21772 4966
rect 21730 4720 21786 4729
rect 21730 4655 21786 4664
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 21928 3942 21956 4490
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 22020 3754 22048 16934
rect 22112 16794 22140 17138
rect 22388 17134 22416 17818
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 22376 17128 22428 17134
rect 23216 17105 23244 17682
rect 22376 17070 22428 17076
rect 23202 17096 23258 17105
rect 23202 17031 23204 17040
rect 23256 17031 23258 17040
rect 23204 17002 23256 17008
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23492 16561 23520 16594
rect 23110 16552 23166 16561
rect 22744 16516 22796 16522
rect 23110 16487 23166 16496
rect 23478 16552 23534 16561
rect 23478 16487 23534 16496
rect 22744 16458 22796 16464
rect 22756 16250 22784 16458
rect 23124 16250 23152 16487
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22756 15609 22784 16186
rect 23124 16153 23152 16186
rect 23110 16144 23166 16153
rect 23110 16079 23166 16088
rect 22742 15600 22798 15609
rect 22742 15535 22798 15544
rect 23204 15564 23256 15570
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 15162 22692 15302
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22558 14784 22614 14793
rect 22558 14719 22614 14728
rect 22572 14414 22600 14719
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22572 14113 22600 14350
rect 22558 14104 22614 14113
rect 22664 14074 22692 14418
rect 22558 14039 22614 14048
rect 22652 14068 22704 14074
rect 22572 13734 22600 14039
rect 22652 14010 22704 14016
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22204 13326 22232 13670
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12986 22232 13262
rect 22572 12986 22600 13398
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22756 12306 22784 15535
rect 23204 15506 23256 15512
rect 23216 14822 23244 15506
rect 23584 15502 23612 19110
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24228 18290 24256 18906
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 23662 17776 23718 17785
rect 23662 17711 23664 17720
rect 23716 17711 23718 17720
rect 23664 17682 23716 17688
rect 24228 17678 24256 18226
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 23860 16726 23888 17614
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24136 17202 24164 17478
rect 24320 17202 24348 18702
rect 24412 18630 24440 19110
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24872 18306 24900 22335
rect 25226 21584 25282 21593
rect 25226 21519 25282 21528
rect 25134 20496 25190 20505
rect 25134 20431 25190 20440
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24964 19242 24992 19654
rect 24952 19236 25004 19242
rect 24952 19178 25004 19184
rect 24964 18970 24992 19178
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 24780 18278 24900 18306
rect 24780 18222 24808 18278
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24780 17649 24808 17682
rect 24766 17640 24822 17649
rect 24766 17575 24822 17584
rect 24780 17338 24808 17575
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24858 17232 24914 17241
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24308 17196 24360 17202
rect 24858 17167 24914 17176
rect 24308 17138 24360 17144
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24044 16794 24072 17002
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23848 16720 23900 16726
rect 23848 16662 23900 16668
rect 23860 16590 23888 16662
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 16182 23888 16526
rect 24136 16250 24164 17138
rect 24320 16794 24348 17138
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23860 15638 23888 16118
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23848 15632 23900 15638
rect 23848 15574 23900 15580
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23308 14958 23336 15370
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23216 13025 23244 14758
rect 23202 13016 23258 13025
rect 23202 12951 23258 12960
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22204 10470 22232 10950
rect 22848 10810 22876 11154
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22192 10464 22244 10470
rect 22190 10432 22192 10441
rect 22284 10464 22336 10470
rect 22244 10432 22246 10441
rect 22284 10406 22336 10412
rect 22190 10367 22246 10376
rect 22296 10266 22324 10406
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22848 10146 22876 10746
rect 22744 10124 22796 10130
rect 22848 10118 22968 10146
rect 22744 10066 22796 10072
rect 22756 9654 22784 10066
rect 22940 10062 22968 10118
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22756 9110 22784 9590
rect 22848 9178 22876 9998
rect 22940 9722 22968 9998
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22664 6633 22692 8434
rect 23216 8090 23244 9046
rect 23308 8537 23336 14894
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23492 13546 23520 13942
rect 23400 13518 23520 13546
rect 23400 13462 23428 13518
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23492 12753 23520 13126
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23478 12744 23534 12753
rect 23478 12679 23480 12688
rect 23532 12679 23534 12688
rect 23480 12650 23532 12656
rect 23860 12442 23888 12786
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10674 23428 10950
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23584 9926 23612 10406
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23584 9586 23612 9862
rect 23754 9616 23810 9625
rect 23572 9580 23624 9586
rect 23754 9551 23810 9560
rect 23572 9522 23624 9528
rect 23400 9042 23520 9058
rect 23388 9036 23520 9042
rect 23440 9030 23520 9036
rect 23388 8978 23440 8984
rect 23294 8528 23350 8537
rect 23294 8463 23350 8472
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 23124 7585 23152 7890
rect 23308 7886 23336 8463
rect 23492 8294 23520 9030
rect 23584 8974 23612 9522
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23584 8566 23612 8910
rect 23676 8634 23704 9386
rect 23768 9382 23796 9551
rect 23860 9518 23888 12242
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23860 9042 23888 9454
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23754 8936 23810 8945
rect 23952 8922 23980 15914
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24136 15706 24164 15846
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24306 15056 24362 15065
rect 24306 14991 24308 15000
rect 24360 14991 24362 15000
rect 24308 14962 24360 14968
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24044 14006 24072 14214
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 24504 13938 24532 14758
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24504 13530 24532 13874
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 12850 24348 13126
rect 24688 12918 24716 13670
rect 24872 13258 24900 17167
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24228 10266 24256 10542
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24228 9994 24256 10202
rect 24216 9988 24268 9994
rect 24216 9930 24268 9936
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 23810 8894 23980 8922
rect 23754 8871 23810 8880
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23110 7576 23166 7585
rect 23492 7546 23520 8230
rect 23110 7511 23112 7520
rect 23164 7511 23166 7520
rect 23480 7540 23532 7546
rect 23112 7482 23164 7488
rect 23480 7482 23532 7488
rect 23124 7451 23152 7482
rect 23768 7206 23796 8871
rect 23938 8528 23994 8537
rect 23938 8463 23940 8472
rect 23992 8463 23994 8472
rect 23940 8434 23992 8440
rect 23952 8362 23980 8434
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23860 7274 23888 7822
rect 24044 7342 24072 8978
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24136 8498 24164 8774
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24228 8401 24256 9318
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23768 6662 23796 7142
rect 24044 7002 24072 7278
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 23756 6656 23808 6662
rect 22650 6624 22706 6633
rect 23756 6598 23808 6604
rect 22650 6559 22706 6568
rect 22928 6248 22980 6254
rect 22928 6190 22980 6196
rect 22940 5846 22968 6190
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 5914 23520 6054
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 22928 5840 22980 5846
rect 23492 5817 23520 5850
rect 22928 5782 22980 5788
rect 23478 5808 23534 5817
rect 22940 5370 22968 5782
rect 23478 5743 23534 5752
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22940 4214 22968 5306
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 21928 3726 22048 3754
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 21652 3194 21680 3606
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21928 2666 21956 3726
rect 23768 3097 23796 6598
rect 24320 3194 24348 12650
rect 24872 12442 24900 12718
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24964 12322 24992 16186
rect 25148 13530 25176 20431
rect 25240 18873 25268 21519
rect 25318 21312 25374 21321
rect 25318 21247 25374 21256
rect 25226 18864 25282 18873
rect 25226 18799 25282 18808
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25240 15201 25268 18362
rect 25226 15192 25282 15201
rect 25226 15127 25282 15136
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25240 14278 25268 14962
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 14074 25268 14214
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25136 13524 25188 13530
rect 25136 13466 25188 13472
rect 25240 13410 25268 13874
rect 25148 13382 25268 13410
rect 25042 12472 25098 12481
rect 25042 12407 25098 12416
rect 24872 12294 24992 12322
rect 24872 10554 24900 12294
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24964 11898 24992 12174
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25056 11801 25084 12407
rect 25148 12238 25176 13382
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25042 11792 25098 11801
rect 25042 11727 25098 11736
rect 24872 10526 24992 10554
rect 24858 10432 24914 10441
rect 24858 10367 24914 10376
rect 24872 10266 24900 10367
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24872 9722 24900 9998
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24584 8356 24636 8362
rect 24584 8298 24636 8304
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24596 6361 24624 8298
rect 24688 7886 24716 8298
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7410 24716 7822
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24688 7206 24716 7346
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24688 6662 24716 7142
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24582 6352 24638 6361
rect 24582 6287 24638 6296
rect 24596 6066 24624 6287
rect 24780 6254 24808 8026
rect 24964 6905 24992 10526
rect 25240 10248 25268 13262
rect 25332 12617 25360 21247
rect 25410 20088 25466 20097
rect 25410 20023 25466 20032
rect 25424 16250 25452 20023
rect 25516 18426 25544 23015
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25502 18320 25558 18329
rect 25502 18255 25558 18264
rect 25516 17241 25544 18255
rect 25502 17232 25558 17241
rect 25502 17167 25558 17176
rect 25502 16960 25558 16969
rect 25502 16895 25558 16904
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25410 15056 25466 15065
rect 25410 14991 25466 15000
rect 25318 12608 25374 12617
rect 25318 12543 25374 12552
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25332 11898 25360 12378
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25148 10220 25268 10248
rect 25320 10260 25372 10266
rect 25148 8809 25176 10220
rect 25320 10202 25372 10208
rect 25332 9722 25360 10202
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25134 8800 25190 8809
rect 25134 8735 25190 8744
rect 25424 8537 25452 14991
rect 25516 14521 25544 16895
rect 25502 14512 25558 14521
rect 25502 14447 25558 14456
rect 25502 12880 25558 12889
rect 25502 12815 25504 12824
rect 25556 12815 25558 12824
rect 25504 12786 25556 12792
rect 25608 12730 25636 23559
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26238 20360 26294 20369
rect 26238 20295 26294 20304
rect 26252 20262 26280 20295
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 27528 20256 27580 20262
rect 27580 20204 27660 20210
rect 27528 20198 27660 20204
rect 27540 20182 27660 20198
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18766 25728 19110
rect 25870 18864 25926 18873
rect 25870 18799 25926 18808
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25700 18290 25728 18702
rect 25780 18624 25832 18630
rect 25780 18566 25832 18572
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25700 18154 25728 18226
rect 25688 18148 25740 18154
rect 25688 18090 25740 18096
rect 25792 18086 25820 18566
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25792 17626 25820 18022
rect 25700 17598 25820 17626
rect 25700 17542 25728 17598
rect 25688 17536 25740 17542
rect 25688 17478 25740 17484
rect 25700 17066 25728 17478
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25700 16454 25728 17002
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25700 15366 25728 16390
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 14793 25728 15302
rect 25780 14952 25832 14958
rect 25778 14920 25780 14929
rect 25832 14920 25834 14929
rect 25778 14855 25834 14864
rect 25686 14784 25742 14793
rect 25686 14719 25742 14728
rect 25686 14648 25742 14657
rect 25686 14583 25742 14592
rect 25700 13433 25728 14583
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25686 13424 25742 13433
rect 25686 13359 25742 13368
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12782 25728 13194
rect 25516 12702 25636 12730
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 25516 12209 25544 12702
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25792 12594 25820 14447
rect 25884 12714 25912 18799
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 27172 17134 27200 18022
rect 27160 17128 27212 17134
rect 26514 17096 26570 17105
rect 27160 17070 27212 17076
rect 26514 17031 26570 17040
rect 26528 16658 26556 17031
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 26344 15042 26372 15302
rect 26160 15014 26372 15042
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 26068 14793 26096 14894
rect 26160 14890 26188 15014
rect 26148 14884 26200 14890
rect 26148 14826 26200 14832
rect 26332 14884 26384 14890
rect 26332 14826 26384 14832
rect 26054 14784 26110 14793
rect 26054 14719 26110 14728
rect 26344 14618 26372 14826
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26436 14113 26464 16458
rect 26528 16250 26556 16594
rect 26606 16552 26662 16561
rect 26606 16487 26662 16496
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26422 14104 26478 14113
rect 26422 14039 26478 14048
rect 26054 13968 26110 13977
rect 26054 13903 26056 13912
rect 26108 13903 26110 13912
rect 26332 13932 26384 13938
rect 26056 13874 26108 13880
rect 26332 13874 26384 13880
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26252 13705 26280 13806
rect 26344 13802 26372 13874
rect 26332 13796 26384 13802
rect 26332 13738 26384 13744
rect 26238 13696 26294 13705
rect 26238 13631 26294 13640
rect 26252 13530 26280 13631
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26252 13433 26280 13466
rect 26238 13424 26294 13433
rect 26238 13359 26294 13368
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26344 12866 26372 13126
rect 26160 12838 26372 12866
rect 25872 12708 25924 12714
rect 25872 12650 25924 12656
rect 25700 12442 25728 12582
rect 25792 12566 25912 12594
rect 25778 12472 25834 12481
rect 25688 12436 25740 12442
rect 25778 12407 25834 12416
rect 25688 12378 25740 12384
rect 25596 12368 25648 12374
rect 25596 12310 25648 12316
rect 25502 12200 25558 12209
rect 25502 12135 25558 12144
rect 25608 11898 25636 12310
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25792 10985 25820 12407
rect 25778 10976 25834 10985
rect 25778 10911 25834 10920
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25608 10062 25636 10406
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25700 9382 25728 10066
rect 25792 9654 25820 10911
rect 25884 10441 25912 12566
rect 26160 12374 26188 12838
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26148 12368 26200 12374
rect 26148 12310 26200 12316
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25870 10432 25926 10441
rect 25870 10367 25926 10376
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 25780 9648 25832 9654
rect 25780 9590 25832 9596
rect 25792 9450 25820 9590
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25700 9178 25728 9318
rect 25976 9178 26004 9454
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 26344 9058 26372 12038
rect 26436 11694 26464 12718
rect 26514 12336 26570 12345
rect 26514 12271 26516 12280
rect 26568 12271 26570 12280
rect 26516 12242 26568 12248
rect 26528 11898 26556 12242
rect 26620 11914 26648 16487
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26712 14521 26740 16390
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26698 14512 26754 14521
rect 26698 14447 26754 14456
rect 26804 14278 26832 15506
rect 27356 15502 27384 16934
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 26988 14929 27016 15438
rect 26974 14920 27030 14929
rect 26974 14855 27030 14864
rect 27250 14920 27306 14929
rect 27250 14855 27306 14864
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26712 12782 26740 13262
rect 26700 12776 26752 12782
rect 26698 12744 26700 12753
rect 26752 12744 26754 12753
rect 26698 12679 26754 12688
rect 26804 12209 26832 14214
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 26884 13388 26936 13394
rect 26884 13330 26936 13336
rect 26896 12986 26924 13330
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26790 12200 26846 12209
rect 26790 12135 26846 12144
rect 26516 11892 26568 11898
rect 26620 11886 26832 11914
rect 26516 11834 26568 11840
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26698 11656 26754 11665
rect 26698 11591 26754 11600
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26514 11248 26570 11257
rect 26514 11183 26516 11192
rect 26568 11183 26570 11192
rect 26516 11154 26568 11160
rect 26528 10810 26556 11154
rect 26620 11121 26648 11494
rect 26712 11354 26740 11591
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26606 11112 26662 11121
rect 26606 11047 26662 11056
rect 26516 10804 26568 10810
rect 26516 10746 26568 10752
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26436 9586 26464 9862
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26436 9110 26464 9522
rect 26620 9518 26648 10406
rect 26698 9888 26754 9897
rect 26698 9823 26754 9832
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26712 9178 26740 9823
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 25884 9030 26372 9058
rect 26424 9104 26476 9110
rect 26424 9046 26476 9052
rect 26514 9072 26570 9081
rect 25410 8528 25466 8537
rect 25410 8463 25466 8472
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 25608 8090 25636 8366
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 24950 6896 25006 6905
rect 24950 6831 25006 6840
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24596 6038 24900 6066
rect 24872 3602 24900 6038
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24308 3188 24360 3194
rect 24308 3130 24360 3136
rect 23754 3088 23810 3097
rect 23754 3023 23810 3032
rect 24320 2990 24348 3130
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21272 2644 21324 2650
rect 21928 2638 22140 2666
rect 21272 2586 21324 2592
rect 22112 2514 22140 2638
rect 24306 2544 24362 2553
rect 22100 2508 22152 2514
rect 24306 2479 24308 2488
rect 22100 2450 22152 2456
rect 24360 2479 24362 2488
rect 24308 2450 24360 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 22020 480 22048 2382
rect 23492 480 23520 2382
rect 24872 480 24900 2858
rect 25148 2514 25176 7210
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25332 6458 25360 6598
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25884 5273 25912 9030
rect 26514 9007 26516 9016
rect 26568 9007 26570 9016
rect 26516 8978 26568 8984
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26528 8634 26556 8978
rect 26698 8664 26754 8673
rect 26516 8628 26568 8634
rect 26698 8599 26754 8608
rect 26516 8570 26568 8576
rect 26330 8392 26386 8401
rect 26330 8327 26386 8336
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26344 6866 26372 8327
rect 26606 8120 26662 8129
rect 26712 8090 26740 8599
rect 26606 8055 26662 8064
rect 26700 8084 26752 8090
rect 26514 7984 26570 7993
rect 26514 7919 26516 7928
rect 26568 7919 26570 7928
rect 26516 7890 26568 7896
rect 26528 7478 26556 7890
rect 26620 7546 26648 8055
rect 26700 8026 26752 8032
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26516 7472 26568 7478
rect 26516 7414 26568 7420
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26436 6225 26464 7278
rect 26698 6896 26754 6905
rect 26698 6831 26754 6840
rect 26712 6730 26740 6831
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26608 6384 26660 6390
rect 26606 6352 26608 6361
rect 26660 6352 26662 6361
rect 26606 6287 26662 6296
rect 26422 6216 26478 6225
rect 26422 6151 26478 6160
rect 26804 5778 26832 11886
rect 26974 10704 27030 10713
rect 26974 10639 27030 10648
rect 26988 10266 27016 10639
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26896 10033 26924 10066
rect 26882 10024 26938 10033
rect 26882 9959 26938 9968
rect 26896 9722 26924 9959
rect 26988 9722 27016 10202
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 26896 9518 26924 9658
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 26988 8566 27016 9046
rect 26976 8560 27028 8566
rect 26976 8502 27028 8508
rect 27172 6458 27200 13738
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 26698 5672 26754 5681
rect 26698 5607 26700 5616
rect 26752 5607 26754 5616
rect 26700 5578 26752 5584
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26804 5370 26832 5714
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 25870 5264 25926 5273
rect 25870 5199 25926 5208
rect 26424 5160 26476 5166
rect 26422 5128 26424 5137
rect 26476 5128 26478 5137
rect 26422 5063 26478 5072
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26514 4720 26570 4729
rect 26514 4655 26516 4664
rect 26568 4655 26570 4664
rect 26516 4626 26568 4632
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26528 4282 26556 4626
rect 26620 4457 26648 4966
rect 26700 4480 26752 4486
rect 26606 4448 26662 4457
rect 26700 4422 26752 4428
rect 26606 4383 26662 4392
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26712 4185 26740 4422
rect 26698 4176 26754 4185
rect 26698 4111 26754 4120
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26514 4040 26570 4049
rect 26436 3641 26464 4014
rect 26514 3975 26570 3984
rect 26422 3632 26478 3641
rect 25320 3596 25372 3602
rect 26528 3602 26556 3975
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26422 3567 26478 3576
rect 26516 3596 26568 3602
rect 25320 3538 25372 3544
rect 26516 3538 26568 3544
rect 25332 3194 25360 3538
rect 25502 3496 25558 3505
rect 25502 3431 25504 3440
rect 25556 3431 25558 3440
rect 25504 3402 25556 3408
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26528 3194 26556 3538
rect 26700 3392 26752 3398
rect 26700 3334 26752 3340
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 921 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 912 25926 921
rect 25870 847 25926 856
rect 26344 480 26372 2382
rect 3974 368 4030 377
rect 3974 303 4030 312
rect 4894 0 4950 480
rect 6366 0 6422 480
rect 7746 0 7802 480
rect 9218 0 9274 480
rect 10598 0 10654 480
rect 12070 0 12126 480
rect 13450 0 13506 480
rect 14922 0 14978 480
rect 16302 0 16358 480
rect 17774 0 17830 480
rect 19154 0 19210 480
rect 20626 0 20682 480
rect 22006 0 22062 480
rect 23478 0 23534 480
rect 24858 0 24914 480
rect 26330 0 26386 480
rect 26620 377 26648 2790
rect 26712 1465 26740 3334
rect 26804 2825 26832 3878
rect 27264 3777 27292 14855
rect 27356 14618 27384 15438
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27448 13938 27476 14758
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27448 13326 27476 13874
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27448 12782 27476 13262
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27448 12442 27476 12718
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27540 10713 27568 12650
rect 27526 10704 27582 10713
rect 27526 10639 27582 10648
rect 27632 9466 27660 20182
rect 27632 9438 27752 9466
rect 27620 9376 27672 9382
rect 27618 9344 27620 9353
rect 27672 9344 27674 9353
rect 27618 9279 27674 9288
rect 27724 7562 27752 9438
rect 27632 7534 27752 7562
rect 27526 7440 27582 7449
rect 27526 7375 27582 7384
rect 27540 7342 27568 7375
rect 27528 7336 27580 7342
rect 27528 7278 27580 7284
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27356 6458 27384 6802
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27250 3768 27306 3777
rect 27250 3703 27306 3712
rect 27264 3126 27292 3703
rect 27252 3120 27304 3126
rect 27252 3062 27304 3068
rect 27526 3088 27582 3097
rect 27632 3074 27660 7534
rect 27712 7472 27764 7478
rect 27710 7440 27712 7449
rect 27764 7440 27766 7449
rect 27710 7375 27766 7384
rect 27632 3046 27752 3074
rect 27526 3023 27582 3032
rect 27540 2990 27568 3023
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 26790 2816 26846 2825
rect 26790 2751 26846 2760
rect 26698 1456 26754 1465
rect 26698 1391 26754 1400
rect 27724 480 27752 3046
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27816 2145 27844 2790
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 27802 2136 27858 2145
rect 27802 2071 27858 2080
rect 29196 480 29224 2246
rect 26606 368 26662 377
rect 26606 303 26662 312
rect 27710 0 27766 480
rect 29182 0 29238 480
<< via2 >>
rect 3330 23568 3386 23624
rect 2410 22344 2466 22400
rect 2318 17740 2374 17776
rect 2318 17720 2320 17740
rect 2320 17720 2372 17740
rect 2372 17720 2374 17740
rect 3054 21800 3110 21856
rect 2870 21256 2926 21312
rect 2870 20032 2926 20088
rect 2686 17856 2742 17912
rect 2410 17448 2466 17504
rect 1490 14068 1546 14104
rect 1490 14048 1492 14068
rect 1492 14048 1544 14068
rect 1544 14048 1546 14068
rect 1950 14728 2006 14784
rect 1490 11600 1546 11656
rect 1582 11076 1638 11112
rect 1582 11056 1584 11076
rect 1584 11056 1636 11076
rect 1636 11056 1638 11076
rect 1398 10376 1454 10432
rect 1398 7384 1454 7440
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1582 8608 1638 8664
rect 1674 7284 1676 7304
rect 1676 7284 1728 7304
rect 1728 7284 1730 7304
rect 1674 7248 1730 7284
rect 1582 6840 1638 6896
rect 1582 6296 1638 6352
rect 1582 5616 1638 5672
rect 2778 12824 2834 12880
rect 2042 11212 2098 11248
rect 2042 11192 2044 11212
rect 2044 11192 2096 11212
rect 2096 11192 2098 11212
rect 2410 10804 2466 10840
rect 2410 10784 2412 10804
rect 2412 10784 2464 10804
rect 2464 10784 2466 10804
rect 2778 10512 2834 10568
rect 3146 19352 3202 19408
rect 3146 17176 3202 17232
rect 25594 23568 25650 23624
rect 3422 23024 3478 23080
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 3882 20576 3938 20632
rect 3514 18264 3570 18320
rect 3054 14184 3110 14240
rect 3054 13912 3110 13968
rect 2962 13368 3018 13424
rect 2962 12824 3018 12880
rect 2870 10376 2926 10432
rect 2042 9444 2098 9480
rect 2042 9424 2044 9444
rect 2044 9424 2096 9444
rect 2096 9424 2098 9444
rect 2686 9832 2742 9888
rect 2042 9016 2098 9072
rect 2410 9560 2466 9616
rect 2686 8084 2742 8120
rect 2686 8064 2688 8084
rect 2688 8064 2740 8084
rect 2740 8064 2742 8084
rect 2502 7948 2558 7984
rect 2502 7928 2504 7948
rect 2504 7928 2556 7948
rect 2556 7928 2558 7948
rect 1858 6860 1914 6896
rect 1858 6840 1860 6860
rect 1860 6840 1912 6860
rect 1912 6840 1914 6860
rect 2410 5888 2466 5944
rect 2594 6024 2650 6080
rect 1766 5072 1822 5128
rect 1582 4392 1638 4448
rect 1398 4020 1400 4040
rect 1400 4020 1452 4040
rect 1452 4020 1454 4040
rect 1398 3984 1454 4020
rect 662 3712 718 3768
rect 2686 3848 2742 3904
rect 1582 1400 1638 1456
rect 3238 13268 3240 13288
rect 3240 13268 3292 13288
rect 3292 13268 3294 13288
rect 3238 13232 3294 13268
rect 3790 17040 3846 17096
rect 3606 14184 3662 14240
rect 3514 13912 3570 13968
rect 3422 11600 3478 11656
rect 3238 10104 3294 10160
rect 7470 20304 7526 20360
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 3974 18808 4030 18864
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 4066 17584 4122 17640
rect 3974 15952 4030 16008
rect 3882 15680 3938 15736
rect 3882 15272 3938 15328
rect 3790 13504 3846 13560
rect 3790 12552 3846 12608
rect 3514 7792 3570 7848
rect 3146 6976 3202 7032
rect 3054 6024 3110 6080
rect 2502 2352 2558 2408
rect 4066 14592 4122 14648
rect 4066 13368 4122 13424
rect 4066 11076 4122 11112
rect 4066 11056 4068 11076
rect 4068 11056 4120 11076
rect 4120 11056 4122 11076
rect 4250 8200 4306 8256
rect 4250 7928 4306 7984
rect 4250 6840 4306 6896
rect 3882 6296 3938 6352
rect 3606 4972 3608 4992
rect 3608 4972 3660 4992
rect 3660 4972 3662 4992
rect 3606 4936 3662 4972
rect 3606 3848 3662 3904
rect 3882 3304 3938 3360
rect 4250 5908 4306 5944
rect 4250 5888 4252 5908
rect 4252 5888 4304 5908
rect 4304 5888 4306 5908
rect 7470 17720 7526 17776
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 4710 16360 4766 16416
rect 4434 15580 4436 15600
rect 4436 15580 4488 15600
rect 4488 15580 4490 15600
rect 4434 15544 4490 15580
rect 4526 15444 4528 15464
rect 4528 15444 4580 15464
rect 4580 15444 4582 15464
rect 4526 15408 4582 15444
rect 4434 14068 4490 14104
rect 4434 14048 4436 14068
rect 4436 14048 4488 14068
rect 4488 14048 4490 14068
rect 7470 17312 7526 17368
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5722 15680 5778 15736
rect 6182 15700 6238 15736
rect 6182 15680 6184 15700
rect 6184 15680 6236 15700
rect 6236 15680 6238 15700
rect 4802 14864 4858 14920
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 6274 14764 6276 14784
rect 6276 14764 6328 14784
rect 6328 14764 6330 14784
rect 6274 14728 6330 14764
rect 5722 14048 5778 14104
rect 6274 14456 6330 14512
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 4434 10512 4490 10568
rect 4618 11328 4674 11384
rect 5262 12180 5264 12200
rect 5264 12180 5316 12200
rect 5316 12180 5318 12200
rect 5262 12144 5318 12180
rect 5078 11636 5080 11656
rect 5080 11636 5132 11656
rect 5132 11636 5134 11656
rect 5078 11600 5134 11636
rect 5354 11464 5410 11520
rect 5354 10784 5410 10840
rect 5446 10648 5502 10704
rect 4802 10412 4804 10432
rect 4804 10412 4856 10432
rect 4856 10412 4858 10432
rect 4802 10376 4858 10412
rect 4894 10104 4950 10160
rect 4986 8492 5042 8528
rect 4986 8472 4988 8492
rect 4988 8472 5040 8492
rect 5040 8472 5042 8492
rect 4986 8084 5042 8120
rect 4986 8064 4988 8084
rect 4988 8064 5040 8084
rect 5040 8064 5042 8084
rect 4710 5616 4766 5672
rect 4802 4528 4858 4584
rect 4618 4120 4674 4176
rect 4342 3440 4398 3496
rect 5354 4528 5410 4584
rect 5722 8336 5778 8392
rect 5630 3984 5686 4040
rect 5170 3712 5226 3768
rect 4250 2624 4306 2680
rect 4066 856 4122 912
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6642 15272 6698 15328
rect 6826 15020 6882 15056
rect 6826 15000 6828 15020
rect 6828 15000 6880 15020
rect 6880 15000 6882 15020
rect 8298 16496 8354 16552
rect 9126 16496 9182 16552
rect 8298 15816 8354 15872
rect 6918 14048 6974 14104
rect 6918 12280 6974 12336
rect 7378 13232 7434 13288
rect 8390 13524 8446 13560
rect 8390 13504 8392 13524
rect 8392 13504 8444 13524
rect 8444 13504 8446 13524
rect 7562 12960 7618 13016
rect 8758 13404 8760 13424
rect 8760 13404 8812 13424
rect 8812 13404 8814 13424
rect 8758 13368 8814 13404
rect 8298 13232 8354 13288
rect 7194 12144 7250 12200
rect 8482 11736 8538 11792
rect 7654 11348 7710 11384
rect 7654 11328 7656 11348
rect 7656 11328 7708 11348
rect 7708 11328 7710 11348
rect 7102 9560 7158 9616
rect 6366 7928 6422 7984
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 7286 8744 7342 8800
rect 7470 5752 7526 5808
rect 7286 4120 7342 4176
rect 5814 2488 5870 2544
rect 7930 11464 7986 11520
rect 7746 11092 7748 11112
rect 7748 11092 7800 11112
rect 7800 11092 7802 11112
rect 7746 11056 7802 11092
rect 7930 11056 7986 11112
rect 8850 12588 8852 12608
rect 8852 12588 8904 12608
rect 8904 12588 8906 12608
rect 8850 12552 8906 12588
rect 7746 5888 7802 5944
rect 8666 10376 8722 10432
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 10690 18672 10746 18728
rect 12714 18708 12716 18728
rect 12716 18708 12768 18728
rect 12768 18708 12770 18728
rect 9954 17076 9956 17096
rect 9956 17076 10008 17096
rect 10008 17076 10010 17096
rect 9954 17040 10010 17076
rect 9218 15000 9274 15056
rect 9770 13912 9826 13968
rect 9862 12844 9918 12880
rect 9862 12824 9864 12844
rect 9864 12824 9916 12844
rect 9916 12824 9918 12844
rect 9034 8336 9090 8392
rect 8850 5636 8906 5672
rect 8850 5616 8852 5636
rect 8852 5616 8904 5636
rect 8904 5616 8906 5636
rect 8298 4936 8354 4992
rect 8574 4664 8630 4720
rect 8298 3576 8354 3632
rect 9126 6196 9128 6216
rect 9128 6196 9180 6216
rect 9180 6196 9182 6216
rect 9126 6160 9182 6196
rect 10046 13388 10102 13424
rect 10046 13368 10048 13388
rect 10048 13368 10100 13388
rect 10100 13368 10102 13388
rect 10138 12708 10194 12744
rect 10138 12688 10140 12708
rect 10140 12688 10192 12708
rect 10192 12688 10194 12708
rect 10414 15272 10470 15328
rect 10506 14068 10562 14104
rect 10506 14048 10508 14068
rect 10508 14048 10560 14068
rect 10560 14048 10562 14068
rect 10598 13812 10600 13832
rect 10600 13812 10652 13832
rect 10652 13812 10654 13832
rect 10322 11192 10378 11248
rect 10598 13776 10654 13812
rect 10138 8200 10194 8256
rect 9954 8064 10010 8120
rect 10414 8780 10416 8800
rect 10416 8780 10468 8800
rect 10468 8780 10470 8800
rect 10414 8744 10470 8780
rect 10506 6976 10562 7032
rect 10138 6704 10194 6760
rect 9586 3984 9642 4040
rect 9402 3848 9458 3904
rect 10414 6296 10470 6352
rect 10322 5908 10378 5944
rect 10322 5888 10324 5908
rect 10324 5888 10376 5908
rect 10376 5888 10378 5908
rect 10322 4528 10378 4584
rect 10230 3712 10286 3768
rect 10138 3440 10194 3496
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 5078 2080 5134 2136
rect 9770 2508 9826 2544
rect 12714 18672 12770 18708
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11702 13504 11758 13560
rect 13910 17312 13966 17368
rect 14186 17584 14242 17640
rect 13082 15544 13138 15600
rect 13082 15272 13138 15328
rect 13082 12824 13138 12880
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10782 11736 10838 11792
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 11334 11192 11390 11248
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 13174 12688 13230 12744
rect 13174 12416 13230 12472
rect 12990 11756 13046 11792
rect 12990 11736 12992 11756
rect 12992 11736 13044 11756
rect 13044 11736 13046 11756
rect 12162 9596 12164 9616
rect 12164 9596 12216 9616
rect 12216 9596 12218 9616
rect 12162 9560 12218 9596
rect 12070 9016 12126 9072
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 11978 8064 12034 8120
rect 12898 8880 12954 8936
rect 13450 13640 13506 13696
rect 13358 12436 13414 12472
rect 13358 12416 13360 12436
rect 13360 12416 13412 12436
rect 13412 12416 13414 12436
rect 13358 11076 13414 11112
rect 14370 16532 14372 16552
rect 14372 16532 14424 16552
rect 14424 16532 14426 16552
rect 14370 16496 14426 16532
rect 14002 15564 14058 15600
rect 14002 15544 14004 15564
rect 14004 15544 14056 15564
rect 14056 15544 14058 15564
rect 14738 18148 14794 18184
rect 14738 18128 14740 18148
rect 14740 18128 14792 18148
rect 14792 18128 14794 18148
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 16578 17176 16634 17232
rect 14646 16940 14648 16960
rect 14648 16940 14700 16960
rect 14700 16940 14702 16960
rect 14646 16904 14702 16940
rect 13358 11056 13360 11076
rect 13360 11056 13412 11076
rect 13412 11056 13414 11076
rect 13266 8336 13322 8392
rect 11794 7928 11850 7984
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 11794 6976 11850 7032
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 11426 4664 11482 4720
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 11610 3984 11666 4040
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 9770 2488 9772 2508
rect 9772 2488 9824 2508
rect 9824 2488 9826 2508
rect 13634 5752 13690 5808
rect 11978 2352 12034 2408
rect 14646 12144 14702 12200
rect 14646 11872 14702 11928
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15198 15952 15254 16008
rect 15474 15952 15530 16008
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 14922 14884 14978 14920
rect 14922 14864 14924 14884
rect 14924 14864 14976 14884
rect 14976 14864 14978 14884
rect 14554 10648 14610 10704
rect 14830 10648 14886 10704
rect 14186 9288 14242 9344
rect 14002 8200 14058 8256
rect 14830 7248 14886 7304
rect 14554 4528 14610 4584
rect 14002 4120 14058 4176
rect 15106 6316 15162 6352
rect 15106 6296 15108 6316
rect 15108 6296 15160 6316
rect 15160 6296 15162 6316
rect 16394 14476 16450 14512
rect 16394 14456 16396 14476
rect 16396 14456 16448 14476
rect 16448 14456 16450 14476
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16210 13932 16266 13968
rect 16210 13912 16212 13932
rect 16212 13912 16264 13932
rect 16264 13912 16266 13932
rect 15842 13232 15898 13288
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 17498 16496 17554 16552
rect 17222 13776 17278 13832
rect 17130 13504 17186 13560
rect 16486 12416 16542 12472
rect 15842 12280 15898 12336
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15750 9560 15806 9616
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 15658 8336 15714 8392
rect 16210 7928 16266 7984
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15382 5072 15438 5128
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 16946 12724 16948 12744
rect 16948 12724 17000 12744
rect 17000 12724 17002 12744
rect 16946 12688 17002 12724
rect 17130 12688 17186 12744
rect 17590 12180 17592 12200
rect 17592 12180 17644 12200
rect 17644 12180 17646 12200
rect 17590 12144 17646 12180
rect 17130 11192 17186 11248
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 19154 19216 19210 19272
rect 18602 19080 18658 19136
rect 18510 17720 18566 17776
rect 18326 12588 18328 12608
rect 18328 12588 18380 12608
rect 18380 12588 18382 12608
rect 18326 12552 18382 12588
rect 18510 10920 18566 10976
rect 18142 9988 18198 10024
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 25502 23024 25558 23080
rect 24858 22344 24914 22400
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 19062 16224 19118 16280
rect 18878 15816 18934 15872
rect 18694 13096 18750 13152
rect 19062 15816 19118 15872
rect 18878 12008 18934 12064
rect 18786 11600 18842 11656
rect 18786 11192 18842 11248
rect 19338 17332 19394 17368
rect 19338 17312 19340 17332
rect 19340 17312 19392 17332
rect 19392 17312 19394 17332
rect 19522 16088 19578 16144
rect 19338 13912 19394 13968
rect 19154 13640 19210 13696
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20258 15408 20314 15464
rect 19614 14864 19670 14920
rect 19614 13776 19670 13832
rect 19430 12688 19486 12744
rect 19062 12008 19118 12064
rect 18602 10104 18658 10160
rect 18142 9968 18144 9988
rect 18144 9968 18196 9988
rect 18196 9968 18198 9988
rect 18418 9424 18474 9480
rect 18602 9016 18658 9072
rect 19706 9324 19708 9344
rect 19708 9324 19760 9344
rect 19760 9324 19762 9344
rect 19706 9288 19762 9324
rect 19798 8200 19854 8256
rect 16578 7384 16634 7440
rect 17222 6740 17224 6760
rect 17224 6740 17276 6760
rect 17276 6740 17278 6760
rect 17222 6704 17278 6740
rect 16854 6568 16910 6624
rect 16762 6180 16818 6216
rect 16762 6160 16764 6180
rect 16764 6160 16816 6180
rect 16816 6160 16818 6180
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20810 15000 20866 15056
rect 20166 14048 20222 14104
rect 20166 12960 20222 13016
rect 20074 8084 20130 8120
rect 20074 8064 20076 8084
rect 20076 8064 20128 8084
rect 20128 8064 20130 8084
rect 19890 7520 19946 7576
rect 16854 5616 16910 5672
rect 16302 2488 16358 2544
rect 19890 5752 19946 5808
rect 20718 12688 20774 12744
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 21270 12688 21326 12744
rect 20810 12552 20866 12608
rect 20718 12008 20774 12064
rect 20534 8472 20590 8528
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 21270 8880 21326 8936
rect 21270 8336 21326 8392
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 21270 7948 21326 7984
rect 21270 7928 21272 7948
rect 21272 7928 21324 7948
rect 21324 7928 21326 7948
rect 23478 18164 23480 18184
rect 23480 18164 23532 18184
rect 23532 18164 23534 18184
rect 23478 18128 23534 18164
rect 21730 13640 21786 13696
rect 21730 13096 21786 13152
rect 21638 12008 21694 12064
rect 20442 6976 20498 7032
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 21178 3984 21234 4040
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 21362 3732 21418 3768
rect 21362 3712 21364 3732
rect 21364 3712 21416 3732
rect 21416 3712 21418 3732
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 21822 8744 21878 8800
rect 21730 4664 21786 4720
rect 23202 17060 23258 17096
rect 23202 17040 23204 17060
rect 23204 17040 23256 17060
rect 23256 17040 23258 17060
rect 23110 16496 23166 16552
rect 23478 16496 23534 16552
rect 23110 16088 23166 16144
rect 22742 15544 22798 15600
rect 22558 14728 22614 14784
rect 22558 14048 22614 14104
rect 23662 17740 23718 17776
rect 23662 17720 23664 17740
rect 23664 17720 23716 17740
rect 23716 17720 23718 17740
rect 25226 21528 25282 21584
rect 25134 20440 25190 20496
rect 24766 17584 24822 17640
rect 24858 17176 24914 17232
rect 23202 12960 23258 13016
rect 22190 10412 22192 10432
rect 22192 10412 22244 10432
rect 22244 10412 22246 10432
rect 22190 10376 22246 10412
rect 23478 12708 23534 12744
rect 23478 12688 23480 12708
rect 23480 12688 23532 12708
rect 23532 12688 23534 12708
rect 23754 9560 23810 9616
rect 23294 8472 23350 8528
rect 23754 8880 23810 8936
rect 24306 15020 24362 15056
rect 24306 15000 24308 15020
rect 24308 15000 24360 15020
rect 24360 15000 24362 15020
rect 23110 7540 23166 7576
rect 23110 7520 23112 7540
rect 23112 7520 23164 7540
rect 23164 7520 23166 7540
rect 23938 8492 23994 8528
rect 23938 8472 23940 8492
rect 23940 8472 23992 8492
rect 23992 8472 23994 8492
rect 24214 8336 24270 8392
rect 22650 6568 22706 6624
rect 23478 5752 23534 5808
rect 25318 21256 25374 21312
rect 25226 18808 25282 18864
rect 25226 15136 25282 15192
rect 25042 12416 25098 12472
rect 25042 11736 25098 11792
rect 24858 10376 24914 10432
rect 24582 6296 24638 6352
rect 25410 20032 25466 20088
rect 25502 18264 25558 18320
rect 25502 17176 25558 17232
rect 25502 16904 25558 16960
rect 25410 15000 25466 15056
rect 25318 12552 25374 12608
rect 25134 8744 25190 8800
rect 25502 14456 25558 14512
rect 25502 12844 25558 12880
rect 25502 12824 25504 12844
rect 25504 12824 25556 12844
rect 25556 12824 25558 12844
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 26238 20304 26294 20360
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25870 18808 25926 18864
rect 25778 14900 25780 14920
rect 25780 14900 25832 14920
rect 25832 14900 25834 14920
rect 25778 14864 25834 14900
rect 25686 14728 25742 14784
rect 25686 14592 25742 14648
rect 25778 14456 25834 14512
rect 25686 13368 25742 13424
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 26514 17040 26570 17096
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 26054 14728 26110 14784
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 26606 16496 26662 16552
rect 26422 14048 26478 14104
rect 26054 13932 26110 13968
rect 26054 13912 26056 13932
rect 26056 13912 26108 13932
rect 26108 13912 26110 13932
rect 26238 13640 26294 13696
rect 26238 13368 26294 13424
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25778 12416 25834 12472
rect 25502 12144 25558 12200
rect 25778 10920 25834 10976
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25870 10376 25926 10432
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26514 12300 26570 12336
rect 26514 12280 26516 12300
rect 26516 12280 26568 12300
rect 26568 12280 26570 12300
rect 26698 14456 26754 14512
rect 26974 14864 27030 14920
rect 27250 14864 27306 14920
rect 26698 12724 26700 12744
rect 26700 12724 26752 12744
rect 26752 12724 26754 12744
rect 26698 12688 26754 12724
rect 26790 12144 26846 12200
rect 26698 11600 26754 11656
rect 26514 11212 26570 11248
rect 26514 11192 26516 11212
rect 26516 11192 26568 11212
rect 26568 11192 26570 11212
rect 26606 11056 26662 11112
rect 26698 9832 26754 9888
rect 26514 9036 26570 9072
rect 25410 8472 25466 8528
rect 24950 6840 25006 6896
rect 23754 3032 23810 3088
rect 24306 2508 24362 2544
rect 24306 2488 24308 2508
rect 24308 2488 24360 2508
rect 24360 2488 24362 2508
rect 26514 9016 26516 9036
rect 26516 9016 26568 9036
rect 26568 9016 26570 9036
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26698 8608 26754 8664
rect 26330 8336 26386 8392
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26606 8064 26662 8120
rect 26514 7948 26570 7984
rect 26514 7928 26516 7948
rect 26516 7928 26568 7948
rect 26568 7928 26570 7948
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26698 6840 26754 6896
rect 26606 6332 26608 6352
rect 26608 6332 26660 6352
rect 26660 6332 26662 6352
rect 26606 6296 26662 6332
rect 26422 6160 26478 6216
rect 26974 10648 27030 10704
rect 26882 9968 26938 10024
rect 26698 5636 26754 5672
rect 26698 5616 26700 5636
rect 26700 5616 26752 5636
rect 26752 5616 26754 5636
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25870 5208 25926 5264
rect 26422 5108 26424 5128
rect 26424 5108 26476 5128
rect 26476 5108 26478 5128
rect 26422 5072 26478 5108
rect 26514 4684 26570 4720
rect 26514 4664 26516 4684
rect 26516 4664 26568 4684
rect 26568 4664 26570 4684
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26606 4392 26662 4448
rect 26698 4120 26754 4176
rect 26514 3984 26570 4040
rect 26422 3576 26478 3632
rect 25502 3460 25558 3496
rect 25502 3440 25504 3460
rect 25504 3440 25556 3460
rect 25556 3440 25558 3460
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 856 25926 912
rect 3974 312 4030 368
rect 27526 10648 27582 10704
rect 27618 9324 27620 9344
rect 27620 9324 27672 9344
rect 27672 9324 27674 9344
rect 27618 9288 27674 9324
rect 27526 7384 27582 7440
rect 27250 3712 27306 3768
rect 27526 3032 27582 3088
rect 27710 7420 27712 7440
rect 27712 7420 27764 7440
rect 27764 7420 27766 7440
rect 27710 7384 27766 7420
rect 26790 2760 26846 2816
rect 26698 1400 26754 1456
rect 27802 2080 27858 2136
rect 26606 312 26662 368
<< metal3 >>
rect 0 23626 480 23656
rect 3325 23626 3391 23629
rect 0 23624 3391 23626
rect 0 23568 3330 23624
rect 3386 23568 3391 23624
rect 0 23566 3391 23568
rect 0 23536 480 23566
rect 3325 23563 3391 23566
rect 25589 23626 25655 23629
rect 29520 23626 30000 23656
rect 25589 23624 30000 23626
rect 25589 23568 25594 23624
rect 25650 23568 30000 23624
rect 25589 23566 30000 23568
rect 25589 23563 25655 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3417 23082 3483 23085
rect 0 23080 3483 23082
rect 0 23024 3422 23080
rect 3478 23024 3483 23080
rect 0 23022 3483 23024
rect 0 22992 480 23022
rect 3417 23019 3483 23022
rect 25497 23082 25563 23085
rect 29520 23082 30000 23112
rect 25497 23080 30000 23082
rect 25497 23024 25502 23080
rect 25558 23024 30000 23080
rect 25497 23022 30000 23024
rect 25497 23019 25563 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2405 22402 2471 22405
rect 0 22400 2471 22402
rect 0 22344 2410 22400
rect 2466 22344 2471 22400
rect 0 22342 2471 22344
rect 0 22312 480 22342
rect 2405 22339 2471 22342
rect 24853 22402 24919 22405
rect 29520 22402 30000 22432
rect 24853 22400 30000 22402
rect 24853 22344 24858 22400
rect 24914 22344 30000 22400
rect 24853 22342 30000 22344
rect 24853 22339 24919 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3049 21858 3115 21861
rect 29520 21858 30000 21888
rect 0 21856 3115 21858
rect 0 21800 3054 21856
rect 3110 21800 3115 21856
rect 0 21798 3115 21800
rect 0 21768 480 21798
rect 3049 21795 3115 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 25221 21586 25287 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 25221 21584 26434 21586
rect 25221 21528 25226 21584
rect 25282 21528 26434 21584
rect 25221 21526 26434 21528
rect 25221 21523 25287 21526
rect 0 21314 480 21344
rect 2865 21314 2931 21317
rect 0 21312 2931 21314
rect 0 21256 2870 21312
rect 2926 21256 2931 21312
rect 0 21254 2931 21256
rect 0 21224 480 21254
rect 2865 21251 2931 21254
rect 25313 21314 25379 21317
rect 29520 21314 30000 21344
rect 25313 21312 30000 21314
rect 25313 21256 25318 21312
rect 25374 21256 30000 21312
rect 25313 21254 30000 21256
rect 25313 21251 25379 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3877 20634 3943 20637
rect 29520 20634 30000 20664
rect 0 20632 3943 20634
rect 0 20576 3882 20632
rect 3938 20576 3943 20632
rect 0 20574 3943 20576
rect 0 20544 480 20574
rect 3877 20571 3943 20574
rect 26374 20574 30000 20634
rect 25129 20498 25195 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25129 20496 26434 20498
rect 25129 20440 25134 20496
rect 25190 20440 26434 20496
rect 25129 20438 26434 20440
rect 25129 20435 25195 20438
rect 7465 20362 7531 20365
rect 26233 20362 26299 20365
rect 7465 20360 26299 20362
rect 7465 20304 7470 20360
rect 7526 20304 26238 20360
rect 26294 20304 26299 20360
rect 7465 20302 26299 20304
rect 7465 20299 7531 20302
rect 26233 20299 26299 20302
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 2865 20090 2931 20093
rect 0 20088 2931 20090
rect 0 20032 2870 20088
rect 2926 20032 2931 20088
rect 0 20030 2931 20032
rect 0 20000 480 20030
rect 2865 20027 2931 20030
rect 25405 20090 25471 20093
rect 29520 20090 30000 20120
rect 25405 20088 30000 20090
rect 25405 20032 25410 20088
rect 25466 20032 30000 20088
rect 25405 20030 30000 20032
rect 25405 20027 25471 20030
rect 29520 20000 30000 20030
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19410 480 19440
rect 3141 19410 3207 19413
rect 29520 19410 30000 19440
rect 0 19408 3207 19410
rect 0 19352 3146 19408
rect 3202 19352 3207 19408
rect 0 19350 3207 19352
rect 0 19320 480 19350
rect 3141 19347 3207 19350
rect 25822 19350 30000 19410
rect 19149 19274 19215 19277
rect 25822 19274 25882 19350
rect 29520 19320 30000 19350
rect 19149 19272 25882 19274
rect 19149 19216 19154 19272
rect 19210 19216 25882 19272
rect 19149 19214 25882 19216
rect 19149 19211 19215 19214
rect 18597 19140 18663 19141
rect 18597 19138 18644 19140
rect 18552 19136 18644 19138
rect 18552 19080 18602 19136
rect 18552 19078 18644 19080
rect 18597 19076 18644 19078
rect 18708 19076 18714 19140
rect 18597 19075 18663 19076
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 3969 18866 4035 18869
rect 0 18864 4035 18866
rect 0 18808 3974 18864
rect 4030 18808 4035 18864
rect 0 18806 4035 18808
rect 0 18776 480 18806
rect 3969 18803 4035 18806
rect 18638 18804 18644 18868
rect 18708 18866 18714 18868
rect 25221 18866 25287 18869
rect 18708 18864 25287 18866
rect 18708 18808 25226 18864
rect 25282 18808 25287 18864
rect 18708 18806 25287 18808
rect 18708 18804 18714 18806
rect 25221 18803 25287 18806
rect 25865 18866 25931 18869
rect 29520 18866 30000 18896
rect 25865 18864 30000 18866
rect 25865 18808 25870 18864
rect 25926 18808 30000 18864
rect 25865 18806 30000 18808
rect 25865 18803 25931 18806
rect 29520 18776 30000 18806
rect 10685 18730 10751 18733
rect 12709 18730 12775 18733
rect 10685 18728 12775 18730
rect 10685 18672 10690 18728
rect 10746 18672 12714 18728
rect 12770 18672 12775 18728
rect 10685 18670 12775 18672
rect 10685 18667 10751 18670
rect 12709 18667 12775 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 3509 18322 3575 18325
rect 0 18320 3575 18322
rect 0 18264 3514 18320
rect 3570 18264 3575 18320
rect 0 18262 3575 18264
rect 0 18232 480 18262
rect 3509 18259 3575 18262
rect 25497 18322 25563 18325
rect 29520 18322 30000 18352
rect 25497 18320 30000 18322
rect 25497 18264 25502 18320
rect 25558 18264 30000 18320
rect 25497 18262 30000 18264
rect 25497 18259 25563 18262
rect 29520 18232 30000 18262
rect 14733 18186 14799 18189
rect 23473 18186 23539 18189
rect 14733 18184 23539 18186
rect 14733 18128 14738 18184
rect 14794 18128 23478 18184
rect 23534 18128 23539 18184
rect 14733 18126 23539 18128
rect 14733 18123 14799 18126
rect 23473 18123 23539 18126
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 2681 17914 2747 17917
rect 2681 17912 7666 17914
rect 2681 17856 2686 17912
rect 2742 17856 7666 17912
rect 2681 17854 7666 17856
rect 2681 17851 2747 17854
rect 2313 17778 2379 17781
rect 7465 17778 7531 17781
rect 2313 17776 7531 17778
rect 2313 17720 2318 17776
rect 2374 17720 7470 17776
rect 7526 17720 7531 17776
rect 2313 17718 7531 17720
rect 7606 17778 7666 17854
rect 18505 17778 18571 17781
rect 23657 17778 23723 17781
rect 7606 17776 23723 17778
rect 7606 17720 18510 17776
rect 18566 17720 23662 17776
rect 23718 17720 23723 17776
rect 7606 17718 23723 17720
rect 2313 17715 2379 17718
rect 7465 17715 7531 17718
rect 18505 17715 18571 17718
rect 23657 17715 23723 17718
rect 0 17642 480 17672
rect 4061 17642 4127 17645
rect 14181 17642 14247 17645
rect 0 17640 4127 17642
rect 0 17584 4066 17640
rect 4122 17584 4127 17640
rect 0 17582 4127 17584
rect 0 17552 480 17582
rect 4061 17579 4127 17582
rect 5766 17640 14247 17642
rect 5766 17584 14186 17640
rect 14242 17584 14247 17640
rect 5766 17582 14247 17584
rect 2405 17506 2471 17509
rect 5766 17506 5826 17582
rect 14181 17579 14247 17582
rect 24761 17642 24827 17645
rect 29520 17642 30000 17672
rect 24761 17640 30000 17642
rect 24761 17584 24766 17640
rect 24822 17584 30000 17640
rect 24761 17582 30000 17584
rect 24761 17579 24827 17582
rect 29520 17552 30000 17582
rect 2405 17504 5826 17506
rect 2405 17448 2410 17504
rect 2466 17448 5826 17504
rect 2405 17446 5826 17448
rect 2405 17443 2471 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 7465 17370 7531 17373
rect 13905 17370 13971 17373
rect 19333 17370 19399 17373
rect 7465 17368 13971 17370
rect 7465 17312 7470 17368
rect 7526 17312 13910 17368
rect 13966 17312 13971 17368
rect 7465 17310 13971 17312
rect 7465 17307 7531 17310
rect 13905 17307 13971 17310
rect 16990 17368 19399 17370
rect 16990 17312 19338 17368
rect 19394 17312 19399 17368
rect 16990 17310 19399 17312
rect 3141 17234 3207 17237
rect 16573 17234 16639 17237
rect 16990 17234 17050 17310
rect 19333 17307 19399 17310
rect 24853 17234 24919 17237
rect 25497 17234 25563 17237
rect 3141 17232 17050 17234
rect 3141 17176 3146 17232
rect 3202 17176 16578 17232
rect 16634 17176 17050 17232
rect 3141 17174 17050 17176
rect 17174 17232 25563 17234
rect 17174 17176 24858 17232
rect 24914 17176 25502 17232
rect 25558 17176 25563 17232
rect 17174 17174 25563 17176
rect 3141 17171 3207 17174
rect 16573 17171 16639 17174
rect 0 17098 480 17128
rect 3785 17098 3851 17101
rect 0 17096 3851 17098
rect 0 17040 3790 17096
rect 3846 17040 3851 17096
rect 0 17038 3851 17040
rect 0 17008 480 17038
rect 3785 17035 3851 17038
rect 9949 17098 10015 17101
rect 17174 17098 17234 17174
rect 24853 17171 24919 17174
rect 25497 17171 25563 17174
rect 23197 17098 23263 17101
rect 26509 17098 26575 17101
rect 29520 17098 30000 17128
rect 9949 17096 17234 17098
rect 9949 17040 9954 17096
rect 10010 17040 17234 17096
rect 9949 17038 17234 17040
rect 17358 17096 26575 17098
rect 17358 17040 23202 17096
rect 23258 17040 26514 17096
rect 26570 17040 26575 17096
rect 17358 17038 26575 17040
rect 9949 17035 10015 17038
rect 14641 16962 14707 16965
rect 17358 16962 17418 17038
rect 23197 17035 23263 17038
rect 26509 17035 26575 17038
rect 26742 17038 30000 17098
rect 14641 16960 17418 16962
rect 14641 16904 14646 16960
rect 14702 16904 17418 16960
rect 14641 16902 17418 16904
rect 25497 16962 25563 16965
rect 26742 16962 26802 17038
rect 29520 17008 30000 17038
rect 25497 16960 26802 16962
rect 25497 16904 25502 16960
rect 25558 16904 26802 16960
rect 25497 16902 26802 16904
rect 14641 16899 14707 16902
rect 25497 16899 25563 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 8293 16554 8359 16557
rect 9121 16554 9187 16557
rect 14365 16554 14431 16557
rect 17493 16554 17559 16557
rect 8293 16552 14290 16554
rect 8293 16496 8298 16552
rect 8354 16496 9126 16552
rect 9182 16496 14290 16552
rect 8293 16494 14290 16496
rect 8293 16491 8359 16494
rect 9121 16491 9187 16494
rect 0 16418 480 16448
rect 4705 16418 4771 16421
rect 0 16416 4771 16418
rect 0 16360 4710 16416
rect 4766 16360 4771 16416
rect 0 16358 4771 16360
rect 0 16328 480 16358
rect 4705 16355 4771 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 14230 16146 14290 16494
rect 14365 16552 17559 16554
rect 14365 16496 14370 16552
rect 14426 16496 17498 16552
rect 17554 16496 17559 16552
rect 14365 16494 17559 16496
rect 14365 16491 14431 16494
rect 17493 16491 17559 16494
rect 23105 16554 23171 16557
rect 23473 16554 23539 16557
rect 26601 16554 26667 16557
rect 23105 16552 26667 16554
rect 23105 16496 23110 16552
rect 23166 16496 23478 16552
rect 23534 16496 26606 16552
rect 26662 16496 26667 16552
rect 23105 16494 26667 16496
rect 23105 16491 23171 16494
rect 23473 16491 23539 16494
rect 26601 16491 26667 16494
rect 29520 16418 30000 16448
rect 26374 16358 30000 16418
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 19057 16282 19123 16285
rect 19057 16280 19810 16282
rect 19057 16224 19062 16280
rect 19118 16224 19810 16280
rect 19057 16222 19810 16224
rect 19057 16219 19123 16222
rect 19517 16146 19583 16149
rect 14230 16144 19583 16146
rect 14230 16088 19522 16144
rect 19578 16088 19583 16144
rect 14230 16086 19583 16088
rect 19750 16146 19810 16222
rect 23105 16146 23171 16149
rect 19750 16144 23171 16146
rect 19750 16088 23110 16144
rect 23166 16088 23171 16144
rect 19750 16086 23171 16088
rect 19517 16083 19583 16086
rect 23105 16083 23171 16086
rect 3969 16010 4035 16013
rect 15193 16010 15259 16013
rect 3969 16008 15259 16010
rect 3969 15952 3974 16008
rect 4030 15952 15198 16008
rect 15254 15952 15259 16008
rect 3969 15950 15259 15952
rect 3969 15947 4035 15950
rect 15193 15947 15259 15950
rect 15469 16010 15535 16013
rect 26374 16010 26434 16358
rect 29520 16328 30000 16358
rect 15469 16008 26434 16010
rect 15469 15952 15474 16008
rect 15530 15952 26434 16008
rect 15469 15950 26434 15952
rect 15469 15947 15535 15950
rect 0 15874 480 15904
rect 8293 15874 8359 15877
rect 18873 15874 18939 15877
rect 19057 15874 19123 15877
rect 29520 15874 30000 15904
rect 0 15872 8359 15874
rect 0 15816 8298 15872
rect 8354 15816 8359 15872
rect 0 15814 8359 15816
rect 0 15784 480 15814
rect 8293 15811 8359 15814
rect 11470 15872 19123 15874
rect 11470 15816 18878 15872
rect 18934 15816 19062 15872
rect 19118 15816 19123 15872
rect 11470 15814 19123 15816
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 3877 15738 3943 15741
rect 5717 15738 5783 15741
rect 6177 15738 6243 15741
rect 3877 15736 6243 15738
rect 3877 15680 3882 15736
rect 3938 15680 5722 15736
rect 5778 15680 6182 15736
rect 6238 15680 6243 15736
rect 3877 15678 6243 15680
rect 3877 15675 3943 15678
rect 5717 15675 5783 15678
rect 6177 15675 6243 15678
rect 4429 15602 4495 15605
rect 11470 15602 11530 15814
rect 18873 15811 18939 15814
rect 19057 15811 19123 15814
rect 25822 15814 30000 15874
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 15743 21264 15744
rect 4429 15600 11530 15602
rect 4429 15544 4434 15600
rect 4490 15544 11530 15600
rect 4429 15542 11530 15544
rect 13077 15602 13143 15605
rect 13997 15602 14063 15605
rect 22737 15602 22803 15605
rect 13077 15600 22803 15602
rect 13077 15544 13082 15600
rect 13138 15544 14002 15600
rect 14058 15544 22742 15600
rect 22798 15544 22803 15600
rect 13077 15542 22803 15544
rect 4429 15539 4495 15542
rect 13077 15539 13143 15542
rect 13997 15539 14063 15542
rect 22737 15539 22803 15542
rect 4521 15466 4587 15469
rect 20253 15466 20319 15469
rect 25822 15466 25882 15814
rect 29520 15784 30000 15814
rect 4521 15464 10610 15466
rect 4521 15408 4526 15464
rect 4582 15408 10610 15464
rect 4521 15406 10610 15408
rect 4521 15403 4587 15406
rect 0 15330 480 15360
rect 3877 15330 3943 15333
rect 0 15328 3943 15330
rect 0 15272 3882 15328
rect 3938 15272 3943 15328
rect 0 15270 3943 15272
rect 0 15240 480 15270
rect 3877 15267 3943 15270
rect 6637 15330 6703 15333
rect 10409 15330 10475 15333
rect 6637 15328 10475 15330
rect 6637 15272 6642 15328
rect 6698 15272 10414 15328
rect 10470 15272 10475 15328
rect 6637 15270 10475 15272
rect 10550 15330 10610 15406
rect 20253 15464 25882 15466
rect 20253 15408 20258 15464
rect 20314 15408 25882 15464
rect 20253 15406 25882 15408
rect 20253 15403 20319 15406
rect 13077 15330 13143 15333
rect 29520 15330 30000 15360
rect 10550 15328 13143 15330
rect 10550 15272 13082 15328
rect 13138 15272 13143 15328
rect 10550 15270 13143 15272
rect 6637 15267 6703 15270
rect 10409 15267 10475 15270
rect 13077 15267 13143 15270
rect 26374 15270 30000 15330
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 15199 26264 15200
rect 25078 15132 25084 15196
rect 25148 15194 25154 15196
rect 25221 15194 25287 15197
rect 25148 15192 25287 15194
rect 25148 15136 25226 15192
rect 25282 15136 25287 15192
rect 25148 15134 25287 15136
rect 25148 15132 25154 15134
rect 25221 15131 25287 15134
rect 6821 15058 6887 15061
rect 9213 15058 9279 15061
rect 6821 15056 9279 15058
rect 6821 15000 6826 15056
rect 6882 15000 9218 15056
rect 9274 15000 9279 15056
rect 6821 14998 9279 15000
rect 6821 14995 6887 14998
rect 9213 14995 9279 14998
rect 20805 15058 20871 15061
rect 24301 15058 24367 15061
rect 20805 15056 24367 15058
rect 20805 15000 20810 15056
rect 20866 15000 24306 15056
rect 24362 15000 24367 15056
rect 20805 14998 24367 15000
rect 20805 14995 20871 14998
rect 24301 14995 24367 14998
rect 25405 15058 25471 15061
rect 26374 15058 26434 15270
rect 29520 15240 30000 15270
rect 25405 15056 26434 15058
rect 25405 15000 25410 15056
rect 25466 15000 26434 15056
rect 25405 14998 26434 15000
rect 25405 14995 25471 14998
rect 4797 14922 4863 14925
rect 14917 14922 14983 14925
rect 4797 14920 14983 14922
rect 4797 14864 4802 14920
rect 4858 14864 14922 14920
rect 14978 14864 14983 14920
rect 4797 14862 14983 14864
rect 4797 14859 4863 14862
rect 14917 14859 14983 14862
rect 19609 14922 19675 14925
rect 25773 14922 25839 14925
rect 26969 14922 27035 14925
rect 27245 14922 27311 14925
rect 19609 14920 27311 14922
rect 19609 14864 19614 14920
rect 19670 14864 25778 14920
rect 25834 14864 26974 14920
rect 27030 14864 27250 14920
rect 27306 14864 27311 14920
rect 19609 14862 27311 14864
rect 19609 14859 19675 14862
rect 25773 14859 25839 14862
rect 26969 14859 27035 14862
rect 27245 14859 27311 14862
rect 1945 14786 2011 14789
rect 6269 14786 6335 14789
rect 1945 14784 6335 14786
rect 1945 14728 1950 14784
rect 2006 14728 6274 14784
rect 6330 14728 6335 14784
rect 1945 14726 6335 14728
rect 1945 14723 2011 14726
rect 6269 14723 6335 14726
rect 22553 14786 22619 14789
rect 25681 14786 25747 14789
rect 26049 14786 26115 14789
rect 22553 14784 26115 14786
rect 22553 14728 22558 14784
rect 22614 14728 25686 14784
rect 25742 14728 26054 14784
rect 26110 14728 26115 14784
rect 22553 14726 26115 14728
rect 22553 14723 22619 14726
rect 25681 14723 25747 14726
rect 26049 14723 26115 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 4061 14650 4127 14653
rect 0 14648 4127 14650
rect 0 14592 4066 14648
rect 4122 14592 4127 14648
rect 0 14590 4127 14592
rect 0 14560 480 14590
rect 4061 14587 4127 14590
rect 25681 14650 25747 14653
rect 29520 14650 30000 14680
rect 25681 14648 30000 14650
rect 25681 14592 25686 14648
rect 25742 14592 30000 14648
rect 25681 14590 30000 14592
rect 25681 14587 25747 14590
rect 29520 14560 30000 14590
rect 6269 14514 6335 14517
rect 16389 14514 16455 14517
rect 25497 14514 25563 14517
rect 6269 14512 25563 14514
rect 6269 14456 6274 14512
rect 6330 14456 16394 14512
rect 16450 14456 25502 14512
rect 25558 14456 25563 14512
rect 6269 14454 25563 14456
rect 6269 14451 6335 14454
rect 16389 14451 16455 14454
rect 25497 14451 25563 14454
rect 25773 14514 25839 14517
rect 26693 14514 26759 14517
rect 25773 14512 26759 14514
rect 25773 14456 25778 14512
rect 25834 14456 26698 14512
rect 26754 14456 26759 14512
rect 25773 14454 26759 14456
rect 25773 14451 25839 14454
rect 26693 14451 26759 14454
rect 3049 14242 3115 14245
rect 3601 14242 3667 14245
rect 1350 14240 3667 14242
rect 1350 14184 3054 14240
rect 3110 14184 3606 14240
rect 3662 14184 3667 14240
rect 1350 14182 3667 14184
rect 0 14106 480 14136
rect 1350 14106 1410 14182
rect 3049 14179 3115 14182
rect 3601 14179 3667 14182
rect 5944 14176 6264 14177
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 0 14046 1410 14106
rect 1485 14106 1551 14109
rect 4429 14106 4495 14109
rect 5717 14106 5783 14109
rect 1485 14104 5783 14106
rect 1485 14048 1490 14104
rect 1546 14048 4434 14104
rect 4490 14048 5722 14104
rect 5778 14048 5783 14104
rect 1485 14046 5783 14048
rect 0 14016 480 14046
rect 1485 14043 1551 14046
rect 4429 14043 4495 14046
rect 5717 14043 5783 14046
rect 6913 14106 6979 14109
rect 10501 14106 10567 14109
rect 6913 14104 10567 14106
rect 6913 14048 6918 14104
rect 6974 14048 10506 14104
rect 10562 14048 10567 14104
rect 6913 14046 10567 14048
rect 6913 14043 6979 14046
rect 10501 14043 10567 14046
rect 20161 14106 20227 14109
rect 22553 14106 22619 14109
rect 20161 14104 22619 14106
rect 20161 14048 20166 14104
rect 20222 14048 22558 14104
rect 22614 14048 22619 14104
rect 20161 14046 22619 14048
rect 20161 14043 20227 14046
rect 22553 14043 22619 14046
rect 26417 14106 26483 14109
rect 29520 14106 30000 14136
rect 26417 14104 30000 14106
rect 26417 14048 26422 14104
rect 26478 14048 30000 14104
rect 26417 14046 30000 14048
rect 26417 14043 26483 14046
rect 29520 14016 30000 14046
rect 3049 13970 3115 13973
rect 3509 13970 3575 13973
rect 9765 13972 9831 13973
rect 9765 13970 9812 13972
rect 3049 13968 9812 13970
rect 3049 13912 3054 13968
rect 3110 13912 3514 13968
rect 3570 13912 9770 13968
rect 3049 13910 9812 13912
rect 3049 13907 3115 13910
rect 3509 13907 3575 13910
rect 9765 13908 9812 13910
rect 9876 13908 9882 13972
rect 16205 13970 16271 13973
rect 19333 13970 19399 13973
rect 16205 13968 19399 13970
rect 16205 13912 16210 13968
rect 16266 13912 19338 13968
rect 19394 13912 19399 13968
rect 16205 13910 19399 13912
rect 9765 13907 9831 13908
rect 16205 13907 16271 13910
rect 19333 13907 19399 13910
rect 25630 13908 25636 13972
rect 25700 13970 25706 13972
rect 26049 13970 26115 13973
rect 25700 13968 26115 13970
rect 25700 13912 26054 13968
rect 26110 13912 26115 13968
rect 25700 13910 26115 13912
rect 25700 13908 25706 13910
rect 26049 13907 26115 13910
rect 10593 13834 10659 13837
rect 17217 13834 17283 13837
rect 19609 13834 19675 13837
rect 10593 13832 19675 13834
rect 10593 13776 10598 13832
rect 10654 13776 17222 13832
rect 17278 13776 19614 13832
rect 19670 13776 19675 13832
rect 10593 13774 19675 13776
rect 10593 13771 10659 13774
rect 17217 13771 17283 13774
rect 19609 13771 19675 13774
rect 13445 13698 13511 13701
rect 19149 13698 19215 13701
rect 13445 13696 19215 13698
rect 13445 13640 13450 13696
rect 13506 13640 19154 13696
rect 19210 13640 19215 13696
rect 13445 13638 19215 13640
rect 13445 13635 13511 13638
rect 19149 13635 19215 13638
rect 21725 13698 21791 13701
rect 26233 13698 26299 13701
rect 21725 13696 26299 13698
rect 21725 13640 21730 13696
rect 21786 13640 26238 13696
rect 26294 13640 26299 13696
rect 21725 13638 26299 13640
rect 21725 13635 21791 13638
rect 26233 13635 26299 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 3785 13562 3851 13565
rect 8385 13562 8451 13565
rect 3785 13560 8451 13562
rect 3785 13504 3790 13560
rect 3846 13504 8390 13560
rect 8446 13504 8451 13560
rect 3785 13502 8451 13504
rect 3785 13499 3851 13502
rect 8385 13499 8451 13502
rect 11697 13562 11763 13565
rect 17125 13562 17191 13565
rect 11697 13560 17191 13562
rect 11697 13504 11702 13560
rect 11758 13504 17130 13560
rect 17186 13504 17191 13560
rect 11697 13502 17191 13504
rect 11697 13499 11763 13502
rect 17125 13499 17191 13502
rect 0 13426 480 13456
rect 2957 13426 3023 13429
rect 0 13424 3023 13426
rect 0 13368 2962 13424
rect 3018 13368 3023 13424
rect 0 13366 3023 13368
rect 0 13336 480 13366
rect 2957 13363 3023 13366
rect 4061 13426 4127 13429
rect 8753 13426 8819 13429
rect 4061 13424 8819 13426
rect 4061 13368 4066 13424
rect 4122 13368 8758 13424
rect 8814 13368 8819 13424
rect 4061 13366 8819 13368
rect 4061 13363 4127 13366
rect 8753 13363 8819 13366
rect 10041 13426 10107 13429
rect 25681 13426 25747 13429
rect 10041 13424 25747 13426
rect 10041 13368 10046 13424
rect 10102 13368 25686 13424
rect 25742 13368 25747 13424
rect 10041 13366 25747 13368
rect 10041 13363 10107 13366
rect 25681 13363 25747 13366
rect 26233 13426 26299 13429
rect 29520 13426 30000 13456
rect 26233 13424 30000 13426
rect 26233 13368 26238 13424
rect 26294 13368 30000 13424
rect 26233 13366 30000 13368
rect 26233 13363 26299 13366
rect 29520 13336 30000 13366
rect 3233 13290 3299 13293
rect 7373 13290 7439 13293
rect 3233 13288 7439 13290
rect 3233 13232 3238 13288
rect 3294 13232 7378 13288
rect 7434 13232 7439 13288
rect 3233 13230 7439 13232
rect 3233 13227 3299 13230
rect 7373 13227 7439 13230
rect 8293 13290 8359 13293
rect 15837 13290 15903 13293
rect 8293 13288 15903 13290
rect 8293 13232 8298 13288
rect 8354 13232 15842 13288
rect 15898 13232 15903 13288
rect 8293 13230 15903 13232
rect 8293 13227 8359 13230
rect 15837 13227 15903 13230
rect 18689 13154 18755 13157
rect 21725 13154 21791 13157
rect 18689 13152 21791 13154
rect 18689 13096 18694 13152
rect 18750 13096 21730 13152
rect 21786 13096 21791 13152
rect 18689 13094 21791 13096
rect 18689 13091 18755 13094
rect 21725 13091 21791 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 7557 13018 7623 13021
rect 20161 13018 20227 13021
rect 23197 13018 23263 13021
rect 6502 13016 9874 13018
rect 6502 12960 7562 13016
rect 7618 12960 9874 13016
rect 6502 12958 9874 12960
rect 0 12882 480 12912
rect 2773 12882 2839 12885
rect 0 12880 2839 12882
rect 0 12824 2778 12880
rect 2834 12824 2839 12880
rect 0 12822 2839 12824
rect 0 12792 480 12822
rect 2773 12819 2839 12822
rect 2957 12882 3023 12885
rect 6502 12882 6562 12958
rect 7557 12955 7623 12958
rect 2957 12880 6562 12882
rect 2957 12824 2962 12880
rect 3018 12824 6562 12880
rect 2957 12822 6562 12824
rect 9814 12885 9874 12958
rect 20161 13016 25698 13018
rect 20161 12960 20166 13016
rect 20222 12960 23202 13016
rect 23258 12960 25698 13016
rect 20161 12958 25698 12960
rect 20161 12955 20227 12958
rect 23197 12955 23263 12958
rect 9814 12882 9923 12885
rect 13077 12882 13143 12885
rect 25497 12882 25563 12885
rect 9814 12880 11714 12882
rect 9814 12824 9862 12880
rect 9918 12824 11714 12880
rect 9814 12822 11714 12824
rect 2957 12819 3023 12822
rect 9857 12819 9923 12822
rect 10133 12746 10199 12749
rect 10133 12744 11530 12746
rect 10133 12688 10138 12744
rect 10194 12688 11530 12744
rect 10133 12686 11530 12688
rect 10133 12683 10199 12686
rect 3785 12610 3851 12613
rect 8845 12610 8911 12613
rect 3785 12608 8911 12610
rect 3785 12552 3790 12608
rect 3846 12552 8850 12608
rect 8906 12552 8911 12608
rect 3785 12550 8911 12552
rect 3785 12547 3851 12550
rect 8845 12547 8911 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 11470 12474 11530 12686
rect 11654 12610 11714 12822
rect 13077 12880 25563 12882
rect 13077 12824 13082 12880
rect 13138 12824 25502 12880
rect 25558 12824 25563 12880
rect 13077 12822 25563 12824
rect 25638 12882 25698 12958
rect 29520 12882 30000 12912
rect 25638 12822 30000 12882
rect 13077 12819 13143 12822
rect 25497 12819 25563 12822
rect 29520 12792 30000 12822
rect 13169 12746 13235 12749
rect 16941 12746 17007 12749
rect 13169 12744 17007 12746
rect 13169 12688 13174 12744
rect 13230 12688 16946 12744
rect 17002 12688 17007 12744
rect 13169 12686 17007 12688
rect 13169 12683 13235 12686
rect 16941 12683 17007 12686
rect 17125 12746 17191 12749
rect 19425 12746 19491 12749
rect 20713 12746 20779 12749
rect 17125 12744 20779 12746
rect 17125 12688 17130 12744
rect 17186 12688 19430 12744
rect 19486 12688 20718 12744
rect 20774 12688 20779 12744
rect 17125 12686 20779 12688
rect 17125 12683 17191 12686
rect 19425 12683 19491 12686
rect 20713 12683 20779 12686
rect 21265 12746 21331 12749
rect 23473 12746 23539 12749
rect 21265 12744 23539 12746
rect 21265 12688 21270 12744
rect 21326 12688 23478 12744
rect 23534 12688 23539 12744
rect 21265 12686 23539 12688
rect 21265 12683 21331 12686
rect 23473 12683 23539 12686
rect 25078 12684 25084 12748
rect 25148 12746 25154 12748
rect 26693 12746 26759 12749
rect 25148 12744 26759 12746
rect 25148 12688 26698 12744
rect 26754 12688 26759 12744
rect 25148 12686 26759 12688
rect 25148 12684 25154 12686
rect 26693 12683 26759 12686
rect 18321 12610 18387 12613
rect 20805 12610 20871 12613
rect 11654 12608 20871 12610
rect 11654 12552 18326 12608
rect 18382 12552 20810 12608
rect 20866 12552 20871 12608
rect 11654 12550 20871 12552
rect 18321 12547 18387 12550
rect 20805 12547 20871 12550
rect 25313 12610 25379 12613
rect 25313 12608 25514 12610
rect 25313 12552 25318 12608
rect 25374 12552 25514 12608
rect 25313 12550 25514 12552
rect 25313 12547 25379 12550
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 13169 12474 13235 12477
rect 11470 12472 13235 12474
rect 11470 12416 13174 12472
rect 13230 12416 13235 12472
rect 11470 12414 13235 12416
rect 13169 12411 13235 12414
rect 13353 12474 13419 12477
rect 16481 12474 16547 12477
rect 25037 12476 25103 12477
rect 25037 12474 25084 12476
rect 13353 12472 16547 12474
rect 13353 12416 13358 12472
rect 13414 12416 16486 12472
rect 16542 12416 16547 12472
rect 13353 12414 16547 12416
rect 24992 12472 25084 12474
rect 24992 12416 25042 12472
rect 24992 12414 25084 12416
rect 13353 12411 13419 12414
rect 16481 12411 16547 12414
rect 25037 12412 25084 12414
rect 25148 12412 25154 12476
rect 25454 12474 25514 12550
rect 25773 12474 25839 12477
rect 25454 12472 25839 12474
rect 25454 12416 25778 12472
rect 25834 12416 25839 12472
rect 25454 12414 25839 12416
rect 25037 12411 25103 12412
rect 25773 12411 25839 12414
rect 0 12338 480 12368
rect 6913 12338 6979 12341
rect 0 12336 6979 12338
rect 0 12280 6918 12336
rect 6974 12280 6979 12336
rect 0 12278 6979 12280
rect 0 12248 480 12278
rect 6913 12275 6979 12278
rect 15837 12338 15903 12341
rect 26509 12338 26575 12341
rect 29520 12338 30000 12368
rect 15837 12336 26575 12338
rect 15837 12280 15842 12336
rect 15898 12280 26514 12336
rect 26570 12280 26575 12336
rect 15837 12278 26575 12280
rect 15837 12275 15903 12278
rect 26509 12275 26575 12278
rect 26926 12278 30000 12338
rect 5257 12202 5323 12205
rect 7189 12202 7255 12205
rect 5257 12200 7255 12202
rect 5257 12144 5262 12200
rect 5318 12144 7194 12200
rect 7250 12144 7255 12200
rect 5257 12142 7255 12144
rect 5257 12139 5323 12142
rect 7189 12139 7255 12142
rect 14641 12202 14707 12205
rect 17585 12202 17651 12205
rect 25497 12202 25563 12205
rect 26785 12202 26851 12205
rect 26926 12202 26986 12278
rect 29520 12248 30000 12278
rect 14641 12200 17418 12202
rect 14641 12144 14646 12200
rect 14702 12144 17418 12200
rect 14641 12142 17418 12144
rect 14641 12139 14707 12142
rect 17358 12066 17418 12142
rect 17585 12200 25563 12202
rect 17585 12144 17590 12200
rect 17646 12144 25502 12200
rect 25558 12144 25563 12200
rect 17585 12142 25563 12144
rect 17585 12139 17651 12142
rect 25497 12139 25563 12142
rect 25822 12200 26986 12202
rect 25822 12144 26790 12200
rect 26846 12144 26986 12200
rect 25822 12142 26986 12144
rect 18873 12066 18939 12069
rect 19057 12066 19123 12069
rect 17358 12064 19123 12066
rect 17358 12008 18878 12064
rect 18934 12008 19062 12064
rect 19118 12008 19123 12064
rect 17358 12006 19123 12008
rect 18873 12003 18939 12006
rect 19057 12003 19123 12006
rect 20713 12066 20779 12069
rect 21633 12066 21699 12069
rect 25822 12066 25882 12142
rect 26785 12139 26851 12142
rect 20713 12064 25882 12066
rect 20713 12008 20718 12064
rect 20774 12008 21638 12064
rect 21694 12008 25882 12064
rect 20713 12006 25882 12008
rect 20713 12003 20779 12006
rect 21633 12003 21699 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 14641 11930 14707 11933
rect 12758 11928 14707 11930
rect 12758 11872 14646 11928
rect 14702 11872 14707 11928
rect 12758 11870 14707 11872
rect 8477 11794 8543 11797
rect 10777 11794 10843 11797
rect 12758 11794 12818 11870
rect 14641 11867 14707 11870
rect 8477 11792 12818 11794
rect 8477 11736 8482 11792
rect 8538 11736 10782 11792
rect 10838 11736 12818 11792
rect 8477 11734 12818 11736
rect 12985 11794 13051 11797
rect 25037 11794 25103 11797
rect 12985 11792 25103 11794
rect 12985 11736 12990 11792
rect 13046 11736 25042 11792
rect 25098 11736 25103 11792
rect 12985 11734 25103 11736
rect 8477 11731 8543 11734
rect 10777 11731 10843 11734
rect 12985 11731 13051 11734
rect 25037 11731 25103 11734
rect 0 11658 480 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 480 11598
rect 1485 11595 1551 11598
rect 3417 11658 3483 11661
rect 5073 11658 5139 11661
rect 18781 11658 18847 11661
rect 3417 11656 18847 11658
rect 3417 11600 3422 11656
rect 3478 11600 5078 11656
rect 5134 11600 18786 11656
rect 18842 11600 18847 11656
rect 3417 11598 18847 11600
rect 3417 11595 3483 11598
rect 5073 11595 5139 11598
rect 18781 11595 18847 11598
rect 26693 11658 26759 11661
rect 29520 11658 30000 11688
rect 26693 11656 30000 11658
rect 26693 11600 26698 11656
rect 26754 11600 30000 11656
rect 26693 11598 30000 11600
rect 26693 11595 26759 11598
rect 29520 11568 30000 11598
rect 5349 11522 5415 11525
rect 7925 11522 7991 11525
rect 5349 11520 7991 11522
rect 5349 11464 5354 11520
rect 5410 11464 7930 11520
rect 7986 11464 7991 11520
rect 5349 11462 7991 11464
rect 5349 11459 5415 11462
rect 7925 11459 7991 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 4613 11386 4679 11389
rect 7649 11386 7715 11389
rect 4613 11384 7715 11386
rect 4613 11328 4618 11384
rect 4674 11328 7654 11384
rect 7710 11328 7715 11384
rect 4613 11326 7715 11328
rect 4613 11323 4679 11326
rect 7649 11323 7715 11326
rect 2037 11250 2103 11253
rect 10317 11250 10383 11253
rect 11329 11250 11395 11253
rect 17125 11250 17191 11253
rect 2037 11248 11395 11250
rect 2037 11192 2042 11248
rect 2098 11192 10322 11248
rect 10378 11192 11334 11248
rect 11390 11192 11395 11248
rect 2037 11190 11395 11192
rect 2037 11187 2103 11190
rect 10317 11187 10383 11190
rect 11329 11187 11395 11190
rect 11470 11248 17191 11250
rect 11470 11192 17130 11248
rect 17186 11192 17191 11248
rect 11470 11190 17191 11192
rect 0 11114 480 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 480 11054
rect 1577 11051 1643 11054
rect 4061 11114 4127 11117
rect 7741 11114 7807 11117
rect 4061 11112 7807 11114
rect 4061 11056 4066 11112
rect 4122 11056 7746 11112
rect 7802 11056 7807 11112
rect 4061 11054 7807 11056
rect 4061 11051 4127 11054
rect 7741 11051 7807 11054
rect 7925 11114 7991 11117
rect 11470 11114 11530 11190
rect 17125 11187 17191 11190
rect 18781 11250 18847 11253
rect 26509 11250 26575 11253
rect 18781 11248 26575 11250
rect 18781 11192 18786 11248
rect 18842 11192 26514 11248
rect 26570 11192 26575 11248
rect 18781 11190 26575 11192
rect 18781 11187 18847 11190
rect 26509 11187 26575 11190
rect 13353 11116 13419 11117
rect 7925 11112 11530 11114
rect 7925 11056 7930 11112
rect 7986 11056 11530 11112
rect 7925 11054 11530 11056
rect 7925 11051 7991 11054
rect 13302 11052 13308 11116
rect 13372 11114 13419 11116
rect 26601 11114 26667 11117
rect 29520 11114 30000 11144
rect 13372 11112 13464 11114
rect 13414 11056 13464 11112
rect 13372 11054 13464 11056
rect 26601 11112 30000 11114
rect 26601 11056 26606 11112
rect 26662 11056 30000 11112
rect 26601 11054 30000 11056
rect 13372 11052 13419 11054
rect 13353 11051 13419 11052
rect 26601 11051 26667 11054
rect 29520 11024 30000 11054
rect 18505 10978 18571 10981
rect 25773 10978 25839 10981
rect 18505 10976 25839 10978
rect 18505 10920 18510 10976
rect 18566 10920 25778 10976
rect 25834 10920 25839 10976
rect 18505 10918 25839 10920
rect 18505 10915 18571 10918
rect 25773 10915 25839 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 2405 10842 2471 10845
rect 5349 10842 5415 10845
rect 2405 10840 5415 10842
rect 2405 10784 2410 10840
rect 2466 10784 5354 10840
rect 5410 10784 5415 10840
rect 2405 10782 5415 10784
rect 2405 10779 2471 10782
rect 5349 10779 5415 10782
rect 5441 10706 5507 10709
rect 14549 10706 14615 10709
rect 5441 10704 14615 10706
rect 5441 10648 5446 10704
rect 5502 10648 14554 10704
rect 14610 10648 14615 10704
rect 5441 10646 14615 10648
rect 5441 10643 5507 10646
rect 14549 10643 14615 10646
rect 14825 10706 14891 10709
rect 26969 10706 27035 10709
rect 27521 10706 27587 10709
rect 14825 10704 27587 10706
rect 14825 10648 14830 10704
rect 14886 10648 26974 10704
rect 27030 10648 27526 10704
rect 27582 10648 27587 10704
rect 14825 10646 27587 10648
rect 14825 10643 14891 10646
rect 26969 10643 27035 10646
rect 27521 10643 27587 10646
rect 2773 10570 2839 10573
rect 4429 10570 4495 10573
rect 2773 10568 4495 10570
rect 2773 10512 2778 10568
rect 2834 10512 4434 10568
rect 4490 10512 4495 10568
rect 2773 10510 4495 10512
rect 2773 10507 2839 10510
rect 4429 10507 4495 10510
rect 0 10434 480 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 480 10374
rect 1393 10371 1459 10374
rect 2865 10434 2931 10437
rect 4797 10434 4863 10437
rect 8661 10434 8727 10437
rect 2865 10432 8727 10434
rect 2865 10376 2870 10432
rect 2926 10376 4802 10432
rect 4858 10376 8666 10432
rect 8722 10376 8727 10432
rect 2865 10374 8727 10376
rect 2865 10371 2931 10374
rect 4797 10371 4863 10374
rect 8661 10371 8727 10374
rect 22185 10434 22251 10437
rect 24853 10434 24919 10437
rect 22185 10432 24919 10434
rect 22185 10376 22190 10432
rect 22246 10376 24858 10432
rect 24914 10376 24919 10432
rect 22185 10374 24919 10376
rect 22185 10371 22251 10374
rect 24853 10371 24919 10374
rect 25865 10434 25931 10437
rect 29520 10434 30000 10464
rect 25865 10432 30000 10434
rect 25865 10376 25870 10432
rect 25926 10376 30000 10432
rect 25865 10374 30000 10376
rect 25865 10371 25931 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 3233 10162 3299 10165
rect 4889 10162 4955 10165
rect 18597 10162 18663 10165
rect 3233 10160 18663 10162
rect 3233 10104 3238 10160
rect 3294 10104 4894 10160
rect 4950 10104 18602 10160
rect 18658 10104 18663 10160
rect 3233 10102 18663 10104
rect 3233 10099 3299 10102
rect 4889 10099 4955 10102
rect 18597 10099 18663 10102
rect 18137 10026 18203 10029
rect 26877 10026 26943 10029
rect 18137 10024 26943 10026
rect 18137 9968 18142 10024
rect 18198 9968 26882 10024
rect 26938 9968 26943 10024
rect 18137 9966 26943 9968
rect 18137 9963 18203 9966
rect 26877 9963 26943 9966
rect 0 9890 480 9920
rect 2681 9890 2747 9893
rect 0 9888 2747 9890
rect 0 9832 2686 9888
rect 2742 9832 2747 9888
rect 0 9830 2747 9832
rect 0 9800 480 9830
rect 2681 9827 2747 9830
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 2405 9618 2471 9621
rect 7097 9618 7163 9621
rect 12157 9618 12223 9621
rect 2405 9616 12223 9618
rect 2405 9560 2410 9616
rect 2466 9560 7102 9616
rect 7158 9560 12162 9616
rect 12218 9560 12223 9616
rect 2405 9558 12223 9560
rect 2405 9555 2471 9558
rect 7097 9555 7163 9558
rect 12157 9555 12223 9558
rect 15745 9618 15811 9621
rect 23749 9618 23815 9621
rect 15745 9616 23815 9618
rect 15745 9560 15750 9616
rect 15806 9560 23754 9616
rect 23810 9560 23815 9616
rect 15745 9558 23815 9560
rect 15745 9555 15811 9558
rect 23749 9555 23815 9558
rect 2037 9482 2103 9485
rect 18413 9482 18479 9485
rect 2037 9480 18479 9482
rect 2037 9424 2042 9480
rect 2098 9424 18418 9480
rect 18474 9424 18479 9480
rect 2037 9422 18479 9424
rect 2037 9419 2103 9422
rect 18413 9419 18479 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 14181 9346 14247 9349
rect 19701 9346 19767 9349
rect 14181 9344 19767 9346
rect 14181 9288 14186 9344
rect 14242 9288 19706 9344
rect 19762 9288 19767 9344
rect 14181 9286 19767 9288
rect 14181 9283 14247 9286
rect 19701 9283 19767 9286
rect 27613 9346 27679 9349
rect 29520 9346 30000 9376
rect 27613 9344 30000 9346
rect 27613 9288 27618 9344
rect 27674 9288 30000 9344
rect 27613 9286 30000 9288
rect 27613 9283 27679 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 2037 9074 2103 9077
rect 12065 9074 12131 9077
rect 2037 9072 12131 9074
rect 2037 9016 2042 9072
rect 2098 9016 12070 9072
rect 12126 9016 12131 9072
rect 2037 9014 12131 9016
rect 2037 9011 2103 9014
rect 12065 9011 12131 9014
rect 18597 9074 18663 9077
rect 26509 9074 26575 9077
rect 18597 9072 26575 9074
rect 18597 9016 18602 9072
rect 18658 9016 26514 9072
rect 26570 9016 26575 9072
rect 18597 9014 26575 9016
rect 18597 9011 18663 9014
rect 26509 9011 26575 9014
rect 12893 8938 12959 8941
rect 21265 8938 21331 8941
rect 23749 8938 23815 8941
rect 12893 8936 17970 8938
rect 12893 8880 12898 8936
rect 12954 8880 17970 8936
rect 12893 8878 17970 8880
rect 12893 8875 12959 8878
rect 7281 8802 7347 8805
rect 10409 8802 10475 8805
rect 7281 8800 10475 8802
rect 7281 8744 7286 8800
rect 7342 8744 10414 8800
rect 10470 8744 10475 8800
rect 7281 8742 10475 8744
rect 17910 8802 17970 8878
rect 21265 8936 23815 8938
rect 21265 8880 21270 8936
rect 21326 8880 23754 8936
rect 23810 8880 23815 8936
rect 21265 8878 23815 8880
rect 21265 8875 21331 8878
rect 23749 8875 23815 8878
rect 21817 8802 21883 8805
rect 25129 8802 25195 8805
rect 17910 8800 25195 8802
rect 17910 8744 21822 8800
rect 21878 8744 25134 8800
rect 25190 8744 25195 8800
rect 17910 8742 25195 8744
rect 7281 8739 7347 8742
rect 10409 8739 10475 8742
rect 21817 8739 21883 8742
rect 25129 8739 25195 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1577 8666 1643 8669
rect 0 8664 1643 8666
rect 0 8608 1582 8664
rect 1638 8608 1643 8664
rect 0 8606 1643 8608
rect 0 8576 480 8606
rect 1577 8603 1643 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 4981 8532 5047 8533
rect 4981 8530 5028 8532
rect 4936 8528 5028 8530
rect 4936 8472 4986 8528
rect 4936 8470 5028 8472
rect 4981 8468 5028 8470
rect 5092 8468 5098 8532
rect 20529 8530 20595 8533
rect 23289 8530 23355 8533
rect 20529 8528 23355 8530
rect 20529 8472 20534 8528
rect 20590 8472 23294 8528
rect 23350 8472 23355 8528
rect 20529 8470 23355 8472
rect 4981 8467 5047 8468
rect 20529 8467 20595 8470
rect 23289 8467 23355 8470
rect 23933 8530 23999 8533
rect 25405 8530 25471 8533
rect 23933 8528 25471 8530
rect 23933 8472 23938 8528
rect 23994 8472 25410 8528
rect 25466 8472 25471 8528
rect 23933 8470 25471 8472
rect 23933 8467 23999 8470
rect 25405 8467 25471 8470
rect 5717 8394 5783 8397
rect 9029 8394 9095 8397
rect 13261 8394 13327 8397
rect 15653 8394 15719 8397
rect 21265 8394 21331 8397
rect 5717 8392 21331 8394
rect 5717 8336 5722 8392
rect 5778 8336 9034 8392
rect 9090 8336 13266 8392
rect 13322 8336 15658 8392
rect 15714 8336 21270 8392
rect 21326 8336 21331 8392
rect 5717 8334 21331 8336
rect 5717 8331 5783 8334
rect 9029 8331 9095 8334
rect 13261 8331 13327 8334
rect 15653 8331 15719 8334
rect 21265 8331 21331 8334
rect 24209 8394 24275 8397
rect 26325 8394 26391 8397
rect 24209 8392 26391 8394
rect 24209 8336 24214 8392
rect 24270 8336 26330 8392
rect 26386 8336 26391 8392
rect 24209 8334 26391 8336
rect 24209 8331 24275 8334
rect 26325 8331 26391 8334
rect 4245 8258 4311 8261
rect 10133 8258 10199 8261
rect 4245 8256 10199 8258
rect 4245 8200 4250 8256
rect 4306 8200 10138 8256
rect 10194 8200 10199 8256
rect 4245 8198 10199 8200
rect 4245 8195 4311 8198
rect 10133 8195 10199 8198
rect 13997 8258 14063 8261
rect 19793 8258 19859 8261
rect 13997 8256 19859 8258
rect 13997 8200 14002 8256
rect 14058 8200 19798 8256
rect 19854 8200 19859 8256
rect 13997 8198 19859 8200
rect 13997 8195 14063 8198
rect 19793 8195 19859 8198
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 2681 8122 2747 8125
rect 0 8120 2747 8122
rect 0 8064 2686 8120
rect 2742 8064 2747 8120
rect 0 8062 2747 8064
rect 0 8032 480 8062
rect 2681 8059 2747 8062
rect 4981 8122 5047 8125
rect 9949 8122 10015 8125
rect 4981 8120 10015 8122
rect 4981 8064 4986 8120
rect 5042 8064 9954 8120
rect 10010 8064 10015 8120
rect 4981 8062 10015 8064
rect 4981 8059 5047 8062
rect 9949 8059 10015 8062
rect 11973 8122 12039 8125
rect 20069 8122 20135 8125
rect 11973 8120 20135 8122
rect 11973 8064 11978 8120
rect 12034 8064 20074 8120
rect 20130 8064 20135 8120
rect 11973 8062 20135 8064
rect 11973 8059 12039 8062
rect 20069 8059 20135 8062
rect 26601 8122 26667 8125
rect 29520 8122 30000 8152
rect 26601 8120 30000 8122
rect 26601 8064 26606 8120
rect 26662 8064 30000 8120
rect 26601 8062 30000 8064
rect 26601 8059 26667 8062
rect 29520 8032 30000 8062
rect 2497 7986 2563 7989
rect 4245 7986 4311 7989
rect 2497 7984 4311 7986
rect 2497 7928 2502 7984
rect 2558 7928 4250 7984
rect 4306 7928 4311 7984
rect 2497 7926 4311 7928
rect 2497 7923 2563 7926
rect 4245 7923 4311 7926
rect 6361 7986 6427 7989
rect 11789 7986 11855 7989
rect 16205 7986 16271 7989
rect 6361 7984 11855 7986
rect 6361 7928 6366 7984
rect 6422 7928 11794 7984
rect 11850 7928 11855 7984
rect 6361 7926 11855 7928
rect 6361 7923 6427 7926
rect 11789 7923 11855 7926
rect 11976 7984 16271 7986
rect 11976 7928 16210 7984
rect 16266 7928 16271 7984
rect 11976 7926 16271 7928
rect 3509 7850 3575 7853
rect 11976 7850 12036 7926
rect 16205 7923 16271 7926
rect 21265 7986 21331 7989
rect 26509 7986 26575 7989
rect 21265 7984 26575 7986
rect 21265 7928 21270 7984
rect 21326 7928 26514 7984
rect 26570 7928 26575 7984
rect 21265 7926 26575 7928
rect 21265 7923 21331 7926
rect 26509 7923 26575 7926
rect 3509 7848 12036 7850
rect 3509 7792 3514 7848
rect 3570 7792 12036 7848
rect 3509 7790 12036 7792
rect 3509 7787 3575 7790
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 19885 7578 19951 7581
rect 23105 7578 23171 7581
rect 19885 7576 23171 7578
rect 19885 7520 19890 7576
rect 19946 7520 23110 7576
rect 23166 7520 23171 7576
rect 19885 7518 23171 7520
rect 19885 7515 19951 7518
rect 23105 7515 23171 7518
rect 0 7442 480 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 480 7382
rect 1393 7379 1459 7382
rect 16573 7442 16639 7445
rect 27521 7442 27587 7445
rect 16573 7440 27587 7442
rect 16573 7384 16578 7440
rect 16634 7384 27526 7440
rect 27582 7384 27587 7440
rect 16573 7382 27587 7384
rect 16573 7379 16639 7382
rect 27521 7379 27587 7382
rect 27705 7442 27771 7445
rect 29520 7442 30000 7472
rect 27705 7440 30000 7442
rect 27705 7384 27710 7440
rect 27766 7384 30000 7440
rect 27705 7382 30000 7384
rect 27705 7379 27771 7382
rect 29520 7352 30000 7382
rect 1669 7306 1735 7309
rect 14825 7306 14891 7309
rect 1669 7304 14891 7306
rect 1669 7248 1674 7304
rect 1730 7248 14830 7304
rect 14886 7248 14891 7304
rect 1669 7246 14891 7248
rect 1669 7243 1735 7246
rect 14825 7243 14891 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 3141 7034 3207 7037
rect 10501 7034 10567 7037
rect 3141 7032 10567 7034
rect 3141 6976 3146 7032
rect 3202 6976 10506 7032
rect 10562 6976 10567 7032
rect 3141 6974 10567 6976
rect 3141 6971 3207 6974
rect 10501 6971 10567 6974
rect 11789 7034 11855 7037
rect 20437 7034 20503 7037
rect 11789 7032 20503 7034
rect 11789 6976 11794 7032
rect 11850 6976 20442 7032
rect 20498 6976 20503 7032
rect 11789 6974 20503 6976
rect 11789 6971 11855 6974
rect 20437 6971 20503 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 1853 6898 1919 6901
rect 4245 6898 4311 6901
rect 24945 6898 25011 6901
rect 1853 6896 4311 6898
rect 1853 6840 1858 6896
rect 1914 6840 4250 6896
rect 4306 6840 4311 6896
rect 1853 6838 4311 6840
rect 1853 6835 1919 6838
rect 4245 6835 4311 6838
rect 17358 6896 25011 6898
rect 17358 6840 24950 6896
rect 25006 6840 25011 6896
rect 17358 6838 25011 6840
rect 10133 6762 10199 6765
rect 17217 6762 17283 6765
rect 17358 6762 17418 6838
rect 24945 6835 25011 6838
rect 26693 6898 26759 6901
rect 29520 6898 30000 6928
rect 26693 6896 30000 6898
rect 26693 6840 26698 6896
rect 26754 6840 30000 6896
rect 26693 6838 30000 6840
rect 26693 6835 26759 6838
rect 29520 6808 30000 6838
rect 10133 6760 17418 6762
rect 10133 6704 10138 6760
rect 10194 6704 17222 6760
rect 17278 6704 17418 6760
rect 10133 6702 17418 6704
rect 10133 6699 10199 6702
rect 17217 6699 17283 6702
rect 16849 6626 16915 6629
rect 22645 6626 22711 6629
rect 16849 6624 22711 6626
rect 16849 6568 16854 6624
rect 16910 6568 22650 6624
rect 22706 6568 22711 6624
rect 16849 6566 22711 6568
rect 16849 6563 16915 6566
rect 22645 6563 22711 6566
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 3877 6354 3943 6357
rect 10409 6354 10475 6357
rect 15101 6354 15167 6357
rect 24577 6354 24643 6357
rect 3877 6352 24643 6354
rect 3877 6296 3882 6352
rect 3938 6296 10414 6352
rect 10470 6296 15106 6352
rect 15162 6296 24582 6352
rect 24638 6296 24643 6352
rect 3877 6294 24643 6296
rect 3877 6291 3943 6294
rect 10409 6291 10475 6294
rect 15101 6291 15167 6294
rect 24577 6291 24643 6294
rect 26601 6354 26667 6357
rect 29520 6354 30000 6384
rect 26601 6352 30000 6354
rect 26601 6296 26606 6352
rect 26662 6296 30000 6352
rect 26601 6294 30000 6296
rect 26601 6291 26667 6294
rect 29520 6264 30000 6294
rect 9121 6218 9187 6221
rect 16757 6218 16823 6221
rect 26417 6218 26483 6221
rect 9121 6216 26483 6218
rect 9121 6160 9126 6216
rect 9182 6160 16762 6216
rect 16818 6160 26422 6216
rect 26478 6160 26483 6216
rect 9121 6158 26483 6160
rect 9121 6155 9187 6158
rect 16757 6155 16823 6158
rect 26417 6155 26483 6158
rect 2589 6082 2655 6085
rect 3049 6082 3115 6085
rect 2589 6080 3115 6082
rect 2589 6024 2594 6080
rect 2650 6024 3054 6080
rect 3110 6024 3115 6080
rect 2589 6022 3115 6024
rect 2589 6019 2655 6022
rect 3049 6019 3115 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 2405 5946 2471 5949
rect 4245 5946 4311 5949
rect 2405 5944 4311 5946
rect 2405 5888 2410 5944
rect 2466 5888 4250 5944
rect 4306 5888 4311 5944
rect 2405 5886 4311 5888
rect 2405 5883 2471 5886
rect 4245 5883 4311 5886
rect 7741 5946 7807 5949
rect 10317 5946 10383 5949
rect 7741 5944 10383 5946
rect 7741 5888 7746 5944
rect 7802 5888 10322 5944
rect 10378 5888 10383 5944
rect 7741 5886 10383 5888
rect 7741 5883 7807 5886
rect 10317 5883 10383 5886
rect 7465 5810 7531 5813
rect 13629 5810 13695 5813
rect 7465 5808 13695 5810
rect 7465 5752 7470 5808
rect 7526 5752 13634 5808
rect 13690 5752 13695 5808
rect 7465 5750 13695 5752
rect 7465 5747 7531 5750
rect 13629 5747 13695 5750
rect 19885 5810 19951 5813
rect 23473 5810 23539 5813
rect 19885 5808 23539 5810
rect 19885 5752 19890 5808
rect 19946 5752 23478 5808
rect 23534 5752 23539 5808
rect 19885 5750 23539 5752
rect 19885 5747 19951 5750
rect 23473 5747 23539 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 4705 5674 4771 5677
rect 8845 5674 8911 5677
rect 16849 5674 16915 5677
rect 4705 5672 16915 5674
rect 4705 5616 4710 5672
rect 4766 5616 8850 5672
rect 8906 5616 16854 5672
rect 16910 5616 16915 5672
rect 4705 5614 16915 5616
rect 4705 5611 4771 5614
rect 8845 5611 8911 5614
rect 16849 5611 16915 5614
rect 26693 5674 26759 5677
rect 29520 5674 30000 5704
rect 26693 5672 30000 5674
rect 26693 5616 26698 5672
rect 26754 5616 30000 5672
rect 26693 5614 30000 5616
rect 26693 5611 26759 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 25865 5266 25931 5269
rect 25865 5264 26618 5266
rect 25865 5208 25870 5264
rect 25926 5208 26618 5264
rect 25865 5206 26618 5208
rect 25865 5203 25931 5206
rect 0 5130 480 5160
rect 1761 5130 1827 5133
rect 0 5128 1827 5130
rect 0 5072 1766 5128
rect 1822 5072 1827 5128
rect 0 5070 1827 5072
rect 0 5040 480 5070
rect 1761 5067 1827 5070
rect 15377 5130 15443 5133
rect 26417 5130 26483 5133
rect 15377 5128 26483 5130
rect 15377 5072 15382 5128
rect 15438 5072 26422 5128
rect 26478 5072 26483 5128
rect 15377 5070 26483 5072
rect 26558 5130 26618 5206
rect 29520 5130 30000 5160
rect 26558 5070 30000 5130
rect 15377 5067 15443 5070
rect 26417 5067 26483 5070
rect 29520 5040 30000 5070
rect 3601 4994 3667 4997
rect 8293 4994 8359 4997
rect 3601 4992 8359 4994
rect 3601 4936 3606 4992
rect 3662 4936 8298 4992
rect 8354 4936 8359 4992
rect 3601 4934 8359 4936
rect 3601 4931 3667 4934
rect 8293 4931 8359 4934
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 8569 4722 8635 4725
rect 11421 4722 11487 4725
rect 8569 4720 11487 4722
rect 8569 4664 8574 4720
rect 8630 4664 11426 4720
rect 11482 4664 11487 4720
rect 8569 4662 11487 4664
rect 8569 4659 8635 4662
rect 11421 4659 11487 4662
rect 21725 4722 21791 4725
rect 26509 4722 26575 4725
rect 21725 4720 26575 4722
rect 21725 4664 21730 4720
rect 21786 4664 26514 4720
rect 26570 4664 26575 4720
rect 21725 4662 26575 4664
rect 21725 4659 21791 4662
rect 26509 4659 26575 4662
rect 4797 4586 4863 4589
rect 5349 4586 5415 4589
rect 10317 4586 10383 4589
rect 14549 4586 14615 4589
rect 4797 4584 14615 4586
rect 4797 4528 4802 4584
rect 4858 4528 5354 4584
rect 5410 4528 10322 4584
rect 10378 4528 14554 4584
rect 14610 4528 14615 4584
rect 4797 4526 14615 4528
rect 4797 4523 4863 4526
rect 5349 4523 5415 4526
rect 10317 4523 10383 4526
rect 14549 4523 14615 4526
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 26601 4450 26667 4453
rect 29520 4450 30000 4480
rect 26601 4448 30000 4450
rect 26601 4392 26606 4448
rect 26662 4392 30000 4448
rect 26601 4390 30000 4392
rect 26601 4387 26667 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 4613 4178 4679 4181
rect 7281 4178 7347 4181
rect 13997 4178 14063 4181
rect 4613 4176 14063 4178
rect 4613 4120 4618 4176
rect 4674 4120 7286 4176
rect 7342 4120 14002 4176
rect 14058 4120 14063 4176
rect 4613 4118 14063 4120
rect 4613 4115 4679 4118
rect 7281 4115 7347 4118
rect 13997 4115 14063 4118
rect 26693 4176 26759 4181
rect 26693 4120 26698 4176
rect 26754 4120 26759 4176
rect 26693 4115 26759 4120
rect 1393 4042 1459 4045
rect 5625 4042 5691 4045
rect 1393 4040 5691 4042
rect 1393 3984 1398 4040
rect 1454 3984 5630 4040
rect 5686 3984 5691 4040
rect 1393 3982 5691 3984
rect 1393 3979 1459 3982
rect 5625 3979 5691 3982
rect 9581 4042 9647 4045
rect 11605 4042 11671 4045
rect 9581 4040 11671 4042
rect 9581 3984 9586 4040
rect 9642 3984 11610 4040
rect 11666 3984 11671 4040
rect 9581 3982 11671 3984
rect 9581 3979 9647 3982
rect 11605 3979 11671 3982
rect 21173 4042 21239 4045
rect 26509 4042 26575 4045
rect 21173 4040 26575 4042
rect 21173 3984 21178 4040
rect 21234 3984 26514 4040
rect 26570 3984 26575 4040
rect 21173 3982 26575 3984
rect 21173 3979 21239 3982
rect 26509 3979 26575 3982
rect 0 3906 480 3936
rect 2681 3906 2747 3909
rect 0 3904 2747 3906
rect 0 3848 2686 3904
rect 2742 3848 2747 3904
rect 0 3846 2747 3848
rect 0 3816 480 3846
rect 2681 3843 2747 3846
rect 3601 3906 3667 3909
rect 9397 3906 9463 3909
rect 3601 3904 9463 3906
rect 3601 3848 3606 3904
rect 3662 3848 9402 3904
rect 9458 3848 9463 3904
rect 3601 3846 9463 3848
rect 26696 3906 26756 4115
rect 29520 3906 30000 3936
rect 26696 3846 30000 3906
rect 3601 3843 3667 3846
rect 9397 3843 9463 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 657 3770 723 3773
rect 790 3770 796 3772
rect 657 3768 796 3770
rect 657 3712 662 3768
rect 718 3712 796 3768
rect 657 3710 796 3712
rect 657 3707 723 3710
rect 790 3708 796 3710
rect 860 3708 866 3772
rect 5165 3770 5231 3773
rect 10225 3770 10291 3773
rect 5165 3768 10291 3770
rect 5165 3712 5170 3768
rect 5226 3712 10230 3768
rect 10286 3712 10291 3768
rect 5165 3710 10291 3712
rect 5165 3707 5231 3710
rect 10225 3707 10291 3710
rect 21357 3770 21423 3773
rect 27245 3770 27311 3773
rect 21357 3768 27311 3770
rect 21357 3712 21362 3768
rect 21418 3712 27250 3768
rect 27306 3712 27311 3768
rect 21357 3710 27311 3712
rect 21357 3707 21423 3710
rect 27245 3707 27311 3710
rect 8293 3634 8359 3637
rect 26417 3634 26483 3637
rect 8293 3632 26483 3634
rect 8293 3576 8298 3632
rect 8354 3576 26422 3632
rect 26478 3576 26483 3632
rect 8293 3574 26483 3576
rect 8293 3571 8359 3574
rect 26417 3571 26483 3574
rect 4337 3498 4403 3501
rect 10133 3498 10199 3501
rect 4337 3496 10199 3498
rect 4337 3440 4342 3496
rect 4398 3440 10138 3496
rect 10194 3440 10199 3496
rect 4337 3438 10199 3440
rect 4337 3435 4403 3438
rect 10133 3435 10199 3438
rect 25497 3498 25563 3501
rect 25497 3496 27538 3498
rect 25497 3440 25502 3496
rect 25558 3440 27538 3496
rect 25497 3438 27538 3440
rect 25497 3435 25563 3438
rect 0 3362 480 3392
rect 3877 3362 3943 3365
rect 0 3360 3943 3362
rect 0 3304 3882 3360
rect 3938 3304 3943 3360
rect 0 3302 3943 3304
rect 27478 3362 27538 3438
rect 29520 3362 30000 3392
rect 27478 3302 30000 3362
rect 0 3272 480 3302
rect 3877 3299 3943 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 23749 3090 23815 3093
rect 27521 3090 27587 3093
rect 23749 3088 27587 3090
rect 23749 3032 23754 3088
rect 23810 3032 27526 3088
rect 27582 3032 27587 3088
rect 23749 3030 27587 3032
rect 23749 3027 23815 3030
rect 27521 3027 27587 3030
rect 26785 2818 26851 2821
rect 26785 2816 26986 2818
rect 26785 2760 26790 2816
rect 26846 2760 26986 2816
rect 26785 2758 26986 2760
rect 26785 2755 26851 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 4245 2682 4311 2685
rect 0 2680 4311 2682
rect 0 2624 4250 2680
rect 4306 2624 4311 2680
rect 0 2622 4311 2624
rect 26926 2682 26986 2758
rect 29520 2682 30000 2712
rect 26926 2622 30000 2682
rect 0 2592 480 2622
rect 4245 2619 4311 2622
rect 29520 2592 30000 2622
rect 5809 2546 5875 2549
rect 9765 2546 9831 2549
rect 5809 2544 9831 2546
rect 5809 2488 5814 2544
rect 5870 2488 9770 2544
rect 9826 2488 9831 2544
rect 5809 2486 9831 2488
rect 5809 2483 5875 2486
rect 9765 2483 9831 2486
rect 16297 2546 16363 2549
rect 24301 2546 24367 2549
rect 16297 2544 24367 2546
rect 16297 2488 16302 2544
rect 16358 2488 24306 2544
rect 24362 2488 24367 2544
rect 16297 2486 24367 2488
rect 16297 2483 16363 2486
rect 24301 2483 24367 2486
rect 2497 2410 2563 2413
rect 11973 2410 12039 2413
rect 2497 2408 12039 2410
rect 2497 2352 2502 2408
rect 2558 2352 11978 2408
rect 12034 2352 12039 2408
rect 2497 2350 12039 2352
rect 2497 2347 2563 2350
rect 11973 2347 12039 2350
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 5073 2138 5139 2141
rect 0 2136 5139 2138
rect 0 2080 5078 2136
rect 5134 2080 5139 2136
rect 0 2078 5139 2080
rect 0 2048 480 2078
rect 5073 2075 5139 2078
rect 27797 2138 27863 2141
rect 29520 2138 30000 2168
rect 27797 2136 30000 2138
rect 27797 2080 27802 2136
rect 27858 2080 30000 2136
rect 27797 2078 30000 2080
rect 27797 2075 27863 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 26693 1458 26759 1461
rect 29520 1458 30000 1488
rect 26693 1456 30000 1458
rect 26693 1400 26698 1456
rect 26754 1400 30000 1456
rect 26693 1398 30000 1400
rect 26693 1395 26759 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 4061 914 4127 917
rect 0 912 4127 914
rect 0 856 4066 912
rect 4122 856 4127 912
rect 0 854 4127 856
rect 0 824 480 854
rect 4061 851 4127 854
rect 25865 914 25931 917
rect 29520 914 30000 944
rect 25865 912 30000 914
rect 25865 856 25870 912
rect 25926 856 30000 912
rect 25865 854 30000 856
rect 25865 851 25931 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 3969 370 4035 373
rect 0 368 4035 370
rect 0 312 3974 368
rect 4030 312 4035 368
rect 0 310 4035 312
rect 0 280 480 310
rect 3969 307 4035 310
rect 26601 370 26667 373
rect 29520 370 30000 400
rect 26601 368 30000 370
rect 26601 312 26606 368
rect 26662 312 30000 368
rect 26601 310 30000 312
rect 26601 307 26667 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 18644 19136 18708 19140
rect 18644 19080 18658 19136
rect 18658 19080 18708 19136
rect 18644 19076 18708 19080
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 18644 18804 18708 18868
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 25084 15132 25148 15196
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 9812 13968 9876 13972
rect 9812 13912 9826 13968
rect 9826 13912 9876 13968
rect 9812 13908 9876 13912
rect 25636 13908 25700 13972
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 25084 12684 25148 12748
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 25084 12472 25148 12476
rect 25084 12416 25098 12472
rect 25098 12416 25148 12472
rect 25084 12412 25148 12416
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 13308 11112 13372 11116
rect 13308 11056 13358 11112
rect 13358 11056 13372 11112
rect 13308 11052 13372 11056
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 5028 8528 5092 8532
rect 5028 8472 5042 8528
rect 5042 8472 5092 8528
rect 5028 8468 5092 8472
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 796 3708 860 3772
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 18643 19140 18709 19141
rect 18643 19076 18644 19140
rect 18708 19076 18709 19140
rect 18643 19075 18709 19076
rect 18646 18869 18706 19075
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 18643 18868 18709 18869
rect 18643 18804 18644 18868
rect 18708 18804 18709 18868
rect 18643 18803 18709 18804
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 13307 11116 13373 11117
rect 13307 11052 13308 11116
rect 13372 11052 13373 11116
rect 13307 11051 13373 11052
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 13310 3858 13370 11051
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 18646 8618 18706 18803
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25083 15196 25149 15197
rect 25083 15132 25084 15196
rect 25148 15132 25149 15196
rect 25083 15131 25149 15132
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 25086 12749 25146 15131
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25083 12748 25149 12749
rect 25083 12684 25084 12748
rect 25148 12684 25149 12748
rect 25083 12683 25149 12684
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 25086 12477 25146 12683
rect 25083 12476 25149 12477
rect 25083 12412 25084 12476
rect 25148 12412 25149 12476
rect 25083 12411 25149 12412
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 9726 13972 9962 14058
rect 9726 13908 9812 13972
rect 9812 13908 9876 13972
rect 9876 13908 9962 13972
rect 9726 13822 9962 13908
rect 4942 8532 5178 8618
rect 4942 8468 5028 8532
rect 5028 8468 5092 8532
rect 5092 8468 5178 8532
rect 4942 8382 5178 8468
rect 710 3772 946 3858
rect 710 3708 796 3772
rect 796 3708 860 3772
rect 860 3708 946 3772
rect 710 3622 946 3708
rect 25550 13972 25786 14058
rect 25550 13908 25636 13972
rect 25636 13908 25700 13972
rect 25700 13908 25786 13972
rect 25550 13822 25786 13908
rect 18558 8382 18794 8618
rect 13222 3622 13458 3858
<< metal5 >>
rect 9684 14058 25828 14100
rect 9684 13822 9726 14058
rect 9962 13822 25550 14058
rect 25786 13822 25828 14058
rect 9684 13780 25828 13822
rect 4900 8618 18836 8660
rect 4900 8382 4942 8618
rect 5178 8382 18558 8618
rect 18794 8382 18836 8618
rect 4900 8340 18836 8382
rect 668 3858 13500 3900
rect 668 3622 710 3858
rect 946 3622 13222 3858
rect 13458 3622 13500 3858
rect 668 3580 13500 3622
use sky130_fd_sc_hd__fill_2  FILLER_1_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_49 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 1604681595
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7544 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6900 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80
timestamp 1604681595
transform 1 0 8464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_92
timestamp 1604681595
transform 1 0 9568 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11132 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1604681595
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1604681595
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1604681595
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16376 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_164
timestamp 1604681595
transform 1 0 16192 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_146
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_158
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_176
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_170
timestamp 1604681595
transform 1 0 16744 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1604681595
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_195
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18492 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1604681595
transform 1 0 19872 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_192
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_216
timestamp 1604681595
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_224
timestamp 1604681595
transform 1 0 21712 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1604681595
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24288 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_266
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp 1604681595
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_48
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_60
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_2_127
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_139
timestamp 1604681595
transform 1 0 13892 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1604681595
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18124 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1604681595
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_173
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_224
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_236
timestamp 1604681595
transform 1 0 22816 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_248
timestamp 1604681595
transform 1 0 23920 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_260
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1604681595
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1604681595
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_72
timestamp 1604681595
transform 1 0 7728 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_94
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1604681595
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_235
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1604681595
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_287
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_52
timestamp 1604681595
transform 1 0 5888 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_60
timestamp 1604681595
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_65
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_101
timestamp 1604681595
transform 1 0 10396 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_104
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_139
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_144
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1604681595
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_186
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_198
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_236
timestamp 1604681595
transform 1 0 22816 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_248
timestamp 1604681595
transform 1 0 23920 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_260
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_272
timestamp 1604681595
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_14
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 4048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_24
timestamp 1604681595
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1604681595
transform 1 0 3680 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1604681595
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_90
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_102
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_161
timestamp 1604681595
transform 1 0 15916 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_192
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_203
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_229
timestamp 1604681595
transform 1 0 22172 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_234
timestamp 1604681595
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_238
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_287
timestamp 1604681595
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_25
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1604681595
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_40
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5980 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1604681595
transform 1 0 5888 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_49
timestamp 1604681595
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_99
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_109
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_134
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp 1604681595
transform 1 0 13156 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_142
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_143
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_131
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_160
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_156
timestamp 1604681595
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_162
timestamp 1604681595
transform 1 0 16008 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_158
timestamp 1604681595
transform 1 0 15640 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1604681595
transform 1 0 16560 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_194
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_199
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1604681595
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 21620 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1604681595
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23920 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_237
timestamp 1604681595
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_267
timestamp 1604681595
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_287
timestamp 1604681595
transform 1 0 27508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_14
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_18
timestamp 1604681595
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1604681595
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_39
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_72
timestamp 1604681595
transform 1 0 7728 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604681595
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1604681595
transform 1 0 16560 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_181
timestamp 1604681595
transform 1 0 17756 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_244
timestamp 1604681595
transform 1 0 23552 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1604681595
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_255
timestamp 1604681595
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_52
timestamp 1604681595
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1604681595
transform 1 0 6256 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1604681595
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1604681595
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1604681595
transform 1 0 8924 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1604681595
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_99
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_112
timestamp 1604681595
transform 1 0 11408 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_139
timestamp 1604681595
transform 1 0 13892 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_145
timestamp 1604681595
transform 1 0 14444 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14720 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_167
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_192
timestamp 1604681595
transform 1 0 18768 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_231
timestamp 1604681595
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_235
timestamp 1604681595
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_270
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_274
timestamp 1604681595
transform 1 0 26312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604681595
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604681595
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_291
timestamp 1604681595
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1604681595
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_14
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_19
timestamp 1604681595
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_50
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_57
timestamp 1604681595
transform 1 0 6348 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12052 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_106
timestamp 1604681595
transform 1 0 10856 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1604681595
transform 1 0 11592 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp 1604681595
transform 1 0 11960 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_138
timestamp 1604681595
transform 1 0 13800 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1604681595
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1604681595
transform 1 0 16560 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_188
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_194
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_236
timestamp 1604681595
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_240
timestamp 1604681595
transform 1 0 23184 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1604681595
transform 1 0 24380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_268
timestamp 1604681595
transform 1 0 25760 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_19
timestamp 1604681595
transform 1 0 2852 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1604681595
transform 1 0 3220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_34
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1604681595
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1604681595
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7360 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_77
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1604681595
transform 1 0 9752 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1604681595
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_126
timestamp 1604681595
transform 1 0 12696 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_138
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_150
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1604681595
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1604681595
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_207
timestamp 1604681595
transform 1 0 20148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_219
timestamp 1604681595
transform 1 0 21252 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_227
timestamp 1604681595
transform 1 0 21988 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_262
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 27508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_285
timestamp 1604681595
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_289
timestamp 1604681595
transform 1 0 27692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1604681595
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1604681595
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp 1604681595
transform 1 0 5980 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604681595
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_104
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1604681595
transform 1 0 11040 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1604681595
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1604681595
transform 1 0 13708 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17388 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_168
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_176
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_186
timestamp 1604681595
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_194
timestamp 1604681595
transform 1 0 18952 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_223
timestamp 1604681595
transform 1 0 21620 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23000 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_233
timestamp 1604681595
transform 1 0 22540 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_237
timestamp 1604681595
transform 1 0 22908 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_247
timestamp 1604681595
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1604681595
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_260
timestamp 1604681595
transform 1 0 25024 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_268
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_284
timestamp 1604681595
transform 1 0 27232 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1604681595
transform 1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_22
timestamp 1604681595
transform 1 0 3128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_38
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_42
timestamp 1604681595
transform 1 0 4968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_52
timestamp 1604681595
transform 1 0 5888 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_70
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_72
timestamp 1604681595
transform 1 0 7728 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_92
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_107
timestamp 1604681595
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1604681595
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1604681595
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp 1604681595
transform 1 0 17296 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_167
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_213
timestamp 1604681595
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1604681595
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_234
timestamp 1604681595
transform 1 0 22632 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_230
timestamp 1604681595
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22356 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp 1604681595
transform 1 0 23828 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1604681595
transform 1 0 23552 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_240
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1604681595
transform 1 0 24472 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_264
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_260
timestamp 1604681595
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1604681595
transform 1 0 26680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 26864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_290
timestamp 1604681595
transform 1 0 27784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_282
timestamp 1604681595
transform 1 0 27048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 27416 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_285
timestamp 1604681595
transform 1 0 27324 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 27968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_294
timestamp 1604681595
transform 1 0 28152 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1604681595
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1604681595
transform 1 0 28428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp 1604681595
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_45
timestamp 1604681595
transform 1 0 5244 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_77
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_101
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_148
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_166
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_190
timestamp 1604681595
transform 1 0 18584 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_234
timestamp 1604681595
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_238
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 24196 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 26680 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_49
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_76
timestamp 1604681595
transform 1 0 8096 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_123
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1604681595
transform 1 0 13524 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_180
timestamp 1604681595
transform 1 0 17664 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1604681595
transform 1 0 19228 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1604681595
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_223
timestamp 1604681595
transform 1 0 21620 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_246
timestamp 1604681595
transform 1 0 23736 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1604681595
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_52
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604681595
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13340 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1604681595
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_260
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_268
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 26404 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 27324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_279
timestamp 1604681595
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_283
timestamp 1604681595
transform 1 0 27140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_287
timestamp 1604681595
transform 1 0 27508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_10
timestamp 1604681595
transform 1 0 2024 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4600 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_47
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_69
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_81
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_101
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_113
timestamp 1604681595
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_160
timestamp 1604681595
transform 1 0 15824 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_172
timestamp 1604681595
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_183
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_195
timestamp 1604681595
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_199
timestamp 1604681595
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1604681595
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_234
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_248
timestamp 1604681595
transform 1 0 23920 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_256
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 27048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_280
timestamp 1604681595
transform 1 0 26864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_284
timestamp 1604681595
transform 1 0 27232 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604681595
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_23
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_50
timestamp 1604681595
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_80
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_73
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_115
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1604681595
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_153
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1604681595
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1604681595
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_174
timestamp 1604681595
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_179
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1604681595
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1604681595
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_204
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_209
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_221
timestamp 1604681595
transform 1 0 21436 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_227
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1604681595
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_231
timestamp 1604681595
transform 1 0 22356 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1604681595
transform 1 0 22632 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23736 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_20_258
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_255
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_255
timestamp 1604681595
transform 1 0 24564 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_269
timestamp 1604681595
transform 1 0 25852 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_266
timestamp 1604681595
transform 1 0 25576 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_263
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_280
timestamp 1604681595
transform 1 0 26864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 27048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 27232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_285
timestamp 1604681595
transform 1 0 27324 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_287
timestamp 1604681595
transform 1 0 27508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1604681595
transform 1 0 28428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_11
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1604681595
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1604681595
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_78
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_100
timestamp 1604681595
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1604681595
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1604681595
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20148 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_192
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1604681595
transform 1 0 19872 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_226
timestamp 1604681595
transform 1 0 21896 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_235
timestamp 1604681595
transform 1 0 22724 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1604681595
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1604681595
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24656 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_252
timestamp 1604681595
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_265
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 26220 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 26036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_282
timestamp 1604681595
transform 1 0 27048 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_294
timestamp 1604681595
transform 1 0 28152 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1604681595
transform 1 0 28520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_22
timestamp 1604681595
transform 1 0 3128 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1604681595
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_57
timestamp 1604681595
transform 1 0 6348 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_74
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1604681595
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_86
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp 1604681595
transform 1 0 12236 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_158
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_171
timestamp 1604681595
transform 1 0 16836 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22540 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_252
timestamp 1604681595
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_256
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_268
timestamp 1604681595
transform 1 0 25760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 26680 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 27048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 26036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_273
timestamp 1604681595
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_280
timestamp 1604681595
transform 1 0 26864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_284
timestamp 1604681595
transform 1 0 27232 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_13
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1604681595
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_49
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1604681595
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_103
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1604681595
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15088 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_161
timestamp 1604681595
transform 1 0 15916 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_198
timestamp 1604681595
transform 1 0 19320 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1604681595
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_214
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_226
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_235
timestamp 1604681595
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_239
timestamp 1604681595
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1604681595
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23276 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_250
timestamp 1604681595
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_263
timestamp 1604681595
transform 1 0 25300 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26036 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_23_290
timestamp 1604681595
transform 1 0 27784 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1604681595
transform 1 0 28520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_26
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1604681595
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5796 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_49
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_122
timestamp 1604681595
transform 1 0 12328 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1604681595
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_158
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16652 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_188
timestamp 1604681595
transform 1 0 18400 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_194
timestamp 1604681595
transform 1 0 18952 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1604681595
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1604681595
transform 1 0 20148 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_223
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22908 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_235
timestamp 1604681595
transform 1 0 22724 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1604681595
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1604681595
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_254
timestamp 1604681595
transform 1 0 24472 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1604681595
transform 1 0 25576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_270
timestamp 1604681595
transform 1 0 25944 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_285
timestamp 1604681595
transform 1 0 27324 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1604681595
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1604681595
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_35
timestamp 1604681595
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_76
timestamp 1604681595
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13708 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1604681595
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_146
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_163
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_195
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_270
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_278
timestamp 1604681595
transform 1 0 26680 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_290
timestamp 1604681595
transform 1 0 27784 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1604681595
transform 1 0 28520 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1604681595
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_22
timestamp 1604681595
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_22
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_26
timestamp 1604681595
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1604681595
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1604681595
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_30
timestamp 1604681595
transform 1 0 3864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_55
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_92
timestamp 1604681595
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_88
timestamp 1604681595
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_100
timestamp 1604681595
transform 1 0 10304 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_110
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_109
timestamp 1604681595
transform 1 0 11132 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp 1604681595
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1604681595
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_156
timestamp 1604681595
transform 1 0 15456 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_152
timestamp 1604681595
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_162
timestamp 1604681595
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1604681595
transform 1 0 16652 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1604681595
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_204
timestamp 1604681595
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1604681595
transform 1 0 20976 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_224
timestamp 1604681595
transform 1 0 21712 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_223
timestamp 1604681595
transform 1 0 21620 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_229
timestamp 1604681595
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_237
timestamp 1604681595
transform 1 0 22908 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_242
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_262
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 1604681595
transform 1 0 25852 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1604681595
transform 1 0 25484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1604681595
transform 1 0 24380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_272
timestamp 1604681595
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_280
timestamp 1604681595
transform 1 0 26864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_289
timestamp 1604681595
transform 1 0 27692 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_292
timestamp 1604681595
transform 1 0 27968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1604681595
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp 1604681595
transform 1 0 28428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_21
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1604681595
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10120 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9936 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_107
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_119
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_128
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_162
timestamp 1604681595
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_182
timestamp 1604681595
transform 1 0 17848 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_188
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1604681595
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_219
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23184 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_232
timestamp 1604681595
transform 1 0 22448 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_238
timestamp 1604681595
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1604681595
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1604681595
transform 1 0 25484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1604681595
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604681595
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_50
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_58
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_84
timestamp 1604681595
transform 1 0 8832 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_96
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_105
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1604681595
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1604681595
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1604681595
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1604681595
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1604681595
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_227
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_254
timestamp 1604681595
transform 1 0 24472 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_287
timestamp 1604681595
transform 1 0 27508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_14
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_26
timestamp 1604681595
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604681595
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_51
timestamp 1604681595
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1604681595
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_79
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_83
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604681595
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1604681595
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18860 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 22816 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_245
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1604681595
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_257
timestamp 1604681595
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_260
timestamp 1604681595
transform 1 0 25024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604681595
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_78
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_100
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_112
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15088 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1604681595
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18676 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_200
timestamp 1604681595
transform 1 0 19504 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_224
timestamp 1604681595
transform 1 0 21712 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_249
timestamp 1604681595
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24196 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_253
timestamp 1604681595
transform 1 0 24380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_277
timestamp 1604681595
transform 1 0 26588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_289
timestamp 1604681595
transform 1 0 27692 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1604681595
transform 1 0 28428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_135
timestamp 1604681595
transform 1 0 13524 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_138
timestamp 1604681595
transform 1 0 13800 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1604681595
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 21344 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_219
timestamp 1604681595
transform 1 0 21252 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_224
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_32_236
timestamp 1604681595
transform 1 0 22816 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_242
timestamp 1604681595
transform 1 0 23368 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_262
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1604681595
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604681595
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_131
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_155
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_167
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1604681595
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 22264 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_249
timestamp 1604681595
transform 1 0 24012 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_261
timestamp 1604681595
transform 1 0 25116 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 26036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 26588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_275
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_279
timestamp 1604681595
transform 1 0 26772 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_291
timestamp 1604681595
transform 1 0 27876 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1604681595
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 27710 0 27766 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 7470 23520 7526 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 29182 0 29238 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 22466 23520 22522 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 bottom_grid_pin_11_
port 6 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 bottom_grid_pin_13_
port 8 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 bottom_grid_pin_14_
port 9 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 bottom_grid_pin_15_
port 10 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 bottom_grid_pin_1_
port 11 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 bottom_grid_pin_2_
port 12 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 bottom_grid_pin_3_
port 13 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 bottom_grid_pin_4_
port 14 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 bottom_grid_pin_5_
port 15 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 bottom_grid_pin_6_
port 16 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 bottom_grid_pin_7_
port 17 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_8_
port 18 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 bottom_grid_pin_9_
port 19 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 ccff_head
port 20 nsew default input
rlabel metal2 s 3514 0 3570 480 6 ccff_tail
port 21 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 22 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 23 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 24 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 25 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 26 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 27 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 28 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 29 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 30 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 31 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 32 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 33 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 34 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 35 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 36 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 37 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 38 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 39 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 40 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 41 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 43 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 44 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 45 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 46 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 47 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 48 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 49 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 50 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 51 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 52 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 53 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 54 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 55 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 56 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 57 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 58 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 59 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 60 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 61 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 62 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 63 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 64 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 65 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 66 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 67 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 68 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 69 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 70 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 71 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 72 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 73 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 74 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 75 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 76 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 77 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 78 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 79 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 80 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 81 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 82 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 83 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 84 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 85 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 86 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 87 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 88 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 89 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 90 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 91 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 92 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 93 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 94 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 95 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 96 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 97 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 98 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 99 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 100 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 101 nsew default tristate
rlabel metal2 s 662 0 718 480 6 prog_clk
port 102 nsew default input
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 103 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 104 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
