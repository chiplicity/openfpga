VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 122.000 BY 122.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 118.000 85.010 122.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 118.000 88.230 122.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 34.040 122.000 34.640 ;
    END
  END Test_en_E_in
  PIN Test_en_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 30.640 122.000 31.240 ;
    END
  END Test_en_E_out
  PIN Test_en_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END Test_en_W_in
  PIN Test_en_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END Test_en_W_out
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 27.240 122.000 27.840 ;
    END
  END ccff_tail
  PIN clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 118.000 91.450 122.000 ;
    END
  END clk_0_N_in
  PIN clk_0_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END clk_0_S_in
  PIN prog_clk_0_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 40.840 122.000 41.440 ;
    END
  END prog_clk_0_E_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 37.440 122.000 38.040 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 118.000 94.670 122.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END prog_clk_0_W_out
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 43.560 122.000 44.160 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 46.960 122.000 47.560 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 50.360 122.000 50.960 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 53.760 122.000 54.360 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 57.160 122.000 57.760 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 60.560 122.000 61.160 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 63.280 122.000 63.880 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 66.680 122.000 67.280 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 70.080 122.000 70.680 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 73.480 122.000 74.080 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 76.880 122.000 77.480 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 80.280 122.000 80.880 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 83.000 122.000 83.600 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 86.400 122.000 87.000 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 89.800 122.000 90.400 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 118.000 93.200 122.000 93.800 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 1.400 122.000 2.000 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 96.600 122.000 97.200 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 4.120 122.000 4.720 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 100.000 122.000 100.600 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 7.520 122.000 8.120 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 102.720 122.000 103.320 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 10.920 122.000 11.520 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 106.120 122.000 106.720 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 14.320 122.000 14.920 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 109.520 122.000 110.120 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 17.720 122.000 18.320 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 112.920 122.000 113.520 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 21.120 122.000 21.720 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 116.320 122.000 116.920 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 23.840 122.000 24.440 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 118.000 119.720 122.000 120.320 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 118.000 27.050 122.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 118.000 59.250 122.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 118.000 62.470 122.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 118.000 65.690 122.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 118.000 68.910 122.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 118.000 72.130 122.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 118.000 75.350 122.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 118.000 30.270 122.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 118.000 33.490 122.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 118.000 78.570 122.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 118.000 81.790 122.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 118.000 97.890 122.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.470 118.000 1.750 122.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 118.000 101.110 122.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.230 118.000 4.510 122.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 118.000 104.330 122.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 118.000 7.730 122.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 118.000 107.550 122.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 118.000 10.950 122.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 118.000 110.770 122.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 118.000 14.170 122.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 118.000 113.990 122.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 118.000 17.390 122.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 118.000 36.710 122.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 118.000 117.210 122.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 118.000 20.610 122.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 118.000 120.430 122.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.550 118.000 23.830 122.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 118.000 39.930 122.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 118.000 43.150 122.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 118.000 46.370 122.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 118.000 49.590 122.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 118.000 52.810 122.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 118.000 56.030 122.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.215 10.640 24.815 109.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.705 10.640 43.305 109.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 117.155 110.755 ;
      LAYER met1 ;
        RECT 1.450 9.560 120.450 114.540 ;
      LAYER met2 ;
        RECT 2.030 117.720 3.950 120.205 ;
        RECT 4.790 117.720 7.170 120.205 ;
        RECT 8.010 117.720 10.390 120.205 ;
        RECT 11.230 117.720 13.610 120.205 ;
        RECT 14.450 117.720 16.830 120.205 ;
        RECT 17.670 117.720 20.050 120.205 ;
        RECT 20.890 117.720 23.270 120.205 ;
        RECT 24.110 117.720 26.490 120.205 ;
        RECT 27.330 117.720 29.710 120.205 ;
        RECT 30.550 117.720 32.930 120.205 ;
        RECT 33.770 117.720 36.150 120.205 ;
        RECT 36.990 117.720 39.370 120.205 ;
        RECT 40.210 117.720 42.590 120.205 ;
        RECT 43.430 117.720 45.810 120.205 ;
        RECT 46.650 117.720 49.030 120.205 ;
        RECT 49.870 117.720 52.250 120.205 ;
        RECT 53.090 117.720 55.470 120.205 ;
        RECT 56.310 117.720 58.690 120.205 ;
        RECT 59.530 117.720 61.910 120.205 ;
        RECT 62.750 117.720 65.130 120.205 ;
        RECT 65.970 117.720 68.350 120.205 ;
        RECT 69.190 117.720 71.570 120.205 ;
        RECT 72.410 117.720 74.790 120.205 ;
        RECT 75.630 117.720 78.010 120.205 ;
        RECT 78.850 117.720 81.230 120.205 ;
        RECT 82.070 117.720 84.450 120.205 ;
        RECT 85.290 117.720 87.670 120.205 ;
        RECT 88.510 117.720 90.890 120.205 ;
        RECT 91.730 117.720 94.110 120.205 ;
        RECT 94.950 117.720 97.330 120.205 ;
        RECT 98.170 117.720 100.550 120.205 ;
        RECT 101.390 117.720 103.770 120.205 ;
        RECT 104.610 117.720 106.990 120.205 ;
        RECT 107.830 117.720 110.210 120.205 ;
        RECT 111.050 117.720 113.430 120.205 ;
        RECT 114.270 117.720 116.650 120.205 ;
        RECT 117.490 117.720 119.870 120.205 ;
        RECT 1.480 4.280 120.420 117.720 ;
        RECT 1.480 1.515 8.090 4.280 ;
        RECT 8.930 1.515 25.110 4.280 ;
        RECT 25.950 1.515 42.590 4.280 ;
        RECT 43.430 1.515 60.070 4.280 ;
        RECT 60.910 1.515 77.550 4.280 ;
        RECT 78.390 1.515 95.030 4.280 ;
        RECT 95.870 1.515 112.510 4.280 ;
        RECT 113.350 1.515 120.420 4.280 ;
      LAYER met3 ;
        RECT 4.000 119.320 117.600 120.185 ;
        RECT 4.000 117.320 118.000 119.320 ;
        RECT 4.000 115.920 117.600 117.320 ;
        RECT 4.000 113.920 118.000 115.920 ;
        RECT 4.000 112.520 117.600 113.920 ;
        RECT 4.000 110.520 118.000 112.520 ;
        RECT 4.000 109.120 117.600 110.520 ;
        RECT 4.000 107.120 118.000 109.120 ;
        RECT 4.400 105.720 117.600 107.120 ;
        RECT 4.000 103.720 118.000 105.720 ;
        RECT 4.000 102.320 117.600 103.720 ;
        RECT 4.000 101.000 118.000 102.320 ;
        RECT 4.000 99.600 117.600 101.000 ;
        RECT 4.000 97.600 118.000 99.600 ;
        RECT 4.000 96.200 117.600 97.600 ;
        RECT 4.000 94.200 118.000 96.200 ;
        RECT 4.000 92.800 117.600 94.200 ;
        RECT 4.000 90.800 118.000 92.800 ;
        RECT 4.000 89.400 117.600 90.800 ;
        RECT 4.000 87.400 118.000 89.400 ;
        RECT 4.000 86.000 117.600 87.400 ;
        RECT 4.000 84.000 118.000 86.000 ;
        RECT 4.000 82.600 117.600 84.000 ;
        RECT 4.000 81.280 118.000 82.600 ;
        RECT 4.000 79.880 117.600 81.280 ;
        RECT 4.000 77.880 118.000 79.880 ;
        RECT 4.000 76.520 117.600 77.880 ;
        RECT 4.400 76.480 117.600 76.520 ;
        RECT 4.400 75.120 118.000 76.480 ;
        RECT 4.000 74.480 118.000 75.120 ;
        RECT 4.000 73.080 117.600 74.480 ;
        RECT 4.000 71.080 118.000 73.080 ;
        RECT 4.000 69.680 117.600 71.080 ;
        RECT 4.000 67.680 118.000 69.680 ;
        RECT 4.000 66.280 117.600 67.680 ;
        RECT 4.000 64.280 118.000 66.280 ;
        RECT 4.000 62.880 117.600 64.280 ;
        RECT 4.000 61.560 118.000 62.880 ;
        RECT 4.000 60.160 117.600 61.560 ;
        RECT 4.000 58.160 118.000 60.160 ;
        RECT 4.000 56.760 117.600 58.160 ;
        RECT 4.000 54.760 118.000 56.760 ;
        RECT 4.000 53.360 117.600 54.760 ;
        RECT 4.000 51.360 118.000 53.360 ;
        RECT 4.000 49.960 117.600 51.360 ;
        RECT 4.000 47.960 118.000 49.960 ;
        RECT 4.000 46.560 117.600 47.960 ;
        RECT 4.000 45.920 118.000 46.560 ;
        RECT 4.400 44.560 118.000 45.920 ;
        RECT 4.400 44.520 117.600 44.560 ;
        RECT 4.000 43.160 117.600 44.520 ;
        RECT 4.000 41.840 118.000 43.160 ;
        RECT 4.000 40.440 117.600 41.840 ;
        RECT 4.000 38.440 118.000 40.440 ;
        RECT 4.000 37.040 117.600 38.440 ;
        RECT 4.000 35.040 118.000 37.040 ;
        RECT 4.000 33.640 117.600 35.040 ;
        RECT 4.000 31.640 118.000 33.640 ;
        RECT 4.000 30.240 117.600 31.640 ;
        RECT 4.000 28.240 118.000 30.240 ;
        RECT 4.000 26.840 117.600 28.240 ;
        RECT 4.000 24.840 118.000 26.840 ;
        RECT 4.000 23.440 117.600 24.840 ;
        RECT 4.000 22.120 118.000 23.440 ;
        RECT 4.000 20.720 117.600 22.120 ;
        RECT 4.000 18.720 118.000 20.720 ;
        RECT 4.000 17.320 117.600 18.720 ;
        RECT 4.000 16.000 118.000 17.320 ;
        RECT 4.400 15.320 118.000 16.000 ;
        RECT 4.400 14.600 117.600 15.320 ;
        RECT 4.000 13.920 117.600 14.600 ;
        RECT 4.000 11.920 118.000 13.920 ;
        RECT 4.000 10.520 117.600 11.920 ;
        RECT 4.000 8.520 118.000 10.520 ;
        RECT 4.000 7.120 117.600 8.520 ;
        RECT 4.000 5.120 118.000 7.120 ;
        RECT 4.000 3.720 117.600 5.120 ;
        RECT 4.000 2.400 118.000 3.720 ;
        RECT 4.000 1.535 117.600 2.400 ;
      LAYER met4 ;
        RECT 25.215 10.640 41.305 109.040 ;
        RECT 43.705 10.640 108.265 109.040 ;
  END
END grid_clb
END LIBRARY

