VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__1_
  CLASS BLOCK ;
  FOREIGN cbx_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 85.000 ;
  PIN REGIN_FEEDTHROUGH
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 83.680 100.000 84.280 ;
    END
  END REGIN_FEEDTHROUGH
  PIN REGOUT_FEEDTHROUGH
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 82.600 91.450 85.000 ;
    END
  END REGOUT_FEEDTHROUGH
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.370 82.600 8.650 85.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 82.600 25.210 85.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END bottom_grid_pin_11_
  PIN bottom_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END bottom_grid_pin_12_
  PIN bottom_grid_pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END bottom_grid_pin_13_
  PIN bottom_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.400 ;
    END
  END bottom_grid_pin_14_
  PIN bottom_grid_pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.400 ;
    END
  END bottom_grid_pin_15_
  PIN bottom_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END bottom_grid_pin_1_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END bottom_grid_pin_3_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END bottom_grid_pin_5_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.400 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 2.400 ;
    END
  END bottom_grid_pin_7_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END bottom_grid_pin_8_
  PIN bottom_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END bottom_grid_pin_9_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 2.400 35.320 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 2.400 60.480 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 2.400 62.520 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.400 63.880 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 2.400 40.080 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 2.400 18.320 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.400 6.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.400 11.520 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 51.040 100.000 51.640 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 67.360 100.000 67.960 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 68.720 100.000 69.320 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 70.760 100.000 71.360 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 72.120 100.000 72.720 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 74.160 100.000 74.760 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 75.520 100.000 76.120 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 76.880 100.000 77.480 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 78.920 100.000 79.520 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 80.280 100.000 80.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 82.320 100.000 82.920 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 52.400 100.000 53.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 54.440 100.000 55.040 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 55.800 100.000 56.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 57.840 100.000 58.440 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 59.200 100.000 59.800 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 60.560 100.000 61.160 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 62.600 100.000 63.200 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 63.960 100.000 64.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 66.000 100.000 66.600 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 18.400 100.000 19.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 34.720 100.000 35.320 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 36.080 100.000 36.680 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 38.120 100.000 38.720 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 39.480 100.000 40.080 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 41.520 100.000 42.120 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 42.880 100.000 43.480 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 44.240 100.000 44.840 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 46.280 100.000 46.880 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 47.640 100.000 48.240 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 49.680 100.000 50.280 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 19.760 100.000 20.360 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 21.800 100.000 22.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 23.160 100.000 23.760 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 25.200 100.000 25.800 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 26.560 100.000 27.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 27.920 100.000 28.520 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 29.960 100.000 30.560 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 31.320 100.000 31.920 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 33.360 100.000 33.960 ;
    END
  END chanx_right_out[9]
  PIN clk_1_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 17.040 100.000 17.640 ;
    END
  END clk_1_E_in
  PIN clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 82.600 41.770 85.000 ;
    END
  END clk_1_N_out
  PIN clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END clk_1_S_out
  PIN clk_1_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 2.400 84.280 ;
    END
  END clk_1_W_in
  PIN clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 15.000 100.000 15.600 ;
    END
  END clk_2_E_in
  PIN clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 6.840 100.000 7.440 ;
    END
  END clk_2_E_out
  PIN clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 2.400 74.080 ;
    END
  END clk_2_W_out
  PIN clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 13.640 100.000 14.240 ;
    END
  END clk_3_E_in
  PIN clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 5.480 100.000 6.080 ;
    END
  END clk_3_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END clk_3_W_in
  PIN clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END clk_3_W_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 82.600 58.330 85.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 82.600 74.890 85.000 ;
    END
  END prog_clk_0_W_out
  PIN prog_clk_1_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 11.600 100.000 12.200 ;
    END
  END prog_clk_1_E_in
  PIN prog_clk_1_N_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 3.440 100.000 4.040 ;
    END
  END prog_clk_1_N_out
  PIN prog_clk_1_S_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END prog_clk_1_S_out
  PIN prog_clk_1_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END prog_clk_1_W_in
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 10.240 100.000 10.840 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 2.080 100.000 2.680 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 97.600 8.880 100.000 9.480 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 97.600 0.720 100.000 1.320 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END prog_clk_3_W_out
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.375 10.640 35.975 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.075 73.525 ;
      LAYER met1 ;
        RECT 1.910 5.140 97.450 82.920 ;
      LAYER met2 ;
        RECT 1.940 82.320 8.090 84.165 ;
        RECT 8.930 82.320 24.650 84.165 ;
        RECT 25.490 82.320 41.210 84.165 ;
        RECT 42.050 82.320 57.770 84.165 ;
        RECT 58.610 82.320 74.330 84.165 ;
        RECT 75.170 82.320 90.890 84.165 ;
        RECT 91.730 82.320 97.420 84.165 ;
        RECT 1.940 2.680 97.420 82.320 ;
        RECT 2.490 0.835 5.790 2.680 ;
        RECT 6.630 0.835 10.390 2.680 ;
        RECT 11.230 0.835 14.990 2.680 ;
        RECT 15.830 0.835 19.590 2.680 ;
        RECT 20.430 0.835 24.190 2.680 ;
        RECT 25.030 0.835 28.790 2.680 ;
        RECT 29.630 0.835 33.390 2.680 ;
        RECT 34.230 0.835 37.530 2.680 ;
        RECT 38.370 0.835 42.130 2.680 ;
        RECT 42.970 0.835 46.730 2.680 ;
        RECT 47.570 0.835 51.330 2.680 ;
        RECT 52.170 0.835 55.930 2.680 ;
        RECT 56.770 0.835 60.530 2.680 ;
        RECT 61.370 0.835 65.130 2.680 ;
        RECT 65.970 0.835 69.270 2.680 ;
        RECT 70.110 0.835 73.870 2.680 ;
        RECT 74.710 0.835 78.470 2.680 ;
        RECT 79.310 0.835 83.070 2.680 ;
        RECT 83.910 0.835 87.670 2.680 ;
        RECT 88.510 0.835 92.270 2.680 ;
        RECT 93.110 0.835 96.870 2.680 ;
      LAYER met3 ;
        RECT 2.800 81.920 97.200 84.145 ;
        RECT 2.400 81.280 97.600 81.920 ;
        RECT 2.800 78.520 97.200 81.280 ;
        RECT 2.400 77.880 97.600 78.520 ;
        RECT 2.800 75.120 97.200 77.880 ;
        RECT 2.400 74.480 97.200 75.120 ;
        RECT 2.800 73.760 97.200 74.480 ;
        RECT 2.800 73.120 97.600 73.760 ;
        RECT 2.800 71.720 97.200 73.120 ;
        RECT 2.400 71.080 97.200 71.720 ;
        RECT 2.800 70.360 97.200 71.080 ;
        RECT 2.800 69.720 97.600 70.360 ;
        RECT 2.800 68.320 97.200 69.720 ;
        RECT 2.400 67.680 97.200 68.320 ;
        RECT 2.800 65.600 97.200 67.680 ;
        RECT 2.800 64.960 97.600 65.600 ;
        RECT 2.800 64.920 97.200 64.960 ;
        RECT 2.400 64.280 97.200 64.920 ;
        RECT 2.800 62.200 97.200 64.280 ;
        RECT 2.800 61.560 97.600 62.200 ;
        RECT 2.800 61.520 97.200 61.560 ;
        RECT 2.400 60.880 97.200 61.520 ;
        RECT 2.800 58.120 97.200 60.880 ;
        RECT 2.400 57.480 97.200 58.120 ;
        RECT 2.800 57.440 97.200 57.480 ;
        RECT 2.800 56.800 97.600 57.440 ;
        RECT 2.800 54.720 97.200 56.800 ;
        RECT 2.400 54.080 97.200 54.720 ;
        RECT 2.800 54.040 97.200 54.080 ;
        RECT 2.800 53.400 97.600 54.040 ;
        RECT 2.800 51.320 97.200 53.400 ;
        RECT 2.400 50.680 97.200 51.320 ;
        RECT 2.800 49.280 97.200 50.680 ;
        RECT 2.800 48.640 97.600 49.280 ;
        RECT 2.800 47.920 97.200 48.640 ;
        RECT 2.400 47.280 97.200 47.920 ;
        RECT 2.800 45.880 97.200 47.280 ;
        RECT 2.800 45.240 97.600 45.880 ;
        RECT 2.800 44.520 97.200 45.240 ;
        RECT 2.400 43.880 97.200 44.520 ;
        RECT 2.800 41.120 97.200 43.880 ;
        RECT 2.400 40.480 97.600 41.120 ;
        RECT 2.800 37.720 97.200 40.480 ;
        RECT 2.400 37.080 97.600 37.720 ;
        RECT 2.800 34.320 97.200 37.080 ;
        RECT 2.400 33.680 97.200 34.320 ;
        RECT 2.800 32.960 97.200 33.680 ;
        RECT 2.800 32.320 97.600 32.960 ;
        RECT 2.800 30.920 97.200 32.320 ;
        RECT 2.400 30.280 97.200 30.920 ;
        RECT 2.800 29.560 97.200 30.280 ;
        RECT 2.800 28.920 97.600 29.560 ;
        RECT 2.800 27.520 97.200 28.920 ;
        RECT 2.400 26.880 97.200 27.520 ;
        RECT 2.800 24.800 97.200 26.880 ;
        RECT 2.800 24.160 97.600 24.800 ;
        RECT 2.800 24.120 97.200 24.160 ;
        RECT 2.400 23.480 97.200 24.120 ;
        RECT 2.800 21.400 97.200 23.480 ;
        RECT 2.800 20.760 97.600 21.400 ;
        RECT 2.800 20.720 97.200 20.760 ;
        RECT 2.400 20.080 97.200 20.720 ;
        RECT 2.800 17.320 97.200 20.080 ;
        RECT 2.400 16.680 97.200 17.320 ;
        RECT 2.800 16.640 97.200 16.680 ;
        RECT 2.800 16.000 97.600 16.640 ;
        RECT 2.800 13.920 97.200 16.000 ;
        RECT 2.400 13.280 97.200 13.920 ;
        RECT 2.800 13.240 97.200 13.280 ;
        RECT 2.800 12.600 97.600 13.240 ;
        RECT 2.800 10.520 97.200 12.600 ;
        RECT 2.400 9.880 97.200 10.520 ;
        RECT 2.800 8.480 97.200 9.880 ;
        RECT 2.800 7.840 97.600 8.480 ;
        RECT 2.800 7.120 97.200 7.840 ;
        RECT 2.400 6.480 97.200 7.120 ;
        RECT 2.800 5.080 97.200 6.480 ;
        RECT 2.800 4.440 97.600 5.080 ;
        RECT 2.800 3.720 97.200 4.440 ;
        RECT 2.400 3.080 97.200 3.720 ;
        RECT 2.800 0.855 97.200 3.080 ;
      LAYER met4 ;
        RECT 15.015 10.640 19.145 73.680 ;
        RECT 21.545 10.640 33.975 73.680 ;
        RECT 36.375 10.640 81.585 73.680 ;
  END
END cbx_1__1_
END LIBRARY

