magic
tech sky130A
magscale 1 2
timestamp 1608762747
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 3893 15487 3927 15589
rect 19073 15419 19107 15521
rect 12081 14399 12115 14501
rect 8033 13719 8067 13889
rect 9505 11067 9539 11169
rect 10517 10999 10551 11101
rect 8861 9367 8895 9537
rect 8861 4471 8895 4709
rect 9447 4233 9505 4267
rect 15577 3927 15611 4029
rect 9447 3893 9505 3927
<< viali >>
rect 2053 20009 2087 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 1869 19873 1903 19907
rect 2421 19873 2455 19907
rect 15853 19873 15887 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 15945 19805 15979 19839
rect 16037 19805 16071 19839
rect 2605 19737 2639 19771
rect 15485 19669 15519 19703
rect 20729 19669 20763 19703
rect 2053 19465 2087 19499
rect 5365 19465 5399 19499
rect 15853 19465 15887 19499
rect 19625 19465 19659 19499
rect 20177 19465 20211 19499
rect 7757 19329 7791 19363
rect 1869 19261 1903 19295
rect 2421 19261 2455 19295
rect 3157 19261 3191 19295
rect 5181 19261 5215 19295
rect 5733 19261 5767 19295
rect 8493 19261 8527 19295
rect 10149 19261 10183 19295
rect 12449 19261 12483 19295
rect 14473 19261 14507 19295
rect 18889 19261 18923 19295
rect 19441 19261 19475 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 3424 19193 3458 19227
rect 6009 19193 6043 19227
rect 7481 19193 7515 19227
rect 8738 19193 8772 19227
rect 10394 19193 10428 19227
rect 12716 19193 12750 19227
rect 14740 19193 14774 19227
rect 2605 19125 2639 19159
rect 4537 19125 4571 19159
rect 7113 19125 7147 19159
rect 7573 19125 7607 19159
rect 9873 19125 9907 19159
rect 11529 19125 11563 19159
rect 13829 19125 13863 19159
rect 19073 19125 19107 19159
rect 20729 19125 20763 19159
rect 1961 18921 1995 18955
rect 2513 18921 2547 18955
rect 3065 18921 3099 18955
rect 8033 18921 8067 18955
rect 13093 18921 13127 18955
rect 14473 18921 14507 18955
rect 19533 18921 19567 18955
rect 8769 18853 8803 18887
rect 14565 18853 14599 18887
rect 16028 18853 16062 18887
rect 20177 18853 20211 18887
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2881 18785 2915 18819
rect 4988 18785 5022 18819
rect 6920 18785 6954 18819
rect 8861 18785 8895 18819
rect 11244 18785 11278 18819
rect 12633 18785 12667 18819
rect 13461 18785 13495 18819
rect 15761 18785 15795 18819
rect 19349 18785 19383 18819
rect 19901 18785 19935 18819
rect 4721 18717 4755 18751
rect 6653 18717 6687 18751
rect 8953 18717 8987 18751
rect 10977 18717 11011 18751
rect 13553 18717 13587 18751
rect 13737 18717 13771 18751
rect 14749 18717 14783 18751
rect 12357 18649 12391 18683
rect 14105 18649 14139 18683
rect 6101 18581 6135 18615
rect 8401 18581 8435 18615
rect 17141 18581 17175 18615
rect 7021 18377 7055 18411
rect 10333 18377 10367 18411
rect 1961 18309 1995 18343
rect 13277 18309 13311 18343
rect 20177 18309 20211 18343
rect 3249 18241 3283 18275
rect 7481 18241 7515 18275
rect 7573 18241 7607 18275
rect 8033 18241 8067 18275
rect 8677 18241 8711 18275
rect 10885 18241 10919 18275
rect 13921 18241 13955 18275
rect 15669 18241 15703 18275
rect 16681 18241 16715 18275
rect 1777 18173 1811 18207
rect 3617 18173 3651 18207
rect 3884 18173 3918 18207
rect 7389 18173 7423 18207
rect 16589 18173 16623 18207
rect 18245 18173 18279 18207
rect 18521 18173 18555 18207
rect 19165 18173 19199 18207
rect 19993 18173 20027 18207
rect 20545 18173 20579 18207
rect 8922 18105 8956 18139
rect 10701 18105 10735 18139
rect 13645 18105 13679 18139
rect 2605 18037 2639 18071
rect 2973 18037 3007 18071
rect 3065 18037 3099 18071
rect 4997 18037 5031 18071
rect 10057 18037 10091 18071
rect 10793 18037 10827 18071
rect 13737 18037 13771 18071
rect 15117 18037 15151 18071
rect 15485 18037 15519 18071
rect 15577 18037 15611 18071
rect 16129 18037 16163 18071
rect 16497 18037 16531 18071
rect 19349 18037 19383 18071
rect 20729 18037 20763 18071
rect 1593 17833 1627 17867
rect 2329 17833 2363 17867
rect 2973 17833 3007 17867
rect 9689 17833 9723 17867
rect 12541 17833 12575 17867
rect 13645 17833 13679 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 6929 17765 6963 17799
rect 14013 17765 14047 17799
rect 15669 17765 15703 17799
rect 16856 17765 16890 17799
rect 19993 17765 20027 17799
rect 1409 17697 1443 17731
rect 3341 17697 3375 17731
rect 4721 17697 4755 17731
rect 6653 17697 6687 17731
rect 10057 17697 10091 17731
rect 10149 17697 10183 17731
rect 12449 17697 12483 17731
rect 19717 17697 19751 17731
rect 2421 17629 2455 17663
rect 2605 17629 2639 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 4813 17629 4847 17663
rect 4905 17629 4939 17663
rect 10241 17629 10275 17663
rect 12725 17629 12759 17663
rect 14105 17629 14139 17663
rect 14197 17629 14231 17663
rect 15853 17629 15887 17663
rect 16589 17629 16623 17663
rect 4353 17561 4387 17595
rect 12081 17561 12115 17595
rect 1961 17493 1995 17527
rect 17969 17493 18003 17527
rect 3065 17289 3099 17323
rect 4813 17289 4847 17323
rect 6837 17289 6871 17323
rect 8033 17289 8067 17323
rect 16037 17289 16071 17323
rect 20177 17289 20211 17323
rect 2237 17153 2271 17187
rect 3709 17153 3743 17187
rect 5457 17153 5491 17187
rect 7389 17153 7423 17187
rect 8677 17153 8711 17187
rect 13921 17153 13955 17187
rect 16589 17153 16623 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 3433 17085 3467 17119
rect 10701 17085 10735 17119
rect 13737 17085 13771 17119
rect 18153 17085 18187 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 7297 17017 7331 17051
rect 8401 17017 8435 17051
rect 10968 17017 11002 17051
rect 16405 17017 16439 17051
rect 18420 17017 18454 17051
rect 1685 16949 1719 16983
rect 3525 16949 3559 16983
rect 5181 16949 5215 16983
rect 5273 16949 5307 16983
rect 7205 16949 7239 16983
rect 8493 16949 8527 16983
rect 12081 16949 12115 16983
rect 13369 16949 13403 16983
rect 13829 16949 13863 16983
rect 16497 16949 16531 16983
rect 19533 16949 19567 16983
rect 20729 16949 20763 16983
rect 2513 16745 2547 16779
rect 3065 16745 3099 16779
rect 3433 16745 3467 16779
rect 9045 16745 9079 16779
rect 15301 16745 15335 16779
rect 15761 16745 15795 16779
rect 16313 16745 16347 16779
rect 19901 16745 19935 16779
rect 11897 16677 11931 16711
rect 12970 16677 13004 16711
rect 16773 16677 16807 16711
rect 1777 16609 1811 16643
rect 2329 16609 2363 16643
rect 2881 16609 2915 16643
rect 5089 16609 5123 16643
rect 5356 16609 5390 16643
rect 7665 16609 7699 16643
rect 7932 16609 7966 16643
rect 15669 16609 15703 16643
rect 16681 16609 16715 16643
rect 19717 16609 19751 16643
rect 20269 16609 20303 16643
rect 11989 16541 12023 16575
rect 12081 16541 12115 16575
rect 12725 16541 12759 16575
rect 15945 16541 15979 16575
rect 16957 16541 16991 16575
rect 1961 16473 1995 16507
rect 6469 16405 6503 16439
rect 11529 16405 11563 16439
rect 14105 16405 14139 16439
rect 20453 16405 20487 16439
rect 4997 16201 5031 16235
rect 6837 16201 6871 16235
rect 9873 16201 9907 16235
rect 10333 16201 10367 16235
rect 19441 16201 19475 16235
rect 2329 16065 2363 16099
rect 5549 16065 5583 16099
rect 7389 16065 7423 16099
rect 10793 16065 10827 16099
rect 10977 16065 11011 16099
rect 11897 16065 11931 16099
rect 12449 16065 12483 16099
rect 13921 16065 13955 16099
rect 19993 16065 20027 16099
rect 2053 15997 2087 16031
rect 8493 15997 8527 16031
rect 11805 15997 11839 16031
rect 18061 15997 18095 16031
rect 19809 15997 19843 16031
rect 20545 15997 20579 16031
rect 5457 15929 5491 15963
rect 7205 15929 7239 15963
rect 8760 15929 8794 15963
rect 11713 15929 11747 15963
rect 14166 15929 14200 15963
rect 18306 15929 18340 15963
rect 20821 15929 20855 15963
rect 5365 15861 5399 15895
rect 7297 15861 7331 15895
rect 10701 15861 10735 15895
rect 11345 15861 11379 15895
rect 15301 15861 15335 15895
rect 1961 15657 1995 15691
rect 5457 15657 5491 15691
rect 8585 15657 8619 15691
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 11805 15657 11839 15691
rect 13461 15657 13495 15691
rect 13921 15657 13955 15691
rect 17233 15657 17267 15691
rect 2596 15589 2630 15623
rect 3893 15589 3927 15623
rect 6092 15589 6126 15623
rect 10057 15589 10091 15623
rect 11897 15589 11931 15623
rect 19625 15589 19659 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 4333 15521 4367 15555
rect 5825 15521 5859 15555
rect 8033 15521 8067 15555
rect 8953 15521 8987 15555
rect 13829 15521 13863 15555
rect 15853 15521 15887 15555
rect 16120 15521 16154 15555
rect 18613 15521 18647 15555
rect 18705 15521 18739 15555
rect 19073 15521 19107 15555
rect 20269 15521 20303 15555
rect 3893 15453 3927 15487
rect 4077 15453 4111 15487
rect 9229 15453 9263 15487
rect 10241 15453 10275 15487
rect 12081 15453 12115 15487
rect 14105 15453 14139 15487
rect 18797 15453 18831 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 11437 15385 11471 15419
rect 19073 15385 19107 15419
rect 3709 15317 3743 15351
rect 7205 15317 7239 15351
rect 7849 15317 7883 15351
rect 18245 15317 18279 15351
rect 19257 15317 19291 15351
rect 20453 15317 20487 15351
rect 1961 15113 1995 15147
rect 8677 15113 8711 15147
rect 16957 15113 16991 15147
rect 18889 15113 18923 15147
rect 3525 14977 3559 15011
rect 7021 14977 7055 15011
rect 9321 14977 9355 15011
rect 17509 14977 17543 15011
rect 18429 14977 18463 15011
rect 19441 14977 19475 15011
rect 1777 14909 1811 14943
rect 7288 14909 7322 14943
rect 12817 14909 12851 14943
rect 13461 14909 13495 14943
rect 15117 14909 15151 14943
rect 17325 14909 17359 14943
rect 19257 14909 19291 14943
rect 19993 14909 20027 14943
rect 20729 14909 20763 14943
rect 3792 14841 3826 14875
rect 9045 14841 9079 14875
rect 13728 14841 13762 14875
rect 15362 14841 15396 14875
rect 20269 14841 20303 14875
rect 4905 14773 4939 14807
rect 8401 14773 8435 14807
rect 9137 14773 9171 14807
rect 12633 14773 12667 14807
rect 14841 14773 14875 14807
rect 16497 14773 16531 14807
rect 17417 14773 17451 14807
rect 19349 14773 19383 14807
rect 20913 14773 20947 14807
rect 7021 14569 7055 14603
rect 14933 14569 14967 14603
rect 17601 14569 17635 14603
rect 18153 14569 18187 14603
rect 19901 14569 19935 14603
rect 5632 14501 5666 14535
rect 12081 14501 12115 14535
rect 1777 14433 1811 14467
rect 2973 14433 3007 14467
rect 5365 14433 5399 14467
rect 7389 14433 7423 14467
rect 10609 14433 10643 14467
rect 10876 14433 10910 14467
rect 12532 14433 12566 14467
rect 14289 14433 14323 14467
rect 15117 14433 15151 14467
rect 17509 14433 17543 14467
rect 18521 14433 18555 14467
rect 19717 14433 19751 14467
rect 20269 14433 20303 14467
rect 3065 14365 3099 14399
rect 3249 14365 3283 14399
rect 7481 14365 7515 14399
rect 7573 14365 7607 14399
rect 9137 14365 9171 14399
rect 12081 14365 12115 14399
rect 12265 14365 12299 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 17693 14365 17727 14399
rect 18613 14365 18647 14399
rect 18705 14365 18739 14399
rect 11989 14297 12023 14331
rect 13645 14297 13679 14331
rect 17141 14297 17175 14331
rect 1961 14229 1995 14263
rect 2605 14229 2639 14263
rect 6745 14229 6779 14263
rect 13921 14229 13955 14263
rect 20453 14229 20487 14263
rect 2145 14025 2179 14059
rect 3893 14025 3927 14059
rect 6009 14025 6043 14059
rect 6837 14025 6871 14059
rect 8125 14025 8159 14059
rect 9137 14025 9171 14059
rect 10149 14025 10183 14059
rect 14289 14025 14323 14059
rect 18797 14025 18831 14059
rect 3341 13957 3375 13991
rect 11253 13957 11287 13991
rect 21005 13957 21039 13991
rect 1685 13889 1719 13923
rect 2697 13889 2731 13923
rect 4445 13889 4479 13923
rect 7481 13889 7515 13923
rect 8033 13889 8067 13923
rect 8769 13889 8803 13923
rect 9781 13889 9815 13923
rect 10701 13889 10735 13923
rect 11897 13889 11931 13923
rect 13921 13889 13955 13923
rect 14749 13889 14783 13923
rect 14933 13889 14967 13923
rect 19349 13889 19383 13923
rect 1409 13821 1443 13855
rect 3157 13821 3191 13855
rect 6193 13821 6227 13855
rect 9505 13821 9539 13855
rect 15301 13821 15335 13855
rect 15568 13821 15602 13855
rect 20085 13821 20119 13855
rect 20361 13821 20395 13855
rect 20821 13821 20855 13855
rect 8493 13753 8527 13787
rect 8585 13753 8619 13787
rect 10517 13753 10551 13787
rect 10609 13753 10643 13787
rect 14657 13753 14691 13787
rect 2513 13685 2547 13719
rect 2605 13685 2639 13719
rect 4261 13685 4295 13719
rect 4353 13685 4387 13719
rect 7205 13685 7239 13719
rect 7297 13685 7331 13719
rect 8033 13685 8067 13719
rect 9597 13685 9631 13719
rect 11621 13685 11655 13719
rect 11713 13685 11747 13719
rect 13277 13685 13311 13719
rect 13645 13685 13679 13719
rect 13737 13685 13771 13719
rect 16681 13685 16715 13719
rect 19165 13685 19199 13719
rect 19257 13685 19291 13719
rect 2237 13481 2271 13515
rect 4537 13481 4571 13515
rect 7297 13481 7331 13515
rect 7757 13481 7791 13515
rect 9965 13481 9999 13515
rect 13185 13481 13219 13515
rect 13829 13481 13863 13515
rect 15853 13481 15887 13515
rect 16497 13481 16531 13515
rect 17693 13481 17727 13515
rect 18705 13481 18739 13515
rect 16865 13413 16899 13447
rect 2605 13345 2639 13379
rect 3249 13345 3283 13379
rect 4905 13345 4939 13379
rect 7665 13345 7699 13379
rect 10333 13345 10367 13379
rect 18061 13345 18095 13379
rect 19073 13345 19107 13379
rect 2697 13277 2731 13311
rect 2881 13277 2915 13311
rect 4997 13277 5031 13311
rect 5089 13277 5123 13311
rect 7849 13277 7883 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 13277 13277 13311 13311
rect 13461 13277 13495 13311
rect 15945 13277 15979 13311
rect 16129 13277 16163 13311
rect 16957 13277 16991 13311
rect 17141 13277 17175 13311
rect 18153 13277 18187 13311
rect 18245 13277 18279 13311
rect 19165 13277 19199 13311
rect 19257 13277 19291 13311
rect 15485 13209 15519 13243
rect 12817 13141 12851 13175
rect 2421 12937 2455 12971
rect 4997 12937 5031 12971
rect 7113 12937 7147 12971
rect 8401 12937 8435 12971
rect 12449 12937 12483 12971
rect 16497 12937 16531 12971
rect 18337 12937 18371 12971
rect 7389 12869 7423 12903
rect 14289 12869 14323 12903
rect 15301 12869 15335 12903
rect 3065 12801 3099 12835
rect 5457 12801 5491 12835
rect 5641 12801 5675 12835
rect 7941 12801 7975 12835
rect 8861 12801 8895 12835
rect 8953 12801 8987 12835
rect 13093 12801 13127 12835
rect 14933 12801 14967 12835
rect 15945 12801 15979 12835
rect 17141 12801 17175 12835
rect 18981 12801 19015 12835
rect 20821 12801 20855 12835
rect 2789 12733 2823 12767
rect 5365 12733 5399 12767
rect 7297 12733 7331 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 13829 12733 13863 12767
rect 15669 12733 15703 12767
rect 16865 12733 16899 12767
rect 20729 12733 20763 12767
rect 12909 12665 12943 12699
rect 14657 12665 14691 12699
rect 16957 12665 16991 12699
rect 20637 12665 20671 12699
rect 2881 12597 2915 12631
rect 8769 12597 8803 12631
rect 11345 12597 11379 12631
rect 12817 12597 12851 12631
rect 13645 12597 13679 12631
rect 14749 12597 14783 12631
rect 15761 12597 15795 12631
rect 18705 12597 18739 12631
rect 18797 12597 18831 12631
rect 20269 12597 20303 12631
rect 2237 12393 2271 12427
rect 7573 12393 7607 12427
rect 11161 12393 11195 12427
rect 12449 12393 12483 12427
rect 15301 12393 15335 12427
rect 18153 12393 18187 12427
rect 18521 12393 18555 12427
rect 2605 12257 2639 12291
rect 5181 12257 5215 12291
rect 5273 12257 5307 12291
rect 6193 12257 6227 12291
rect 7941 12257 7975 12291
rect 9689 12257 9723 12291
rect 9945 12257 9979 12291
rect 11529 12257 11563 12291
rect 12357 12257 12391 12291
rect 13452 12257 13486 12291
rect 15669 12257 15703 12291
rect 19432 12257 19466 12291
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 5365 12189 5399 12223
rect 6285 12189 6319 12223
rect 6377 12189 6411 12223
rect 7113 12189 7147 12223
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 11621 12189 11655 12223
rect 11713 12189 11747 12223
rect 12541 12189 12575 12223
rect 13185 12189 13219 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 18613 12189 18647 12223
rect 18705 12189 18739 12223
rect 19165 12189 19199 12223
rect 11069 12121 11103 12155
rect 11989 12121 12023 12155
rect 4813 12053 4847 12087
rect 5825 12053 5859 12087
rect 14565 12053 14599 12087
rect 20545 12053 20579 12087
rect 4353 11849 4387 11883
rect 5549 11849 5583 11883
rect 7113 11849 7147 11883
rect 11529 11849 11563 11883
rect 13829 11849 13863 11883
rect 20361 11849 20395 11883
rect 3709 11781 3743 11815
rect 8493 11781 8527 11815
rect 9873 11781 9907 11815
rect 2329 11713 2363 11747
rect 4813 11713 4847 11747
rect 4905 11713 4939 11747
rect 6101 11713 6135 11747
rect 7757 11713 7791 11747
rect 9137 11713 9171 11747
rect 10517 11713 10551 11747
rect 12081 11713 12115 11747
rect 15945 11713 15979 11747
rect 18981 11713 19015 11747
rect 2596 11645 2630 11679
rect 4721 11645 4755 11679
rect 5917 11645 5951 11679
rect 7481 11645 7515 11679
rect 10333 11645 10367 11679
rect 11897 11645 11931 11679
rect 12456 11645 12490 11679
rect 15761 11645 15795 11679
rect 11345 11577 11379 11611
rect 11989 11577 12023 11611
rect 12716 11577 12750 11611
rect 19248 11577 19282 11611
rect 6009 11509 6043 11543
rect 7573 11509 7607 11543
rect 8861 11509 8895 11543
rect 8953 11509 8987 11543
rect 10241 11509 10275 11543
rect 15393 11509 15427 11543
rect 15853 11509 15887 11543
rect 18061 11509 18095 11543
rect 2513 11305 2547 11339
rect 5181 11305 5215 11339
rect 6009 11305 6043 11339
rect 8033 11305 8067 11339
rect 12449 11305 12483 11339
rect 12909 11305 12943 11339
rect 13461 11305 13495 11339
rect 15301 11305 15335 11339
rect 18889 11305 18923 11339
rect 2881 11237 2915 11271
rect 12817 11237 12851 11271
rect 1777 11169 1811 11203
rect 5273 11169 5307 11203
rect 6377 11169 6411 11203
rect 8217 11169 8251 11203
rect 9505 11169 9539 11203
rect 10609 11169 10643 11203
rect 13645 11169 13679 11203
rect 15669 11169 15703 11203
rect 17500 11169 17534 11203
rect 19257 11169 19291 11203
rect 2973 11101 3007 11135
rect 3065 11101 3099 11135
rect 5457 11101 5491 11135
rect 6469 11101 6503 11135
rect 6561 11101 6595 11135
rect 1961 11033 1995 11067
rect 9505 11033 9539 11067
rect 10517 11101 10551 11135
rect 13001 11101 13035 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 17233 11101 17267 11135
rect 19349 11101 19383 11135
rect 19441 11101 19475 11135
rect 11897 11033 11931 11067
rect 18613 11033 18647 11067
rect 4813 10965 4847 10999
rect 10517 10965 10551 10999
rect 2513 10761 2547 10795
rect 5733 10761 5767 10795
rect 6837 10761 6871 10795
rect 14013 10761 14047 10795
rect 18061 10761 18095 10795
rect 16957 10693 16991 10727
rect 1961 10625 1995 10659
rect 3065 10625 3099 10659
rect 4353 10625 4387 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 14565 10625 14599 10659
rect 15485 10625 15519 10659
rect 15577 10625 15611 10659
rect 17509 10625 17543 10659
rect 18613 10625 18647 10659
rect 20177 10625 20211 10659
rect 20361 10625 20395 10659
rect 1777 10557 1811 10591
rect 10241 10557 10275 10591
rect 10508 10557 10542 10591
rect 17417 10557 17451 10591
rect 18429 10557 18463 10591
rect 18521 10557 18555 10591
rect 2881 10489 2915 10523
rect 4620 10489 4654 10523
rect 14381 10489 14415 10523
rect 15393 10489 15427 10523
rect 16037 10489 16071 10523
rect 2973 10421 3007 10455
rect 7205 10421 7239 10455
rect 7849 10421 7883 10455
rect 11621 10421 11655 10455
rect 14473 10421 14507 10455
rect 15025 10421 15059 10455
rect 17325 10421 17359 10455
rect 19717 10421 19751 10455
rect 20085 10421 20119 10455
rect 1961 10217 1995 10251
rect 5457 10217 5491 10251
rect 6285 10217 6319 10251
rect 6653 10217 6687 10251
rect 10149 10217 10183 10251
rect 10701 10217 10735 10251
rect 15301 10217 15335 10251
rect 18245 10217 18279 10251
rect 19993 10217 20027 10251
rect 20913 10217 20947 10251
rect 1777 10081 1811 10115
rect 4344 10081 4378 10115
rect 6745 10081 6779 10115
rect 7553 10081 7587 10115
rect 10057 10081 10091 10115
rect 11704 10081 11738 10115
rect 13349 10081 13383 10115
rect 15669 10081 15703 10115
rect 17132 10081 17166 10115
rect 20085 10081 20119 10115
rect 4077 10013 4111 10047
rect 6929 10013 6963 10047
rect 7297 10013 7331 10047
rect 10241 10013 10275 10047
rect 11437 10013 11471 10047
rect 13093 10013 13127 10047
rect 15761 10013 15795 10047
rect 15853 10013 15887 10047
rect 16865 10013 16899 10047
rect 20177 10013 20211 10047
rect 14473 9945 14507 9979
rect 8677 9877 8711 9911
rect 9689 9877 9723 9911
rect 12817 9877 12851 9911
rect 19625 9877 19659 9911
rect 10333 9673 10367 9707
rect 15669 9673 15703 9707
rect 5733 9605 5767 9639
rect 12541 9605 12575 9639
rect 15393 9605 15427 9639
rect 1961 9537 1995 9571
rect 6377 9537 6411 9571
rect 7573 9537 7607 9571
rect 8861 9537 8895 9571
rect 8953 9537 8987 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 13185 9537 13219 9571
rect 14020 9537 14054 9571
rect 16221 9537 16255 9571
rect 1777 9469 1811 9503
rect 2789 9469 2823 9503
rect 7389 9469 7423 9503
rect 7481 9469 7515 9503
rect 8217 9469 8251 9503
rect 3056 9401 3090 9435
rect 6101 9401 6135 9435
rect 9220 9469 9254 9503
rect 13001 9469 13035 9503
rect 13921 9469 13955 9503
rect 14280 9469 14314 9503
rect 19625 9469 19659 9503
rect 19892 9469 19926 9503
rect 12909 9401 12943 9435
rect 16037 9401 16071 9435
rect 4169 9333 4203 9367
rect 6193 9333 6227 9367
rect 7021 9333 7055 9367
rect 8033 9333 8067 9367
rect 8861 9333 8895 9367
rect 10609 9333 10643 9367
rect 10977 9333 11011 9367
rect 13737 9333 13771 9367
rect 16129 9333 16163 9367
rect 21005 9333 21039 9367
rect 4537 9129 4571 9163
rect 7205 9129 7239 9163
rect 8677 9129 8711 9163
rect 11253 9129 11287 9163
rect 13093 9129 13127 9163
rect 18245 9129 18279 9163
rect 19625 9129 19659 9163
rect 8585 9061 8619 9095
rect 19533 9061 19567 9095
rect 1685 8993 1719 9027
rect 1952 8993 1986 9027
rect 4445 8993 4479 9027
rect 5805 8993 5839 9027
rect 7573 8993 7607 9027
rect 11161 8993 11195 9027
rect 13001 8993 13035 9027
rect 17132 8993 17166 9027
rect 4721 8925 4755 8959
rect 5549 8925 5583 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 8861 8925 8895 8959
rect 11437 8925 11471 8959
rect 13277 8925 13311 8959
rect 16865 8925 16899 8959
rect 19809 8925 19843 8959
rect 6929 8857 6963 8891
rect 8217 8857 8251 8891
rect 3065 8789 3099 8823
rect 4077 8789 4111 8823
rect 10793 8789 10827 8823
rect 12633 8789 12667 8823
rect 19165 8789 19199 8823
rect 5641 8585 5675 8619
rect 6837 8585 6871 8619
rect 9505 8585 9539 8619
rect 13829 8517 13863 8551
rect 16957 8517 16991 8551
rect 18061 8517 18095 8551
rect 2973 8449 3007 8483
rect 7389 8449 7423 8483
rect 8125 8449 8159 8483
rect 17509 8449 17543 8483
rect 18613 8449 18647 8483
rect 2789 8381 2823 8415
rect 4261 8381 4295 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 12449 8381 12483 8415
rect 12716 8381 12750 8415
rect 15853 8381 15887 8415
rect 17325 8381 17359 8415
rect 18521 8381 18555 8415
rect 19257 8381 19291 8415
rect 19524 8381 19558 8415
rect 2697 8313 2731 8347
rect 4506 8313 4540 8347
rect 8392 8313 8426 8347
rect 2329 8245 2363 8279
rect 15669 8245 15703 8279
rect 17417 8245 17451 8279
rect 18429 8245 18463 8279
rect 20637 8245 20671 8279
rect 1409 8041 1443 8075
rect 1869 8041 1903 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 6653 8041 6687 8075
rect 8125 8041 8159 8075
rect 10149 8041 10183 8075
rect 12357 8041 12391 8075
rect 12633 8041 12667 8075
rect 17049 8041 17083 8075
rect 17509 8041 17543 8075
rect 18061 8041 18095 8075
rect 20177 8041 20211 8075
rect 2789 7973 2823 8007
rect 13001 7973 13035 8007
rect 14013 7973 14047 8007
rect 14105 7973 14139 8007
rect 15568 7973 15602 8007
rect 20085 7973 20119 8007
rect 1777 7905 1811 7939
rect 5825 7905 5859 7939
rect 6561 7905 6595 7939
rect 7021 7905 7055 7939
rect 8309 7905 8343 7939
rect 10057 7905 10091 7939
rect 12541 7905 12575 7939
rect 17417 7905 17451 7939
rect 2053 7837 2087 7871
rect 2881 7837 2915 7871
rect 2973 7837 3007 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 10241 7837 10275 7871
rect 10609 7837 10643 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 14197 7837 14231 7871
rect 15301 7837 15335 7871
rect 17601 7837 17635 7871
rect 20361 7837 20395 7871
rect 2421 7701 2455 7735
rect 5641 7701 5675 7735
rect 9689 7701 9723 7735
rect 13645 7701 13679 7735
rect 16681 7701 16715 7735
rect 19717 7701 19751 7735
rect 2237 7497 2271 7531
rect 8677 7497 8711 7531
rect 17601 7497 17635 7531
rect 5733 7429 5767 7463
rect 2697 7361 2731 7395
rect 2881 7361 2915 7395
rect 3249 7361 3283 7395
rect 6377 7361 6411 7395
rect 9321 7361 9355 7395
rect 12817 7361 12851 7395
rect 2605 7293 2639 7327
rect 9137 7293 9171 7327
rect 9689 7293 9723 7327
rect 13277 7293 13311 7327
rect 13544 7293 13578 7327
rect 16221 7293 16255 7327
rect 16488 7293 16522 7327
rect 19349 7293 19383 7327
rect 19616 7293 19650 7327
rect 6101 7225 6135 7259
rect 9956 7225 9990 7259
rect 6193 7157 6227 7191
rect 9045 7157 9079 7191
rect 11069 7157 11103 7191
rect 14657 7157 14691 7191
rect 20729 7157 20763 7191
rect 5825 6953 5859 6987
rect 6193 6953 6227 6987
rect 8217 6953 8251 6987
rect 12909 6953 12943 6987
rect 13001 6953 13035 6987
rect 2513 6885 2547 6919
rect 2973 6885 3007 6919
rect 6285 6817 6319 6851
rect 10609 6817 10643 6851
rect 10876 6817 10910 6851
rect 15301 6817 15335 6851
rect 15568 6817 15602 6851
rect 19165 6817 19199 6851
rect 19432 6817 19466 6851
rect 1869 6749 1903 6783
rect 3065 6749 3099 6783
rect 3157 6749 3191 6783
rect 6469 6749 6503 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 13185 6749 13219 6783
rect 17049 6749 17083 6783
rect 18705 6749 18739 6783
rect 2605 6613 2639 6647
rect 7849 6613 7883 6647
rect 11989 6613 12023 6647
rect 12541 6613 12575 6647
rect 16681 6613 16715 6647
rect 20545 6613 20579 6647
rect 5273 6409 5307 6443
rect 8493 6409 8527 6443
rect 9413 6409 9447 6443
rect 10425 6409 10459 6443
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 5733 6273 5767 6307
rect 5917 6273 5951 6307
rect 7113 6273 7147 6307
rect 10057 6273 10091 6307
rect 11069 6273 11103 6307
rect 13553 6273 13587 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 17233 6273 17267 6307
rect 18613 6273 18647 6307
rect 19625 6273 19659 6307
rect 19717 6273 19751 6307
rect 20729 6273 20763 6307
rect 1961 6205 1995 6239
rect 2697 6205 2731 6239
rect 7369 6205 7403 6239
rect 13461 6205 13495 6239
rect 16957 6205 16991 6239
rect 17049 6205 17083 6239
rect 19533 6205 19567 6239
rect 20637 6205 20671 6239
rect 2942 6137 2976 6171
rect 5641 6137 5675 6171
rect 6285 6137 6319 6171
rect 13369 6137 13403 6171
rect 15485 6137 15519 6171
rect 18521 6137 18555 6171
rect 1593 6069 1627 6103
rect 4077 6069 4111 6103
rect 9781 6069 9815 6103
rect 9873 6069 9907 6103
rect 10793 6069 10827 6103
rect 10885 6069 10919 6103
rect 13001 6069 13035 6103
rect 14013 6069 14047 6103
rect 15117 6069 15151 6103
rect 16589 6069 16623 6103
rect 18061 6069 18095 6103
rect 18429 6069 18463 6103
rect 19165 6069 19199 6103
rect 20177 6069 20211 6103
rect 20545 6069 20579 6103
rect 5457 5865 5491 5899
rect 7113 5865 7147 5899
rect 7481 5865 7515 5899
rect 7941 5865 7975 5899
rect 8861 5865 8895 5899
rect 10149 5865 10183 5899
rect 13277 5865 13311 5899
rect 13369 5865 13403 5899
rect 14657 5865 14691 5899
rect 16221 5865 16255 5899
rect 19349 5865 19383 5899
rect 20085 5865 20119 5899
rect 4322 5797 4356 5831
rect 8953 5797 8987 5831
rect 14565 5797 14599 5831
rect 16313 5797 16347 5831
rect 19257 5797 19291 5831
rect 2605 5729 2639 5763
rect 6000 5729 6034 5763
rect 7849 5729 7883 5763
rect 10517 5729 10551 5763
rect 11253 5729 11287 5763
rect 11509 5729 11543 5763
rect 17489 5729 17523 5763
rect 2697 5661 2731 5695
rect 2789 5661 2823 5695
rect 4077 5661 4111 5695
rect 5733 5661 5767 5695
rect 8033 5661 8067 5695
rect 9045 5661 9079 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 13553 5661 13587 5695
rect 14841 5661 14875 5695
rect 16497 5661 16531 5695
rect 17233 5661 17267 5695
rect 19533 5661 19567 5695
rect 8493 5593 8527 5627
rect 12633 5593 12667 5627
rect 14197 5593 14231 5627
rect 18613 5593 18647 5627
rect 2237 5525 2271 5559
rect 12909 5525 12943 5559
rect 15853 5525 15887 5559
rect 18889 5525 18923 5559
rect 2421 5321 2455 5355
rect 7849 5321 7883 5355
rect 11253 5321 11287 5355
rect 3433 5253 3467 5287
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 2973 5185 3007 5219
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 8401 5185 8435 5219
rect 18797 5185 18831 5219
rect 1777 5117 1811 5151
rect 2789 5117 2823 5151
rect 9873 5117 9907 5151
rect 10140 5117 10174 5151
rect 12541 5117 12575 5151
rect 12808 5117 12842 5151
rect 14197 5117 14231 5151
rect 20545 5117 20579 5151
rect 3801 5049 3835 5083
rect 8217 5049 8251 5083
rect 14442 5049 14476 5083
rect 19042 5049 19076 5083
rect 1409 4981 1443 5015
rect 2881 4981 2915 5015
rect 8309 4981 8343 5015
rect 11529 4981 11563 5015
rect 13921 4981 13955 5015
rect 15577 4981 15611 5015
rect 20177 4981 20211 5015
rect 20729 4981 20763 5015
rect 2329 4777 2363 4811
rect 2789 4777 2823 4811
rect 10609 4777 10643 4811
rect 10977 4777 11011 4811
rect 13461 4777 13495 4811
rect 15853 4777 15887 4811
rect 18061 4777 18095 4811
rect 8861 4709 8895 4743
rect 13369 4709 13403 4743
rect 16948 4709 16982 4743
rect 2697 4641 2731 4675
rect 5365 4641 5399 4675
rect 5457 4641 5491 4675
rect 8309 4641 8343 4675
rect 2881 4573 2915 4607
rect 5641 4573 5675 4607
rect 8401 4573 8435 4607
rect 8585 4573 8619 4607
rect 15761 4641 15795 4675
rect 19165 4641 19199 4675
rect 19432 4641 19466 4675
rect 8953 4573 8987 4607
rect 11069 4573 11103 4607
rect 11161 4573 11195 4607
rect 13645 4573 13679 4607
rect 15945 4573 15979 4607
rect 16681 4573 16715 4607
rect 4997 4437 5031 4471
rect 7941 4437 7975 4471
rect 8861 4437 8895 4471
rect 13001 4437 13035 4471
rect 15393 4437 15427 4471
rect 20545 4437 20579 4471
rect 7573 4233 7607 4267
rect 8585 4233 8619 4267
rect 9413 4233 9447 4267
rect 9505 4233 9539 4267
rect 9597 4165 9631 4199
rect 4629 4097 4663 4131
rect 5089 4097 5123 4131
rect 6009 4097 6043 4131
rect 6193 4097 6227 4131
rect 8033 4097 8067 4131
rect 8217 4097 8251 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 10241 4097 10275 4131
rect 15301 4097 15335 4131
rect 19993 4097 20027 4131
rect 20177 4097 20211 4131
rect 1501 4029 1535 4063
rect 1768 4029 1802 4063
rect 4353 4029 4387 4063
rect 5917 4029 5951 4063
rect 8953 4029 8987 4063
rect 15117 4029 15151 4063
rect 15577 4029 15611 4063
rect 15669 4029 15703 4063
rect 15936 4029 15970 4063
rect 18981 4029 19015 4063
rect 19901 4029 19935 4063
rect 20545 4029 20579 4063
rect 2881 3893 2915 3927
rect 3985 3893 4019 3927
rect 4445 3893 4479 3927
rect 5549 3893 5583 3927
rect 7941 3893 7975 3927
rect 9413 3893 9447 3927
rect 9505 3893 9539 3927
rect 9965 3893 9999 3927
rect 10057 3893 10091 3927
rect 14657 3893 14691 3927
rect 15025 3893 15059 3927
rect 15577 3893 15611 3927
rect 17049 3893 17083 3927
rect 19165 3893 19199 3927
rect 19533 3893 19567 3927
rect 20729 3893 20763 3927
rect 4905 3689 4939 3723
rect 5549 3689 5583 3723
rect 10701 3689 10735 3723
rect 15669 3689 15703 3723
rect 16313 3689 16347 3723
rect 3341 3621 3375 3655
rect 4997 3621 5031 3655
rect 5917 3621 5951 3655
rect 7840 3621 7874 3655
rect 11989 3621 12023 3655
rect 15761 3621 15795 3655
rect 6009 3553 6043 3587
rect 7573 3553 7607 3587
rect 10609 3553 10643 3587
rect 11713 3553 11747 3587
rect 12449 3553 12483 3587
rect 13645 3553 13679 3587
rect 18061 3553 18095 3587
rect 18613 3553 18647 3587
rect 19257 3553 19291 3587
rect 19809 3553 19843 3587
rect 3433 3485 3467 3519
rect 3617 3485 3651 3519
rect 5089 3485 5123 3519
rect 6193 3485 6227 3519
rect 10885 3485 10919 3519
rect 12725 3485 12759 3519
rect 13921 3485 13955 3519
rect 15945 3485 15979 3519
rect 18245 3417 18279 3451
rect 2973 3349 3007 3383
rect 4537 3349 4571 3383
rect 8953 3349 8987 3383
rect 10241 3349 10275 3383
rect 15301 3349 15335 3383
rect 18797 3349 18831 3383
rect 19441 3349 19475 3383
rect 19993 3349 20027 3383
rect 2973 3145 3007 3179
rect 5365 3145 5399 3179
rect 8217 3009 8251 3043
rect 10517 3009 10551 3043
rect 10701 3009 10735 3043
rect 19717 3009 19751 3043
rect 1593 2941 1627 2975
rect 3985 2941 4019 2975
rect 4252 2941 4286 2975
rect 8484 2941 8518 2975
rect 11069 2941 11103 2975
rect 12449 2941 12483 2975
rect 13093 2941 13127 2975
rect 13829 2941 13863 2975
rect 14105 2941 14139 2975
rect 14565 2941 14599 2975
rect 15393 2941 15427 2975
rect 15669 2941 15703 2975
rect 16129 2941 16163 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 18797 2941 18831 2975
rect 19533 2941 19567 2975
rect 20545 2941 20579 2975
rect 1860 2873 1894 2907
rect 10425 2873 10459 2907
rect 11345 2873 11379 2907
rect 13369 2873 13403 2907
rect 17509 2873 17543 2907
rect 18337 2873 18371 2907
rect 19073 2873 19107 2907
rect 9597 2805 9631 2839
rect 10057 2805 10091 2839
rect 12633 2805 12667 2839
rect 14749 2805 14783 2839
rect 16313 2805 16347 2839
rect 20729 2805 20763 2839
rect 3525 2601 3559 2635
rect 4077 2601 4111 2635
rect 4445 2601 4479 2635
rect 4537 2601 4571 2635
rect 6561 2601 6595 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 2412 2533 2446 2567
rect 7205 2533 7239 2567
rect 10149 2533 10183 2567
rect 2145 2465 2179 2499
rect 5181 2465 5215 2499
rect 5448 2465 5482 2499
rect 6929 2465 6963 2499
rect 11713 2465 11747 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16129 2465 16163 2499
rect 16405 2465 16439 2499
rect 16865 2465 16899 2499
rect 17417 2465 17451 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19901 2465 19935 2499
rect 4629 2397 4663 2431
rect 10333 2397 10367 2431
rect 11989 2397 12023 2431
rect 20085 2397 20119 2431
rect 19073 2329 19107 2363
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 13921 2261 13955 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 17049 2261 17083 2295
rect 17601 2261 17635 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2774 20040 2780 20052
rect 2087 20012 2780 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19904 2467 19907
rect 7190 19904 7196 19916
rect 2455 19876 7196 19904
rect 2455 19873 2467 19876
rect 2409 19867 2467 19873
rect 1872 19836 1900 19867
rect 7190 19864 7196 19876
rect 7248 19864 7254 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15252 19876 15853 19904
rect 15252 19864 15258 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 15841 19867 15899 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19978 19904 19984 19916
rect 19939 19876 19984 19904
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20070 19864 20076 19916
rect 20128 19904 20134 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20128 19876 20545 19904
rect 20128 19864 20134 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 5166 19836 5172 19848
rect 1872 19808 5172 19836
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15344 19808 15945 19836
rect 15344 19796 15350 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16022 19796 16028 19848
rect 16080 19836 16086 19848
rect 16080 19808 16125 19836
rect 16080 19796 16086 19808
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 2958 19768 2964 19780
rect 2639 19740 2964 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 2958 19728 2964 19740
rect 3016 19728 3022 19780
rect 15473 19703 15531 19709
rect 15473 19669 15485 19703
rect 15519 19700 15531 19703
rect 17954 19700 17960 19712
rect 15519 19672 17960 19700
rect 15519 19669 15531 19672
rect 15473 19663 15531 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20680 19672 20729 19700
rect 20680 19660 20686 19672
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 2038 19496 2044 19508
rect 1999 19468 2044 19496
rect 2038 19456 2044 19468
rect 2096 19456 2102 19508
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 4120 19468 5365 19496
rect 4120 19456 4126 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5353 19459 5411 19465
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 16022 19496 16028 19508
rect 15887 19468 16028 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 19702 19496 19708 19508
rect 19659 19468 19708 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 20162 19496 20168 19508
rect 20123 19468 20168 19496
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 7742 19360 7748 19372
rect 7703 19332 7748 19360
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 8312 19332 8616 19360
rect 1854 19292 1860 19304
rect 1815 19264 1860 19292
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2409 19295 2467 19301
rect 2409 19261 2421 19295
rect 2455 19261 2467 19295
rect 3142 19292 3148 19304
rect 3103 19264 3148 19292
rect 2409 19255 2467 19261
rect 2424 19224 2452 19255
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 5074 19292 5080 19304
rect 3344 19264 5080 19292
rect 3344 19224 3372 19264
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 5169 19295 5227 19301
rect 5169 19261 5181 19295
rect 5215 19261 5227 19295
rect 5169 19255 5227 19261
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 7006 19292 7012 19304
rect 5767 19264 7012 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 2424 19196 3372 19224
rect 3412 19227 3470 19233
rect 3412 19193 3424 19227
rect 3458 19224 3470 19227
rect 3602 19224 3608 19236
rect 3458 19196 3608 19224
rect 3458 19193 3470 19196
rect 3412 19187 3470 19193
rect 3602 19184 3608 19196
rect 3660 19184 3666 19236
rect 5184 19224 5212 19255
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 8312 19292 8340 19332
rect 8478 19292 8484 19304
rect 7392 19264 8340 19292
rect 8439 19264 8484 19292
rect 5997 19227 6055 19233
rect 5997 19224 6009 19227
rect 5184 19196 6009 19224
rect 5997 19193 6009 19196
rect 6043 19193 6055 19227
rect 7392 19224 7420 19264
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 8588 19292 8616 19332
rect 10134 19292 10140 19304
rect 8588 19264 8892 19292
rect 10095 19264 10140 19292
rect 5997 19187 6055 19193
rect 7024 19196 7420 19224
rect 7469 19227 7527 19233
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2866 19156 2872 19168
rect 2639 19128 2872 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4525 19159 4583 19165
rect 4525 19156 4537 19159
rect 4212 19128 4537 19156
rect 4212 19116 4218 19128
rect 4525 19125 4537 19128
rect 4571 19125 4583 19159
rect 4525 19119 4583 19125
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 7024 19156 7052 19196
rect 7469 19193 7481 19227
rect 7515 19224 7527 19227
rect 7650 19224 7656 19236
rect 7515 19196 7656 19224
rect 7515 19193 7527 19196
rect 7469 19187 7527 19193
rect 7650 19184 7656 19196
rect 7708 19184 7714 19236
rect 7742 19184 7748 19236
rect 7800 19224 7806 19236
rect 8726 19227 8784 19233
rect 8726 19224 8738 19227
rect 7800 19196 8738 19224
rect 7800 19184 7806 19196
rect 8726 19193 8738 19196
rect 8772 19193 8784 19227
rect 8864 19224 8892 19264
rect 10134 19252 10140 19264
rect 10192 19252 10198 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 10836 19264 12449 19292
rect 10836 19252 10842 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 14458 19292 14464 19304
rect 14419 19264 14464 19292
rect 12437 19255 12495 19261
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 17126 19292 17132 19304
rect 14660 19264 17132 19292
rect 12710 19233 12716 19236
rect 10382 19227 10440 19233
rect 10382 19224 10394 19227
rect 8864 19196 10394 19224
rect 8726 19187 8784 19193
rect 10382 19193 10394 19196
rect 10428 19193 10440 19227
rect 12704 19224 12716 19233
rect 10382 19187 10440 19193
rect 11348 19196 11652 19224
rect 12671 19196 12716 19224
rect 5776 19128 7052 19156
rect 7101 19159 7159 19165
rect 5776 19116 5782 19128
rect 7101 19125 7113 19159
rect 7147 19156 7159 19159
rect 7374 19156 7380 19168
rect 7147 19128 7380 19156
rect 7147 19125 7159 19128
rect 7101 19119 7159 19125
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 7558 19156 7564 19168
rect 7519 19128 7564 19156
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 9858 19156 9864 19168
rect 9819 19128 9864 19156
rect 9858 19116 9864 19128
rect 9916 19156 9922 19168
rect 11348 19156 11376 19196
rect 11514 19156 11520 19168
rect 9916 19128 11376 19156
rect 11475 19128 11520 19156
rect 9916 19116 9922 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11624 19156 11652 19196
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 14660 19224 14688 19264
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 19150 19292 19156 19304
rect 18923 19264 19156 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19760 19264 19993 19292
rect 19760 19252 19766 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 19981 19255 20039 19261
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 12820 19196 14688 19224
rect 14728 19227 14786 19233
rect 12820 19156 12848 19196
rect 14728 19193 14740 19227
rect 14774 19224 14786 19227
rect 15562 19224 15568 19236
rect 14774 19196 15568 19224
rect 14774 19193 14786 19196
rect 14728 19187 14786 19193
rect 11624 19128 12848 19156
rect 13817 19159 13875 19165
rect 13817 19125 13829 19159
rect 13863 19156 13875 19159
rect 14752 19156 14780 19187
rect 15562 19184 15568 19196
rect 15620 19184 15626 19236
rect 19058 19156 19064 19168
rect 13863 19128 14780 19156
rect 19019 19128 19064 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 2501 18955 2559 18961
rect 2501 18921 2513 18955
rect 2547 18952 2559 18955
rect 2774 18952 2780 18964
rect 2547 18924 2780 18952
rect 2547 18921 2559 18924
rect 2501 18915 2559 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 3050 18952 3056 18964
rect 3011 18924 3056 18952
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 7742 18912 7748 18964
rect 7800 18952 7806 18964
rect 8021 18955 8079 18961
rect 8021 18952 8033 18955
rect 7800 18924 8033 18952
rect 7800 18912 7806 18924
rect 8021 18921 8033 18924
rect 8067 18921 8079 18955
rect 8021 18915 8079 18921
rect 2884 18856 7972 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 1765 18779 1823 18785
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 2498 18816 2504 18828
rect 2363 18788 2504 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 1780 18680 1808 18779
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 2884 18825 2912 18856
rect 4982 18825 4988 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 4976 18816 4988 18825
rect 4943 18788 4988 18816
rect 2869 18779 2927 18785
rect 4976 18779 4988 18788
rect 4982 18776 4988 18779
rect 5040 18776 5046 18828
rect 6908 18819 6966 18825
rect 6908 18785 6920 18819
rect 6954 18816 6966 18819
rect 7282 18816 7288 18828
rect 6954 18788 7288 18816
rect 6954 18785 6966 18788
rect 6908 18779 6966 18785
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 3142 18708 3148 18760
rect 3200 18748 3206 18760
rect 4706 18748 4712 18760
rect 3200 18720 4712 18748
rect 3200 18708 3206 18720
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 1780 18652 4752 18680
rect 4724 18612 4752 18652
rect 5626 18612 5632 18624
rect 4724 18584 5632 18612
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 6086 18612 6092 18624
rect 6047 18584 6092 18612
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6656 18612 6684 18711
rect 7944 18680 7972 18856
rect 8036 18748 8064 18915
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 10134 18952 10140 18964
rect 8260 18924 10140 18952
rect 8260 18912 8266 18924
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 13081 18955 13139 18961
rect 13081 18921 13093 18955
rect 13127 18952 13139 18955
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 13127 18924 14473 18952
rect 13127 18921 13139 18924
rect 13081 18915 13139 18921
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 14461 18915 14519 18921
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 19300 18924 19533 18952
rect 19300 18912 19306 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 8757 18887 8815 18893
rect 8757 18853 8769 18887
rect 8803 18884 8815 18887
rect 10318 18884 10324 18896
rect 8803 18856 10324 18884
rect 8803 18853 8815 18856
rect 8757 18847 8815 18853
rect 10318 18844 10324 18856
rect 10376 18844 10382 18896
rect 13538 18844 13544 18896
rect 13596 18884 13602 18896
rect 16022 18893 16028 18896
rect 14553 18887 14611 18893
rect 14553 18884 14565 18887
rect 13596 18856 14565 18884
rect 13596 18844 13602 18856
rect 14553 18853 14565 18856
rect 14599 18853 14611 18887
rect 16016 18884 16028 18893
rect 15983 18856 16028 18884
rect 14553 18847 14611 18853
rect 16016 18847 16028 18856
rect 16022 18844 16028 18847
rect 16080 18844 16086 18896
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20165 18887 20223 18893
rect 20165 18884 20177 18887
rect 20036 18856 20177 18884
rect 20036 18844 20042 18856
rect 20165 18853 20177 18856
rect 20211 18853 20223 18887
rect 20165 18847 20223 18853
rect 8849 18819 8907 18825
rect 8849 18785 8861 18819
rect 8895 18816 8907 18819
rect 9674 18816 9680 18828
rect 8895 18788 9680 18816
rect 8895 18785 8907 18788
rect 8849 18779 8907 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11232 18819 11290 18825
rect 11232 18785 11244 18819
rect 11278 18816 11290 18819
rect 11514 18816 11520 18828
rect 11278 18788 11520 18816
rect 11278 18785 11290 18788
rect 11232 18779 11290 18785
rect 11514 18776 11520 18788
rect 11572 18816 11578 18828
rect 12621 18819 12679 18825
rect 11572 18788 12020 18816
rect 11572 18776 11578 18788
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8036 18720 8953 18748
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 10965 18751 11023 18757
rect 10965 18748 10977 18751
rect 10836 18720 10977 18748
rect 10836 18708 10842 18720
rect 10965 18717 10977 18720
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 9950 18680 9956 18692
rect 7944 18652 9956 18680
rect 9950 18640 9956 18652
rect 10008 18640 10014 18692
rect 8202 18612 8208 18624
rect 6656 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8386 18612 8392 18624
rect 8347 18584 8392 18612
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 11992 18612 12020 18788
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 13449 18819 13507 18825
rect 13449 18816 13461 18819
rect 12667 18788 13461 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 13449 18785 13461 18788
rect 13495 18785 13507 18819
rect 13630 18816 13636 18828
rect 13449 18779 13507 18785
rect 13556 18788 13636 18816
rect 13556 18757 13584 18788
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 14458 18776 14464 18828
rect 14516 18816 14522 18828
rect 15749 18819 15807 18825
rect 15749 18816 15761 18819
rect 14516 18788 15761 18816
rect 14516 18776 14522 18788
rect 15749 18785 15761 18788
rect 15795 18816 15807 18819
rect 16574 18816 16580 18828
rect 15795 18788 16580 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18816 19395 18819
rect 19518 18816 19524 18828
rect 19383 18788 19524 18816
rect 19383 18785 19395 18788
rect 19337 18779 19395 18785
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 19610 18776 19616 18828
rect 19668 18816 19674 18828
rect 19889 18819 19947 18825
rect 19889 18816 19901 18819
rect 19668 18788 19901 18816
rect 19668 18776 19674 18788
rect 19889 18785 19901 18788
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13722 18748 13728 18760
rect 13683 18720 13728 18748
rect 13541 18711 13599 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 15562 18748 15568 18760
rect 14783 18720 15568 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 12345 18683 12403 18689
rect 12345 18649 12357 18683
rect 12391 18680 12403 18683
rect 12710 18680 12716 18692
rect 12391 18652 12716 18680
rect 12391 18649 12403 18652
rect 12345 18643 12403 18649
rect 12710 18640 12716 18652
rect 12768 18680 12774 18692
rect 13740 18680 13768 18708
rect 12768 18652 13768 18680
rect 14093 18683 14151 18689
rect 12768 18640 12774 18652
rect 14093 18649 14105 18683
rect 14139 18680 14151 18683
rect 15194 18680 15200 18692
rect 14139 18652 15200 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 14182 18612 14188 18624
rect 11992 18584 14188 18612
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 17126 18612 17132 18624
rect 17087 18584 17132 18612
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 7006 18408 7012 18420
rect 1780 18380 6868 18408
rect 6967 18380 7012 18408
rect 1780 18213 1808 18380
rect 1946 18340 1952 18352
rect 1907 18312 1952 18340
rect 1946 18300 1952 18312
rect 2004 18300 2010 18352
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 3283 18244 3740 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3605 18207 3663 18213
rect 3605 18204 3617 18207
rect 3200 18176 3617 18204
rect 3200 18164 3206 18176
rect 3605 18173 3617 18176
rect 3651 18173 3663 18207
rect 3712 18204 3740 18244
rect 3872 18207 3930 18213
rect 3872 18204 3884 18207
rect 3712 18176 3884 18204
rect 3605 18167 3663 18173
rect 3872 18173 3884 18176
rect 3918 18204 3930 18207
rect 4154 18204 4160 18216
rect 3918 18176 4160 18204
rect 3918 18173 3930 18176
rect 3872 18167 3930 18173
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 1854 18096 1860 18148
rect 1912 18136 1918 18148
rect 5994 18136 6000 18148
rect 1912 18108 6000 18136
rect 1912 18096 1918 18108
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 2590 18068 2596 18080
rect 2551 18040 2596 18068
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3050 18028 3056 18080
rect 3108 18068 3114 18080
rect 4982 18068 4988 18080
rect 3108 18040 3153 18068
rect 4943 18040 4988 18068
rect 3108 18028 3114 18040
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 6840 18068 6868 18380
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 10318 18408 10324 18420
rect 10279 18380 10324 18408
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 20070 18408 20076 18420
rect 13688 18380 20076 18408
rect 13688 18368 13694 18380
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 8386 18340 8392 18352
rect 7484 18312 8392 18340
rect 7484 18281 7512 18312
rect 8386 18300 8392 18312
rect 8444 18300 8450 18352
rect 13265 18343 13323 18349
rect 13265 18309 13277 18343
rect 13311 18340 13323 18343
rect 15102 18340 15108 18352
rect 13311 18312 15108 18340
rect 13311 18309 13323 18312
rect 13265 18303 13323 18309
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 20162 18340 20168 18352
rect 20123 18312 20168 18340
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 7374 18204 7380 18216
rect 7335 18176 7380 18204
rect 7374 18164 7380 18176
rect 7432 18164 7438 18216
rect 7576 18204 7604 18235
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7708 18244 8033 18272
rect 7708 18232 7714 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8021 18235 8079 18241
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8260 18244 8677 18272
rect 8260 18232 8266 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 10042 18232 10048 18284
rect 10100 18272 10106 18284
rect 10873 18275 10931 18281
rect 10873 18272 10885 18275
rect 10100 18244 10885 18272
rect 10100 18232 10106 18244
rect 10873 18241 10885 18244
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13780 18244 13921 18272
rect 13780 18232 13786 18244
rect 13909 18241 13921 18244
rect 13955 18272 13967 18275
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 13955 18244 15669 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 15657 18235 15715 18241
rect 16500 18244 16681 18272
rect 16500 18216 16528 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 9858 18204 9864 18216
rect 7576 18176 9864 18204
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 16482 18204 16488 18216
rect 14240 18176 16488 18204
rect 14240 18164 14246 18176
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 16577 18207 16635 18213
rect 16577 18173 16589 18207
rect 16623 18204 16635 18207
rect 16850 18204 16856 18216
rect 16623 18176 16856 18204
rect 16623 18173 16635 18176
rect 16577 18167 16635 18173
rect 16850 18164 16856 18176
rect 16908 18204 16914 18216
rect 17862 18204 17868 18216
rect 16908 18176 17868 18204
rect 16908 18164 16914 18176
rect 17862 18164 17868 18176
rect 17920 18164 17926 18216
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 18012 18176 18245 18204
rect 18012 18164 18018 18176
rect 18233 18173 18245 18176
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 19153 18207 19211 18213
rect 19153 18204 19165 18207
rect 18555 18176 19165 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 19153 18173 19165 18176
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 19518 18164 19524 18216
rect 19576 18204 19582 18216
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 19576 18176 19993 18204
rect 19576 18164 19582 18176
rect 19981 18173 19993 18176
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20128 18176 20545 18204
rect 20128 18164 20134 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 8754 18096 8760 18148
rect 8812 18136 8818 18148
rect 8910 18139 8968 18145
rect 8910 18136 8922 18139
rect 8812 18108 8922 18136
rect 8812 18096 8818 18108
rect 8910 18105 8922 18108
rect 8956 18105 8968 18139
rect 8910 18099 8968 18105
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11054 18136 11060 18148
rect 10735 18108 11060 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11054 18096 11060 18108
rect 11112 18096 11118 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 12084 18108 13645 18136
rect 9766 18068 9772 18080
rect 6840 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 10468 18040 10793 18068
rect 10468 18028 10474 18040
rect 10781 18037 10793 18040
rect 10827 18068 10839 18071
rect 12084 18068 12112 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 15746 18136 15752 18148
rect 13633 18099 13691 18105
rect 15120 18108 15752 18136
rect 13722 18068 13728 18080
rect 10827 18040 12112 18068
rect 13683 18040 13728 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 15120 18077 15148 18108
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18037 15163 18071
rect 15470 18068 15476 18080
rect 15431 18040 15476 18068
rect 15105 18031 15163 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 15565 18071 15623 18077
rect 15565 18037 15577 18071
rect 15611 18068 15623 18071
rect 16117 18071 16175 18077
rect 16117 18068 16129 18071
rect 15611 18040 16129 18068
rect 15611 18037 15623 18040
rect 15565 18031 15623 18037
rect 16117 18037 16129 18040
rect 16163 18037 16175 18071
rect 16117 18031 16175 18037
rect 16485 18071 16543 18077
rect 16485 18037 16497 18071
rect 16531 18068 16543 18071
rect 16758 18068 16764 18080
rect 16531 18040 16764 18068
rect 16531 18037 16543 18040
rect 16485 18031 16543 18037
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19337 18071 19395 18077
rect 19337 18068 19349 18071
rect 19024 18040 19349 18068
rect 19024 18028 19030 18040
rect 19337 18037 19349 18040
rect 19383 18037 19395 18071
rect 19337 18031 19395 18037
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20680 18040 20729 18068
rect 20680 18028 20686 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2590 17864 2596 17876
rect 2363 17836 2596 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 2958 17864 2964 17876
rect 2919 17836 2964 17864
rect 2958 17824 2964 17836
rect 3016 17824 3022 17876
rect 4982 17864 4988 17876
rect 4080 17836 4988 17864
rect 4080 17796 4108 17836
rect 4982 17824 4988 17836
rect 5040 17824 5046 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12529 17867 12587 17873
rect 12529 17864 12541 17867
rect 11112 17836 12541 17864
rect 11112 17824 11118 17836
rect 12529 17833 12541 17836
rect 12575 17833 12587 17867
rect 12529 17827 12587 17833
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13722 17864 13728 17876
rect 13679 17836 13728 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15746 17864 15752 17876
rect 15707 17836 15752 17864
rect 15746 17824 15752 17836
rect 15804 17824 15810 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 19426 17864 19432 17876
rect 19116 17836 19432 17864
rect 19116 17824 19122 17836
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 2608 17768 4108 17796
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17697 1455 17731
rect 1397 17691 1455 17697
rect 1412 17592 1440 17691
rect 2608 17669 2636 17768
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4212 17768 4936 17796
rect 4212 17756 4218 17768
rect 3326 17728 3332 17740
rect 3287 17700 3332 17728
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 4632 17700 4721 17728
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17629 2651 17663
rect 3418 17660 3424 17672
rect 3379 17632 3424 17660
rect 2593 17623 2651 17629
rect 2424 17592 2452 17623
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 3602 17660 3608 17672
rect 3563 17632 3608 17660
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 4341 17595 4399 17601
rect 4341 17592 4353 17595
rect 1412 17564 2268 17592
rect 2424 17564 4353 17592
rect 1949 17527 2007 17533
rect 1949 17493 1961 17527
rect 1995 17524 2007 17527
rect 2038 17524 2044 17536
rect 1995 17496 2044 17524
rect 1995 17493 2007 17496
rect 1949 17487 2007 17493
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 2240 17524 2268 17564
rect 4341 17561 4353 17564
rect 4387 17561 4399 17595
rect 4632 17592 4660 17700
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 4908 17669 4936 17768
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 5684 17768 6929 17796
rect 5684 17756 5690 17768
rect 6917 17765 6929 17768
rect 6963 17765 6975 17799
rect 14001 17799 14059 17805
rect 14001 17796 14013 17799
rect 6917 17759 6975 17765
rect 10060 17768 14013 17796
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 8018 17728 8024 17740
rect 6687 17700 8024 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10060 17737 10088 17768
rect 14001 17765 14013 17768
rect 14047 17765 14059 17799
rect 14001 17759 14059 17765
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 15657 17799 15715 17805
rect 15657 17796 15669 17799
rect 15160 17768 15669 17796
rect 15160 17756 15166 17768
rect 15657 17765 15669 17768
rect 15703 17765 15715 17799
rect 15657 17759 15715 17765
rect 16844 17799 16902 17805
rect 16844 17765 16856 17799
rect 16890 17796 16902 17799
rect 16942 17796 16948 17808
rect 16890 17768 16948 17796
rect 16890 17765 16902 17768
rect 16844 17759 16902 17765
rect 16942 17756 16948 17768
rect 17000 17756 17006 17808
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20530 17796 20536 17808
rect 20027 17768 20536 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9916 17700 10057 17728
rect 9916 17688 9922 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10318 17728 10324 17740
rect 10183 17700 10324 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 10152 17660 10180 17691
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 13078 17728 13084 17740
rect 12483 17700 13084 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 17310 17688 17316 17740
rect 17368 17728 17374 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 17368 17700 19717 17728
rect 17368 17688 17374 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 9824 17632 10180 17660
rect 10229 17663 10287 17669
rect 9824 17620 9830 17632
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 12710 17660 12716 17672
rect 12671 17632 12716 17660
rect 10229 17623 10287 17629
rect 6730 17592 6736 17604
rect 4632 17564 6736 17592
rect 4341 17555 4399 17561
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 10042 17592 10048 17604
rect 7340 17564 10048 17592
rect 7340 17552 7346 17564
rect 10042 17552 10048 17564
rect 10100 17592 10106 17604
rect 10244 17592 10272 17623
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14240 17632 14285 17660
rect 14240 17620 14246 17632
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15620 17632 15853 17660
rect 15620 17620 15626 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 16574 17660 16580 17672
rect 16487 17632 16580 17660
rect 15841 17623 15899 17629
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 10100 17564 10272 17592
rect 12069 17595 12127 17601
rect 10100 17552 10106 17564
rect 12069 17561 12081 17595
rect 12115 17592 12127 17595
rect 13538 17592 13544 17604
rect 12115 17564 13544 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 10134 17524 10140 17536
rect 2240 17496 10140 17524
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 16592 17524 16620 17620
rect 17770 17524 17776 17536
rect 16592 17496 17776 17524
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 17954 17524 17960 17536
rect 17915 17496 17960 17524
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 4798 17320 4804 17332
rect 4759 17292 4804 17320
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 7558 17320 7564 17332
rect 6871 17292 7564 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8018 17320 8024 17332
rect 7979 17292 8024 17320
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 15528 17292 16037 17320
rect 15528 17280 15534 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 16025 17283 16083 17289
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1504 17156 2237 17184
rect 1504 17125 1532 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3660 17156 3709 17184
rect 3660 17144 3666 17156
rect 3697 17153 3709 17156
rect 3743 17184 3755 17187
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 3743 17156 5457 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 5445 17153 5457 17156
rect 5491 17184 5503 17187
rect 6454 17184 6460 17196
rect 5491 17156 6460 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7340 17156 7389 17184
rect 7340 17144 7346 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17184 8723 17187
rect 8754 17184 8760 17196
rect 8711 17156 8760 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 8754 17144 8760 17156
rect 8812 17144 8818 17196
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 12124 17156 13921 17184
rect 12124 17144 12130 17156
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16577 17187 16635 17193
rect 16577 17184 16589 17187
rect 16540 17156 16589 17184
rect 16540 17144 16546 17156
rect 16577 17153 16589 17156
rect 16623 17153 16635 17187
rect 16577 17147 16635 17153
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 2038 17116 2044 17128
rect 1999 17088 2044 17116
rect 1489 17079 1547 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 3421 17119 3479 17125
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 3510 17116 3516 17128
rect 3467 17088 3516 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10778 17116 10784 17128
rect 10735 17088 10784 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10778 17076 10784 17088
rect 10836 17116 10842 17128
rect 10836 17088 11652 17116
rect 10836 17076 10842 17088
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 7064 17020 7297 17048
rect 7064 17008 7070 17020
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 8386 17048 8392 17060
rect 8347 17020 8392 17048
rect 7285 17011 7343 17017
rect 8386 17008 8392 17020
rect 8444 17008 8450 17060
rect 10962 17057 10968 17060
rect 10956 17011 10968 17057
rect 11020 17048 11026 17060
rect 11624 17048 11652 17088
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 11756 17088 13737 17116
rect 11756 17076 11762 17088
rect 13725 17085 13737 17088
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 18141 17119 18199 17125
rect 18141 17116 18153 17119
rect 17828 17088 18153 17116
rect 17828 17076 17834 17088
rect 18141 17085 18153 17088
rect 18187 17085 18199 17119
rect 18141 17079 18199 17085
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 20162 17116 20168 17128
rect 20027 17088 20168 17116
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 12618 17048 12624 17060
rect 11020 17020 11056 17048
rect 11624 17020 12624 17048
rect 10962 17008 10968 17011
rect 11020 17008 11026 17020
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 13906 17048 13912 17060
rect 13372 17020 13912 17048
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 3513 16983 3571 16989
rect 3513 16949 3525 16983
rect 3559 16980 3571 16983
rect 4246 16980 4252 16992
rect 3559 16952 4252 16980
rect 3559 16949 3571 16952
rect 3513 16943 3571 16949
rect 4246 16940 4252 16952
rect 4304 16980 4310 16992
rect 4706 16980 4712 16992
rect 4304 16952 4712 16980
rect 4304 16940 4310 16952
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 5169 16983 5227 16989
rect 5169 16980 5181 16983
rect 4948 16952 5181 16980
rect 4948 16940 4954 16952
rect 5169 16949 5181 16952
rect 5215 16949 5227 16983
rect 5169 16943 5227 16949
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 5316 16952 5361 16980
rect 5316 16940 5322 16952
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 7193 16983 7251 16989
rect 7193 16980 7205 16983
rect 6696 16952 7205 16980
rect 6696 16940 6702 16952
rect 7193 16949 7205 16952
rect 7239 16949 7251 16983
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 7193 16943 7251 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 12066 16980 12072 16992
rect 12027 16952 12072 16980
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 13372 16989 13400 17020
rect 13906 17008 13912 17020
rect 13964 17008 13970 17060
rect 16393 17051 16451 17057
rect 16393 17017 16405 17051
rect 16439 17048 16451 17051
rect 17678 17048 17684 17060
rect 16439 17020 17684 17048
rect 16439 17017 16451 17020
rect 16393 17011 16451 17017
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 18408 17051 18466 17057
rect 18408 17017 18420 17051
rect 18454 17048 18466 17051
rect 19426 17048 19432 17060
rect 18454 17020 19432 17048
rect 18454 17017 18466 17020
rect 18408 17011 18466 17017
rect 19426 17008 19432 17020
rect 19484 17008 19490 17060
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20548 17048 20576 17079
rect 19760 17020 20576 17048
rect 19760 17008 19766 17020
rect 13357 16983 13415 16989
rect 13357 16949 13369 16983
rect 13403 16949 13415 16983
rect 13357 16943 13415 16949
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16980 13875 16983
rect 15286 16980 15292 16992
rect 13863 16952 15292 16980
rect 13863 16949 13875 16952
rect 13817 16943 13875 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 16482 16980 16488 16992
rect 16443 16952 16488 16980
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 19521 16983 19579 16989
rect 19521 16980 19533 16983
rect 17000 16952 19533 16980
rect 17000 16940 17006 16952
rect 19521 16949 19533 16952
rect 19567 16949 19579 16983
rect 19521 16943 19579 16949
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 20717 16983 20775 16989
rect 20717 16980 20729 16983
rect 20680 16952 20729 16980
rect 20680 16940 20686 16952
rect 20717 16949 20729 16952
rect 20763 16949 20775 16983
rect 20717 16943 20775 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2774 16776 2780 16788
rect 2547 16748 2780 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2924 16748 3065 16776
rect 2924 16736 2930 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 3053 16739 3111 16745
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 3384 16748 3433 16776
rect 3384 16736 3390 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 3421 16739 3479 16745
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 9033 16779 9091 16785
rect 9033 16776 9045 16779
rect 8812 16748 9045 16776
rect 8812 16736 8818 16748
rect 9033 16745 9045 16748
rect 9079 16745 9091 16779
rect 9033 16739 9091 16745
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 15286 16776 15292 16788
rect 12124 16748 12756 16776
rect 15247 16748 15292 16776
rect 12124 16736 12130 16748
rect 8202 16708 8208 16720
rect 7668 16680 8208 16708
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2314 16640 2320 16652
rect 2275 16612 2320 16640
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2866 16640 2872 16652
rect 2827 16612 2872 16640
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 4798 16600 4804 16652
rect 4856 16640 4862 16652
rect 5350 16649 5356 16652
rect 5077 16643 5135 16649
rect 5077 16640 5089 16643
rect 4856 16612 5089 16640
rect 4856 16600 4862 16612
rect 5077 16609 5089 16612
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5344 16603 5356 16649
rect 5408 16640 5414 16652
rect 7668 16649 7696 16680
rect 8202 16668 8208 16680
rect 8260 16668 8266 16720
rect 11885 16711 11943 16717
rect 11885 16677 11897 16711
rect 11931 16708 11943 16711
rect 12434 16708 12440 16720
rect 11931 16680 12440 16708
rect 11931 16677 11943 16680
rect 11885 16671 11943 16677
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 12728 16708 12756 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15795 16748 16313 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 19886 16776 19892 16788
rect 19847 16748 19892 16776
rect 16301 16739 16359 16745
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 12958 16711 13016 16717
rect 12958 16708 12970 16711
rect 12728 16680 12970 16708
rect 12958 16677 12970 16680
rect 13004 16677 13016 16711
rect 12958 16671 13016 16677
rect 16761 16711 16819 16717
rect 16761 16677 16773 16711
rect 16807 16708 16819 16711
rect 16850 16708 16856 16720
rect 16807 16680 16856 16708
rect 16807 16677 16819 16680
rect 16761 16671 16819 16677
rect 16850 16668 16856 16680
rect 16908 16668 16914 16720
rect 19794 16668 19800 16720
rect 19852 16708 19858 16720
rect 19852 16680 20300 16708
rect 19852 16668 19858 16680
rect 7653 16643 7711 16649
rect 5408 16612 5444 16640
rect 5350 16600 5356 16603
rect 5408 16600 5414 16612
rect 7653 16609 7665 16643
rect 7699 16609 7711 16643
rect 7653 16603 7711 16609
rect 7920 16643 7978 16649
rect 7920 16609 7932 16643
rect 7966 16640 7978 16643
rect 9582 16640 9588 16652
rect 7966 16612 9588 16640
rect 7966 16609 7978 16612
rect 7920 16603 7978 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 14148 16612 15669 16640
rect 14148 16600 14154 16612
rect 15657 16609 15669 16612
rect 15703 16640 15715 16643
rect 16022 16640 16028 16652
rect 15703 16612 16028 16640
rect 15703 16609 15715 16612
rect 15657 16603 15715 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16482 16600 16488 16652
rect 16540 16640 16546 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16540 16612 16681 16640
rect 16540 16600 16546 16612
rect 16669 16609 16681 16612
rect 16715 16640 16727 16643
rect 17586 16640 17592 16652
rect 16715 16612 17592 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 19978 16640 19984 16652
rect 19751 16612 19984 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20272 16649 20300 16680
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11974 16572 11980 16584
rect 11204 16544 11980 16572
rect 11204 16532 11210 16544
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 1946 16504 1952 16516
rect 1907 16476 1952 16504
rect 1946 16464 1952 16476
rect 2004 16464 2010 16516
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 12084 16504 12112 16535
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 12676 16544 12725 16572
rect 12676 16532 12682 16544
rect 12713 16541 12725 16544
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16541 15991 16575
rect 16942 16572 16948 16584
rect 16903 16544 16948 16572
rect 15933 16535 15991 16541
rect 15948 16504 15976 16535
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17954 16504 17960 16516
rect 11020 16476 12112 16504
rect 11020 16464 11026 16476
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 11517 16439 11575 16445
rect 11517 16405 11529 16439
rect 11563 16436 11575 16439
rect 11790 16436 11796 16448
rect 11563 16408 11796 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 12084 16436 12112 16476
rect 13648 16476 17960 16504
rect 13648 16436 13676 16476
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 14090 16436 14096 16448
rect 12084 16408 13676 16436
rect 14051 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 20438 16436 20444 16448
rect 20399 16408 20444 16436
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 4985 16235 5043 16241
rect 4985 16201 4997 16235
rect 5031 16232 5043 16235
rect 5258 16232 5264 16244
rect 5031 16204 5264 16232
rect 5031 16201 5043 16204
rect 4985 16195 5043 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6788 16204 6837 16232
rect 6788 16192 6794 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 8496 16204 9536 16232
rect 4890 16124 4896 16176
rect 4948 16164 4954 16176
rect 8496 16164 8524 16204
rect 4948 16136 8524 16164
rect 4948 16124 4954 16136
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 5350 16056 5356 16108
rect 5408 16096 5414 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5408 16068 5549 16096
rect 5408 16056 5414 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 6512 16068 7389 16096
rect 6512 16056 6518 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 9508 16096 9536 16204
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9640 16204 9873 16232
rect 9640 16192 9646 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 11698 16232 11704 16244
rect 10367 16204 11704 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 15378 16232 15384 16244
rect 13924 16204 15384 16232
rect 9950 16124 9956 16176
rect 10008 16164 10014 16176
rect 10008 16136 13860 16164
rect 10008 16124 10014 16136
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 9508 16068 10793 16096
rect 7377 16059 7435 16065
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10781 16059 10839 16065
rect 10962 16056 10968 16068
rect 11020 16096 11026 16108
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11020 16068 11897 16096
rect 11020 16056 11026 16068
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12492 16068 12537 16096
rect 12492 16056 12498 16068
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 6914 16028 6920 16040
rect 2087 16000 6920 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8260 16000 8493 16028
rect 8260 15988 8266 16000
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 8481 15991 8539 15997
rect 8588 16000 11805 16028
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 5442 15960 5448 15972
rect 1820 15932 5448 15960
rect 1820 15920 1826 15932
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 8588 15960 8616 16000
rect 10980 15972 11008 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 13832 16028 13860 16136
rect 13924 16105 13952 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 19426 16232 19432 16244
rect 19387 16204 19432 16232
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16065 13967 16099
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 13909 16059 13967 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 13832 16000 15884 16028
rect 11793 15991 11851 15997
rect 7239 15932 8616 15960
rect 8748 15963 8806 15969
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 8748 15929 8760 15963
rect 8794 15960 8806 15963
rect 10226 15960 10232 15972
rect 8794 15932 10232 15960
rect 8794 15929 8806 15932
rect 8748 15923 8806 15929
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 10962 15920 10968 15972
rect 11020 15920 11026 15972
rect 11701 15963 11759 15969
rect 11701 15929 11713 15963
rect 11747 15960 11759 15963
rect 11974 15960 11980 15972
rect 11747 15932 11980 15960
rect 11747 15929 11759 15932
rect 11701 15923 11759 15929
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 13998 15960 14004 15972
rect 12084 15932 14004 15960
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5224 15864 5365 15892
rect 5224 15852 5230 15864
rect 5353 15861 5365 15864
rect 5399 15892 5411 15895
rect 6822 15892 6828 15904
rect 5399 15864 6828 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7374 15892 7380 15904
rect 7331 15864 7380 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7374 15852 7380 15864
rect 7432 15892 7438 15904
rect 10689 15895 10747 15901
rect 10689 15892 10701 15895
rect 7432 15864 10701 15892
rect 7432 15852 7438 15864
rect 10689 15861 10701 15864
rect 10735 15861 10747 15895
rect 11330 15892 11336 15904
rect 11291 15864 11336 15892
rect 10689 15855 10747 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 12084 15892 12112 15932
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 14090 15920 14096 15972
rect 14148 15969 14154 15972
rect 14148 15963 14212 15969
rect 14148 15929 14166 15963
rect 14200 15929 14212 15963
rect 14148 15923 14212 15929
rect 14148 15920 14154 15923
rect 15286 15892 15292 15904
rect 11480 15864 12112 15892
rect 15247 15864 15292 15892
rect 11480 15852 11486 15864
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15856 15892 15884 16000
rect 15930 15988 15936 16040
rect 15988 16028 15994 16040
rect 17770 16028 17776 16040
rect 15988 16000 17776 16028
rect 15988 15988 15994 16000
rect 17770 15988 17776 16000
rect 17828 16028 17834 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17828 16000 18061 16028
rect 17828 15988 17834 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 15997 19855 16031
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 19797 15991 19855 15997
rect 17218 15920 17224 15972
rect 17276 15960 17282 15972
rect 18294 15963 18352 15969
rect 18294 15960 18306 15963
rect 17276 15932 18306 15960
rect 17276 15920 17282 15932
rect 18294 15929 18306 15932
rect 18340 15929 18352 15963
rect 19812 15960 19840 15991
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 19978 15960 19984 15972
rect 19812 15932 19984 15960
rect 18294 15923 18352 15929
rect 19978 15920 19984 15932
rect 20036 15920 20042 15972
rect 20254 15920 20260 15972
rect 20312 15960 20318 15972
rect 20809 15963 20867 15969
rect 20809 15960 20821 15963
rect 20312 15932 20821 15960
rect 20312 15920 20318 15932
rect 20809 15929 20821 15932
rect 20855 15929 20867 15963
rect 20809 15923 20867 15929
rect 19058 15892 19064 15904
rect 15856 15864 19064 15892
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 5258 15688 5264 15700
rect 2516 15660 5264 15688
rect 2516 15620 2544 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 5408 15660 5457 15688
rect 5408 15648 5414 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 5445 15651 5503 15657
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8536 15660 8585 15688
rect 8536 15648 8542 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9079 15660 9689 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 10134 15688 10140 15700
rect 10095 15660 10140 15688
rect 9677 15651 9735 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 11422 15688 11428 15700
rect 10244 15660 11428 15688
rect 1780 15592 2544 15620
rect 2584 15623 2642 15629
rect 1780 15561 1808 15592
rect 2584 15589 2596 15623
rect 2630 15620 2642 15623
rect 2682 15620 2688 15632
rect 2630 15592 2688 15620
rect 2630 15589 2642 15592
rect 2584 15583 2642 15589
rect 2682 15580 2688 15592
rect 2740 15580 2746 15632
rect 3881 15623 3939 15629
rect 3881 15620 3893 15623
rect 3620 15592 3893 15620
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 3620 15552 3648 15592
rect 3881 15589 3893 15592
rect 3927 15589 3939 15623
rect 3881 15583 3939 15589
rect 6080 15623 6138 15629
rect 6080 15589 6092 15623
rect 6126 15620 6138 15623
rect 6730 15620 6736 15632
rect 6126 15592 6736 15620
rect 6126 15589 6138 15592
rect 6080 15583 6138 15589
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 6880 15592 9076 15620
rect 6880 15580 6886 15592
rect 4321 15555 4379 15561
rect 4321 15552 4333 15555
rect 2363 15524 3648 15552
rect 3712 15524 4333 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 3712 15357 3740 15524
rect 4321 15521 4333 15524
rect 4367 15521 4379 15555
rect 4321 15515 4379 15521
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 4856 15524 5825 15552
rect 4856 15512 4862 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7156 15524 8033 15552
rect 7156 15512 7162 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8938 15552 8944 15564
rect 8899 15524 8944 15552
rect 8021 15515 8079 15521
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9048 15552 9076 15592
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 10008 15592 10057 15620
rect 10008 15580 10014 15592
rect 10045 15589 10057 15592
rect 10091 15589 10103 15623
rect 10045 15583 10103 15589
rect 10244 15552 10272 15660
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 11790 15688 11796 15700
rect 11751 15660 11796 15688
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15657 13507 15691
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 13449 15651 13507 15657
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 11885 15623 11943 15629
rect 11885 15620 11897 15623
rect 11388 15592 11897 15620
rect 11388 15580 11394 15592
rect 11885 15589 11897 15592
rect 11931 15589 11943 15623
rect 13464 15620 13492 15651
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 16666 15688 16672 15700
rect 14056 15660 16672 15688
rect 14056 15648 14062 15660
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 17218 15688 17224 15700
rect 17179 15660 17224 15688
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 20530 15688 20536 15700
rect 17328 15660 20536 15688
rect 17328 15620 17356 15660
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 13464 15592 17356 15620
rect 11885 15583 11943 15589
rect 18506 15580 18512 15632
rect 18564 15620 18570 15632
rect 19613 15623 19671 15629
rect 19613 15620 19625 15623
rect 18564 15592 19625 15620
rect 18564 15580 18570 15592
rect 19613 15589 19625 15592
rect 19659 15589 19671 15623
rect 19613 15583 19671 15589
rect 19702 15580 19708 15632
rect 19760 15580 19766 15632
rect 13817 15555 13875 15561
rect 13817 15552 13829 15555
rect 9048 15524 10272 15552
rect 11440 15524 13829 15552
rect 3881 15487 3939 15493
rect 3881 15453 3893 15487
rect 3927 15484 3939 15487
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 3927 15456 4077 15484
rect 3927 15453 3939 15456
rect 3881 15447 3939 15453
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9582 15484 9588 15496
rect 9263 15456 9588 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 3697 15351 3755 15357
rect 3697 15348 3709 15351
rect 3292 15320 3709 15348
rect 3292 15308 3298 15320
rect 3697 15317 3709 15320
rect 3743 15317 3755 15351
rect 4080 15348 4108 15447
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 10226 15484 10232 15496
rect 10187 15456 10232 15484
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 11440 15425 11468 15524
rect 13817 15521 13829 15524
rect 13863 15521 13875 15555
rect 13817 15515 13875 15521
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 15436 15524 15853 15552
rect 15436 15512 15442 15524
rect 15841 15521 15853 15524
rect 15887 15552 15899 15555
rect 15930 15552 15936 15564
rect 15887 15524 15936 15552
rect 15887 15521 15899 15524
rect 15841 15515 15899 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16108 15555 16166 15561
rect 16108 15521 16120 15555
rect 16154 15552 16166 15555
rect 16390 15552 16396 15564
rect 16154 15524 16396 15552
rect 16154 15521 16166 15524
rect 16108 15515 16166 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 18598 15552 18604 15564
rect 18559 15524 18604 15552
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 19061 15555 19119 15561
rect 18748 15524 18793 15552
rect 18748 15512 18754 15524
rect 19061 15521 19073 15555
rect 19107 15552 19119 15555
rect 19720 15552 19748 15580
rect 20254 15552 20260 15564
rect 19107 15524 19748 15552
rect 20215 15524 20260 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 12066 15484 12072 15496
rect 12027 15456 12072 15484
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 14090 15484 14096 15496
rect 14051 15456 14096 15484
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 18782 15484 18788 15496
rect 18743 15456 18788 15484
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 18932 15456 19717 15484
rect 18932 15444 18938 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 11425 15419 11483 15425
rect 11425 15385 11437 15419
rect 11471 15385 11483 15419
rect 11425 15379 11483 15385
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 19061 15419 19119 15425
rect 19061 15416 19073 15419
rect 12032 15388 15884 15416
rect 12032 15376 12038 15388
rect 4246 15348 4252 15360
rect 4080 15320 4252 15348
rect 3697 15311 3755 15317
rect 4246 15308 4252 15320
rect 4304 15348 4310 15360
rect 4798 15348 4804 15360
rect 4304 15320 4804 15348
rect 4304 15308 4310 15320
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 7193 15351 7251 15357
rect 7193 15317 7205 15351
rect 7239 15348 7251 15351
rect 7282 15348 7288 15360
rect 7239 15320 7288 15348
rect 7239 15317 7251 15320
rect 7193 15311 7251 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 8202 15348 8208 15360
rect 7883 15320 8208 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8202 15308 8208 15320
rect 8260 15348 8266 15360
rect 8570 15348 8576 15360
rect 8260 15320 8576 15348
rect 8260 15308 8266 15320
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 12894 15348 12900 15360
rect 10192 15320 12900 15348
rect 10192 15308 10198 15320
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 15856 15348 15884 15388
rect 16776 15388 19073 15416
rect 16776 15348 16804 15388
rect 19061 15385 19073 15388
rect 19107 15385 19119 15419
rect 19061 15379 19119 15385
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 19812 15416 19840 15447
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 20346 15484 20352 15496
rect 20036 15456 20352 15484
rect 20036 15444 20042 15456
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 19484 15388 19840 15416
rect 19484 15376 19490 15388
rect 15856 15320 16804 15348
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18012 15320 18245 15348
rect 18012 15308 18018 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15348 19303 15351
rect 19978 15348 19984 15360
rect 19291 15320 19984 15348
rect 19291 15317 19303 15320
rect 19245 15311 19303 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20438 15348 20444 15360
rect 20399 15320 20444 15348
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 1946 15144 1952 15156
rect 1907 15116 1952 15144
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 4246 15144 4252 15156
rect 3528 15116 4252 15144
rect 3528 15017 3556 15116
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 8202 15144 8208 15156
rect 7024 15116 8208 15144
rect 7024 15017 7052 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8444 15116 8677 15144
rect 8444 15104 8450 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 16945 15147 17003 15153
rect 13136 15116 14964 15144
rect 13136 15104 13142 15116
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 9582 15008 9588 15020
rect 9355 14980 9588 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 14936 15008 14964 15116
rect 16945 15113 16957 15147
rect 16991 15144 17003 15147
rect 18506 15144 18512 15156
rect 16991 15116 18512 15144
rect 16991 15113 17003 15116
rect 16945 15107 17003 15113
rect 18506 15104 18512 15116
rect 18564 15104 18570 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18877 15147 18935 15153
rect 18877 15144 18889 15147
rect 18748 15116 18889 15144
rect 18748 15104 18754 15116
rect 18877 15113 18889 15116
rect 18923 15113 18935 15147
rect 18877 15107 18935 15113
rect 19168 15116 20760 15144
rect 19168 15076 19196 15116
rect 17144 15048 19196 15076
rect 14936 14980 15240 15008
rect 7282 14949 7288 14952
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 7276 14940 7288 14949
rect 1811 14912 5212 14940
rect 7243 14912 7288 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 3786 14881 3792 14884
rect 3780 14872 3792 14881
rect 3747 14844 3792 14872
rect 3780 14835 3792 14844
rect 3786 14832 3792 14835
rect 3844 14832 3850 14884
rect 5184 14872 5212 14912
rect 7276 14903 7288 14912
rect 7282 14900 7288 14903
rect 7340 14900 7346 14952
rect 12802 14940 12808 14952
rect 12763 14912 12808 14940
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 15010 14940 15016 14952
rect 13495 14912 15016 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 15010 14900 15016 14912
rect 15068 14940 15074 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 15068 14912 15117 14940
rect 15068 14900 15074 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15212 14940 15240 14980
rect 17144 14940 17172 15048
rect 19242 15036 19248 15088
rect 19300 15036 19306 15088
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17276 14980 17509 15008
rect 17276 14968 17282 14980
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 18598 15008 18604 15020
rect 18463 14980 18604 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19260 15008 19288 15036
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 19260 14980 19441 15008
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 15212 14912 17172 14940
rect 17313 14943 17371 14949
rect 15105 14903 15163 14909
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17954 14940 17960 14952
rect 17359 14912 17960 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 19058 14900 19064 14952
rect 19116 14900 19122 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14940 19303 14943
rect 19334 14940 19340 14952
rect 19291 14912 19340 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20732 14949 20760 15116
rect 20717 14943 20775 14949
rect 20717 14909 20729 14943
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 7558 14872 7564 14884
rect 5184 14844 7564 14872
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 9033 14875 9091 14881
rect 9033 14841 9045 14875
rect 9079 14872 9091 14875
rect 10134 14872 10140 14884
rect 9079 14844 10140 14872
rect 9079 14841 9091 14844
rect 9033 14835 9091 14841
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 13722 14881 13728 14884
rect 13716 14872 13728 14881
rect 13683 14844 13728 14872
rect 13716 14835 13728 14844
rect 13722 14832 13728 14835
rect 13780 14832 13786 14884
rect 15350 14875 15408 14881
rect 15350 14872 15362 14875
rect 15120 14844 15362 14872
rect 15120 14816 15148 14844
rect 15350 14841 15362 14844
rect 15396 14841 15408 14875
rect 19076 14872 19104 14900
rect 19702 14872 19708 14884
rect 19076 14844 19708 14872
rect 15350 14835 15408 14841
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 20254 14872 20260 14884
rect 20215 14844 20260 14872
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 2740 14776 4905 14804
rect 2740 14764 2746 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8352 14776 8401 14804
rect 8352 14764 8358 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8389 14767 8447 14773
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8536 14776 9137 14804
rect 8536 14764 8542 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 12618 14804 12624 14816
rect 12579 14776 12624 14804
rect 9125 14767 9183 14773
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 14829 14807 14887 14813
rect 14829 14773 14841 14807
rect 14875 14804 14887 14807
rect 15102 14804 15108 14816
rect 14875 14776 15108 14804
rect 14875 14773 14887 14776
rect 14829 14767 14887 14773
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16485 14807 16543 14813
rect 16485 14804 16497 14807
rect 16448 14776 16497 14804
rect 16448 14764 16454 14776
rect 16485 14773 16497 14776
rect 16531 14773 16543 14807
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 16485 14767 16543 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19116 14776 19349 14804
rect 19116 14764 19122 14776
rect 19337 14773 19349 14776
rect 19383 14804 19395 14807
rect 19794 14804 19800 14816
rect 19383 14776 19800 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 20898 14804 20904 14816
rect 20859 14776 20904 14804
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6972 14572 7021 14600
rect 6972 14560 6978 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 15010 14600 15016 14612
rect 14967 14572 15016 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 15010 14560 15016 14572
rect 15068 14600 15074 14612
rect 15378 14600 15384 14612
rect 15068 14572 15384 14600
rect 15068 14560 15074 14572
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 17589 14603 17647 14609
rect 17589 14569 17601 14603
rect 17635 14600 17647 14603
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17635 14572 18153 14600
rect 17635 14569 17647 14572
rect 17589 14563 17647 14569
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 18141 14563 18199 14569
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 5620 14535 5678 14541
rect 5620 14501 5632 14535
rect 5666 14532 5678 14535
rect 6086 14532 6092 14544
rect 5666 14504 6092 14532
rect 5666 14501 5678 14504
rect 5620 14495 5678 14501
rect 6086 14492 6092 14504
rect 6144 14532 6150 14544
rect 7742 14532 7748 14544
rect 6144 14504 7748 14532
rect 6144 14492 6150 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 10612 14504 12081 14532
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 1728 14436 1777 14464
rect 1728 14424 1734 14436
rect 1765 14433 1777 14436
rect 1811 14433 1823 14467
rect 1765 14427 1823 14433
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2188 14436 2973 14464
rect 2188 14424 2194 14436
rect 2961 14433 2973 14436
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 5350 14464 5356 14476
rect 4856 14436 5356 14464
rect 4856 14424 4862 14436
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14464 7435 14467
rect 8386 14464 8392 14476
rect 7423 14436 8392 14464
rect 7423 14433 7435 14436
rect 7377 14427 7435 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 10612 14473 10640 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 12802 14492 12808 14544
rect 12860 14532 12866 14544
rect 13538 14532 13544 14544
rect 12860 14504 13544 14532
rect 12860 14492 12866 14504
rect 13538 14492 13544 14504
rect 13596 14532 13602 14544
rect 13596 14504 15148 14532
rect 13596 14492 13602 14504
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14433 10655 14467
rect 10597 14427 10655 14433
rect 10864 14467 10922 14473
rect 10864 14433 10876 14467
rect 10910 14464 10922 14467
rect 11882 14464 11888 14476
rect 10910 14436 11888 14464
rect 10910 14433 10922 14436
rect 10864 14427 10922 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12520 14467 12578 14473
rect 12520 14464 12532 14467
rect 11992 14436 12532 14464
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7469 14399 7527 14405
rect 7469 14396 7481 14399
rect 6880 14368 7481 14396
rect 6880 14356 6886 14368
rect 7469 14365 7481 14368
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 10502 14396 10508 14408
rect 9171 14368 10508 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 6288 14300 6868 14328
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 2590 14260 2596 14272
rect 2551 14232 2596 14260
rect 2590 14220 2596 14232
rect 2648 14220 2654 14272
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 6288 14260 6316 14300
rect 6730 14260 6736 14272
rect 3936 14232 6316 14260
rect 6691 14232 6736 14260
rect 3936 14220 3942 14232
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 6840 14260 6868 14300
rect 7282 14288 7288 14340
rect 7340 14328 7346 14340
rect 7576 14328 7604 14359
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11992 14337 12020 14436
rect 12520 14433 12532 14436
rect 12566 14464 12578 14467
rect 13446 14464 13452 14476
rect 12566 14436 13452 14464
rect 12566 14433 12578 14436
rect 12520 14427 12578 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 14274 14464 14280 14476
rect 14235 14436 14280 14464
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 15120 14473 15148 14504
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 17494 14464 17500 14476
rect 17455 14436 17500 14464
rect 15105 14427 15163 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 18506 14464 18512 14476
rect 18467 14436 18512 14464
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20254 14464 20260 14476
rect 20215 14436 20260 14464
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12115 14368 12265 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 14366 14396 14372 14408
rect 14327 14368 14372 14396
rect 12253 14359 12311 14365
rect 7340 14300 7604 14328
rect 11977 14331 12035 14337
rect 7340 14288 7346 14300
rect 11977 14297 11989 14331
rect 12023 14297 12035 14331
rect 11977 14291 12035 14297
rect 10594 14260 10600 14272
rect 6840 14232 10600 14260
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 12268 14260 12296 14359
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 13633 14331 13691 14337
rect 13633 14297 13645 14331
rect 13679 14328 13691 14331
rect 13722 14328 13728 14340
rect 13679 14300 13728 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 13722 14288 13728 14300
rect 13780 14328 13786 14340
rect 14476 14328 14504 14359
rect 17218 14356 17224 14408
rect 17276 14396 17282 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17276 14368 17693 14396
rect 17276 14356 17282 14368
rect 17681 14365 17693 14368
rect 17727 14365 17739 14399
rect 18598 14396 18604 14408
rect 18559 14368 18604 14396
rect 17681 14359 17739 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 18748 14368 18793 14396
rect 18748 14356 18754 14368
rect 13780 14300 14504 14328
rect 17129 14331 17187 14337
rect 13780 14288 13786 14300
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 18874 14328 18880 14340
rect 17175 14300 18880 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 12618 14260 12624 14272
rect 12268 14232 12624 14260
rect 12618 14220 12624 14232
rect 12676 14260 12682 14272
rect 13170 14260 13176 14272
rect 12676 14232 13176 14260
rect 12676 14220 12682 14232
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13909 14263 13967 14269
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 14826 14260 14832 14272
rect 13955 14232 14832 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 16850 14220 16856 14272
rect 16908 14260 16914 14272
rect 19426 14260 19432 14272
rect 16908 14232 19432 14260
rect 16908 14220 16914 14232
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 20438 14260 20444 14272
rect 20399 14232 20444 14260
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2130 14056 2136 14068
rect 2091 14028 2136 14056
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 3108 14028 3893 14056
rect 3108 14016 3114 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5408 14028 6009 14056
rect 5408 14016 5414 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 5997 14019 6055 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7190 14056 7196 14068
rect 6972 14028 7196 14056
rect 6972 14016 6978 14028
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8478 14056 8484 14068
rect 8159 14028 8484 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8996 14028 9137 14056
rect 8996 14016 9002 14028
rect 9125 14025 9137 14028
rect 9171 14025 9183 14059
rect 9125 14019 9183 14025
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 9950 14056 9956 14068
rect 9640 14028 9956 14056
rect 9640 14016 9646 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10134 14056 10140 14068
rect 10095 14028 10140 14056
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 14274 14056 14280 14068
rect 14235 14028 14280 14056
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 14884 14028 17080 14056
rect 14884 14016 14890 14028
rect 3326 13988 3332 14000
rect 3287 13960 3332 13988
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 8294 13948 8300 14000
rect 8352 13988 8358 14000
rect 11241 13991 11299 13997
rect 8352 13960 9812 13988
rect 8352 13948 8358 13960
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2682 13880 2688 13892
rect 2740 13920 2746 13932
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 2740 13892 4445 13920
rect 2740 13880 2746 13892
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4433 13883 4491 13889
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 8772 13929 8800 13960
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 6788 13892 7481 13920
rect 6788 13880 6794 13892
rect 7469 13889 7481 13892
rect 7515 13920 7527 13923
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 7515 13892 8033 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8021 13889 8033 13892
rect 8067 13889 8079 13923
rect 8021 13883 8079 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9784 13929 9812 13960
rect 11241 13957 11253 13991
rect 11287 13988 11299 13991
rect 11287 13960 14780 13988
rect 11287 13957 11299 13960
rect 11241 13951 11299 13957
rect 9769 13923 9827 13929
rect 9272 13892 9352 13920
rect 9272 13880 9278 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2590 13852 2596 13864
rect 1443 13824 2596 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 6086 13852 6092 13864
rect 3191 13824 6092 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 7098 13852 7104 13864
rect 6227 13824 7104 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 9324 13852 9352 13892
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10226 13920 10232 13932
rect 9815 13892 10232 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 10284 13892 10701 13920
rect 10284 13880 10290 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 11882 13920 11888 13932
rect 11795 13892 11888 13920
rect 10689 13883 10747 13889
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 11940 13892 13921 13920
rect 11940 13880 11946 13892
rect 13909 13889 13921 13892
rect 13955 13920 13967 13923
rect 14090 13920 14096 13932
rect 13955 13892 14096 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14752 13929 14780 13960
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9324 13824 9505 13852
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 14936 13852 14964 13883
rect 9493 13815 9551 13821
rect 13280 13824 14688 13852
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 8481 13787 8539 13793
rect 8481 13784 8493 13787
rect 6328 13756 8493 13784
rect 6328 13744 6334 13756
rect 8481 13753 8493 13756
rect 8527 13753 8539 13787
rect 8481 13747 8539 13753
rect 8573 13787 8631 13793
rect 8573 13753 8585 13787
rect 8619 13784 8631 13787
rect 9398 13784 9404 13796
rect 8619 13756 9404 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 10502 13784 10508 13796
rect 10463 13756 10508 13784
rect 10502 13744 10508 13756
rect 10560 13744 10566 13796
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 10652 13756 10697 13784
rect 10796 13756 11744 13784
rect 10652 13744 10658 13756
rect 2222 13676 2228 13728
rect 2280 13716 2286 13728
rect 2501 13719 2559 13725
rect 2501 13716 2513 13719
rect 2280 13688 2513 13716
rect 2280 13676 2286 13688
rect 2501 13685 2513 13688
rect 2547 13685 2559 13719
rect 2501 13679 2559 13685
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 4246 13716 4252 13728
rect 2648 13688 2693 13716
rect 4207 13688 4252 13716
rect 2648 13676 2654 13688
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 7190 13716 7196 13728
rect 4396 13688 4441 13716
rect 7151 13688 7196 13716
rect 4396 13676 4402 13688
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 8021 13719 8079 13725
rect 7340 13688 7385 13716
rect 7340 13676 7346 13688
rect 8021 13685 8033 13719
rect 8067 13716 8079 13719
rect 8938 13716 8944 13728
rect 8067 13688 8944 13716
rect 8067 13685 8079 13688
rect 8021 13679 8079 13685
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9364 13688 9597 13716
rect 9364 13676 9370 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9585 13679 9643 13685
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10796 13716 10824 13756
rect 11606 13716 11612 13728
rect 9732 13688 10824 13716
rect 11567 13688 11612 13716
rect 9732 13676 9738 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11716 13725 11744 13756
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 11790 13716 11796 13728
rect 11747 13688 11796 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 13280 13725 13308 13824
rect 13446 13744 13452 13796
rect 13504 13784 13510 13796
rect 14660 13793 14688 13824
rect 14844 13824 14964 13852
rect 15289 13855 15347 13861
rect 14645 13787 14703 13793
rect 13504 13756 13952 13784
rect 13504 13744 13510 13756
rect 13265 13719 13323 13725
rect 13265 13685 13277 13719
rect 13311 13685 13323 13719
rect 13630 13716 13636 13728
rect 13591 13688 13636 13716
rect 13265 13679 13323 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13725 13719 13783 13725
rect 13725 13685 13737 13719
rect 13771 13716 13783 13719
rect 13814 13716 13820 13728
rect 13771 13688 13820 13716
rect 13771 13685 13783 13688
rect 13725 13679 13783 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 13924 13716 13952 13756
rect 14645 13753 14657 13787
rect 14691 13753 14703 13787
rect 14645 13747 14703 13753
rect 14844 13716 14872 13824
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15378 13852 15384 13864
rect 15335 13824 15384 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15556 13855 15614 13861
rect 15556 13821 15568 13855
rect 15602 13852 15614 13855
rect 16942 13852 16948 13864
rect 15602 13824 16948 13852
rect 15602 13821 15614 13824
rect 15556 13815 15614 13821
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 17052 13852 17080 14028
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 18785 14059 18843 14065
rect 18785 14056 18797 14059
rect 18656 14028 18797 14056
rect 18656 14016 18662 14028
rect 18785 14025 18797 14028
rect 18831 14025 18843 14059
rect 18785 14019 18843 14025
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20993 13991 21051 13997
rect 20993 13988 21005 13991
rect 20680 13960 21005 13988
rect 20680 13948 20686 13960
rect 20993 13957 21005 13960
rect 21039 13957 21051 13991
rect 20993 13951 21051 13957
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19242 13920 19248 13932
rect 19116 13892 19248 13920
rect 19116 13880 19122 13892
rect 19242 13880 19248 13892
rect 19300 13920 19306 13932
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 19300 13892 19349 13920
rect 19300 13880 19306 13892
rect 19337 13889 19349 13892
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 17052 13824 20085 13852
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20395 13824 20821 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 19702 13784 19708 13796
rect 15068 13756 19708 13784
rect 15068 13744 15074 13756
rect 19702 13744 19708 13756
rect 19760 13744 19766 13796
rect 13924 13688 14872 13716
rect 16114 13676 16120 13728
rect 16172 13716 16178 13728
rect 16669 13719 16727 13725
rect 16669 13716 16681 13719
rect 16172 13688 16681 13716
rect 16172 13676 16178 13688
rect 16669 13685 16681 13688
rect 16715 13685 16727 13719
rect 16669 13679 16727 13685
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 19153 13719 19211 13725
rect 19153 13716 19165 13719
rect 17092 13688 19165 13716
rect 17092 13676 17098 13688
rect 19153 13685 19165 13688
rect 19199 13685 19211 13719
rect 19153 13679 19211 13685
rect 19245 13719 19303 13725
rect 19245 13685 19257 13719
rect 19291 13716 19303 13719
rect 19426 13716 19432 13728
rect 19291 13688 19432 13716
rect 19291 13685 19303 13688
rect 19245 13679 19303 13685
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2222 13512 2228 13524
rect 2183 13484 2228 13512
rect 2222 13472 2228 13484
rect 2280 13472 2286 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4396 13484 4537 13512
rect 4396 13472 4402 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 4525 13475 4583 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7392 13484 7757 13512
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 7392 13444 7420 13484
rect 7745 13481 7757 13484
rect 7791 13512 7803 13515
rect 9674 13512 9680 13524
rect 7791 13484 9680 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 9999 13484 13185 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 13630 13472 13636 13524
rect 13688 13512 13694 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13688 13484 13829 13512
rect 13688 13472 13694 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 16485 13515 16543 13521
rect 16485 13512 16497 13515
rect 15887 13484 16497 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 16485 13481 16497 13484
rect 16531 13481 16543 13515
rect 16485 13475 16543 13481
rect 16758 13472 16764 13524
rect 16816 13512 16822 13524
rect 17218 13512 17224 13524
rect 16816 13484 17224 13512
rect 16816 13472 16822 13484
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 17552 13484 17693 13512
rect 17552 13472 17558 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 17681 13475 17739 13481
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18564 13484 18705 13512
rect 18564 13472 18570 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18693 13475 18751 13481
rect 9858 13444 9864 13456
rect 2924 13416 7420 13444
rect 7668 13416 9864 13444
rect 2924 13404 2930 13416
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 3237 13379 3295 13385
rect 3237 13376 3249 13379
rect 2639 13348 3249 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 3237 13345 3249 13348
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 4893 13379 4951 13385
rect 4893 13345 4905 13379
rect 4939 13376 4951 13379
rect 5534 13376 5540 13388
rect 4939 13348 5540 13376
rect 4939 13345 4951 13348
rect 4893 13339 4951 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7668 13385 7696 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 15010 13444 15016 13456
rect 11664 13416 15016 13444
rect 11664 13404 11670 13416
rect 15010 13404 15016 13416
rect 15068 13404 15074 13456
rect 16853 13447 16911 13453
rect 16853 13413 16865 13447
rect 16899 13444 16911 13447
rect 16899 13416 18552 13444
rect 16899 13413 16911 13416
rect 16853 13407 16911 13413
rect 18524 13388 18552 13416
rect 7653 13379 7711 13385
rect 7653 13376 7665 13379
rect 6880 13348 7665 13376
rect 6880 13336 6886 13348
rect 7653 13345 7665 13348
rect 7699 13345 7711 13379
rect 7653 13339 7711 13345
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 10321 13379 10379 13385
rect 10321 13376 10333 13379
rect 9272 13348 10333 13376
rect 9272 13336 9278 13348
rect 10321 13345 10333 13348
rect 10367 13345 10379 13379
rect 10321 13339 10379 13345
rect 13188 13348 13584 13376
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2464 13280 2697 13308
rect 2464 13268 2470 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 2958 13308 2964 13320
rect 2915 13280 2964 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 4982 13308 4988 13320
rect 4943 13280 4988 13308
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 2976 13240 3004 13268
rect 3786 13240 3792 13252
rect 2976 13212 3792 13240
rect 3786 13200 3792 13212
rect 3844 13240 3850 13252
rect 5092 13240 5120 13271
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 7892 13280 7937 13308
rect 7892 13268 7898 13280
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 9364 13280 10425 13308
rect 9364 13268 9370 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 11882 13308 11888 13320
rect 10643 13280 11888 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 13188 13240 13216 13348
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 13265 13271 13323 13277
rect 3844 13212 5120 13240
rect 6932 13212 13216 13240
rect 13280 13240 13308 13271
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13556 13308 13584 13348
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14148 13348 16160 13376
rect 14148 13336 14154 13348
rect 16132 13320 16160 13348
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 18049 13379 18107 13385
rect 18049 13376 18061 13379
rect 18012 13348 18061 13376
rect 18012 13336 18018 13348
rect 18049 13345 18061 13348
rect 18095 13345 18107 13379
rect 18049 13339 18107 13345
rect 18506 13336 18512 13388
rect 18564 13336 18570 13388
rect 18874 13336 18880 13388
rect 18932 13376 18938 13388
rect 19061 13379 19119 13385
rect 19061 13376 19073 13379
rect 18932 13348 19073 13376
rect 18932 13336 18938 13348
rect 19061 13345 19073 13348
rect 19107 13345 19119 13379
rect 19061 13339 19119 13345
rect 15378 13308 15384 13320
rect 13556 13280 15384 13308
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16114 13308 16120 13320
rect 16075 13280 16120 13308
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 16942 13308 16948 13320
rect 16903 13280 16948 13308
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17920 13280 18153 13308
rect 17920 13268 17926 13280
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18690 13308 18696 13320
rect 18279 13280 18696 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 13280 13212 15485 13240
rect 3844 13200 3850 13212
rect 5074 13132 5080 13184
rect 5132 13172 5138 13184
rect 6932 13172 6960 13212
rect 15473 13209 15485 13212
rect 15519 13209 15531 13243
rect 15473 13203 15531 13209
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 18248 13240 18276 13271
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 19153 13311 19211 13317
rect 19153 13308 19165 13311
rect 18892 13280 19165 13308
rect 16448 13212 18276 13240
rect 16448 13200 16454 13212
rect 5132 13144 6960 13172
rect 5132 13132 5138 13144
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 8294 13172 8300 13184
rect 7432 13144 8300 13172
rect 7432 13132 7438 13144
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 12805 13175 12863 13181
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 14366 13172 14372 13184
rect 12851 13144 14372 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 16574 13172 16580 13184
rect 14516 13144 16580 13172
rect 14516 13132 14522 13144
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 18892 13172 18920 13280
rect 19153 13277 19165 13280
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 19260 13240 19288 13271
rect 19116 13212 19288 13240
rect 19116 13200 19122 13212
rect 16816 13144 18920 13172
rect 16816 13132 16822 13144
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2406 12968 2412 12980
rect 2367 12940 2412 12968
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 7098 12968 7104 12980
rect 7059 12940 7104 12968
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 14458 12968 14464 12980
rect 12483 12940 14464 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16485 12971 16543 12977
rect 16485 12968 16497 12971
rect 15988 12940 16497 12968
rect 15988 12928 15994 12940
rect 16485 12937 16497 12940
rect 16531 12937 16543 12971
rect 16485 12931 16543 12937
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16632 12940 17540 12968
rect 16632 12928 16638 12940
rect 7377 12903 7435 12909
rect 7377 12869 7389 12903
rect 7423 12900 7435 12903
rect 14277 12903 14335 12909
rect 7423 12872 8892 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 3050 12832 3056 12844
rect 3011 12804 3056 12832
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5316 12804 5457 12832
rect 5316 12792 5322 12804
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5445 12795 5503 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 6178 12792 6184 12844
rect 6236 12832 6242 12844
rect 7926 12832 7932 12844
rect 6236 12804 7788 12832
rect 7887 12804 7932 12832
rect 6236 12792 6242 12804
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 3142 12764 3148 12776
rect 2823 12736 3148 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 3142 12724 3148 12736
rect 3200 12764 3206 12776
rect 3418 12764 3424 12776
rect 3200 12736 3424 12764
rect 3200 12724 3206 12736
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 5074 12724 5080 12776
rect 5132 12764 5138 12776
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 5132 12736 5365 12764
rect 5132 12724 5138 12736
rect 5353 12733 5365 12736
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 7760 12773 7788 12804
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 8202 12832 8208 12844
rect 7984 12804 8208 12832
rect 7984 12792 7990 12804
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8864 12841 8892 12872
rect 14277 12869 14289 12903
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 15289 12903 15347 12909
rect 15289 12869 15301 12903
rect 15335 12900 15347 12903
rect 17402 12900 17408 12912
rect 15335 12872 17408 12900
rect 15335 12869 15347 12872
rect 15289 12863 15347 12869
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 12158 12832 12164 12844
rect 8996 12804 9041 12832
rect 10612 12804 12164 12832
rect 8996 12792 9002 12804
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 7156 12736 7297 12764
rect 7156 12724 7162 12736
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 10612 12764 10640 12804
rect 12158 12792 12164 12804
rect 12216 12832 12222 12844
rect 13081 12835 13139 12841
rect 12216 12804 13032 12832
rect 12216 12792 12222 12804
rect 7883 12736 10640 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 12452 12696 12480 12724
rect 4120 12668 12480 12696
rect 4120 12656 4126 12668
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12584 12668 12909 12696
rect 12584 12656 12590 12668
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 13004 12696 13032 12804
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13446 12832 13452 12844
rect 13127 12804 13452 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 13814 12764 13820 12776
rect 13775 12736 13820 12764
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14292 12764 14320 12863
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 17512 12900 17540 12940
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 17920 12940 18337 12968
rect 17920 12928 17926 12940
rect 18325 12937 18337 12940
rect 18371 12937 18383 12971
rect 18325 12931 18383 12937
rect 20346 12928 20352 12980
rect 20404 12928 20410 12980
rect 20364 12900 20392 12928
rect 17512 12872 20392 12900
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12832 14979 12835
rect 15102 12832 15108 12844
rect 14967 12804 15108 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16390 12832 16396 12844
rect 15979 12804 16396 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 18748 12804 18981 12832
rect 18748 12792 18754 12804
rect 18969 12801 18981 12804
rect 19015 12832 19027 12835
rect 19058 12832 19064 12844
rect 19015 12804 19064 12832
rect 19015 12801 19027 12804
rect 18969 12795 19027 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 20404 12804 20821 12832
rect 20404 12792 20410 12804
rect 20809 12801 20821 12804
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 14292 12736 15669 12764
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 18874 12764 18880 12776
rect 16899 12736 18880 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20714 12764 20720 12776
rect 19852 12736 20720 12764
rect 19852 12724 19858 12736
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 14645 12699 14703 12705
rect 14645 12696 14657 12699
rect 13004 12668 14657 12696
rect 12897 12659 12955 12665
rect 14645 12665 14657 12668
rect 14691 12665 14703 12699
rect 14645 12659 14703 12665
rect 16945 12699 17003 12705
rect 16945 12665 16957 12699
rect 16991 12696 17003 12699
rect 17034 12696 17040 12708
rect 16991 12668 17040 12696
rect 16991 12665 17003 12668
rect 16945 12659 17003 12665
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 17586 12656 17592 12708
rect 17644 12696 17650 12708
rect 20622 12696 20628 12708
rect 17644 12668 18828 12696
rect 20583 12668 20628 12696
rect 17644 12656 17650 12668
rect 18800 12640 18828 12668
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 2869 12631 2927 12637
rect 2869 12597 2881 12631
rect 2915 12628 2927 12631
rect 6638 12628 6644 12640
rect 2915 12600 6644 12628
rect 2915 12597 2927 12600
rect 2869 12591 2927 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 8754 12628 8760 12640
rect 8715 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 11333 12631 11391 12637
rect 11333 12597 11345 12631
rect 11379 12628 11391 12631
rect 11882 12628 11888 12640
rect 11379 12600 11888 12628
rect 11379 12597 11391 12600
rect 11333 12591 11391 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12802 12628 12808 12640
rect 12763 12600 12808 12628
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 13538 12588 13544 12640
rect 13596 12628 13602 12640
rect 13633 12631 13691 12637
rect 13633 12628 13645 12631
rect 13596 12600 13645 12628
rect 13596 12588 13602 12600
rect 13633 12597 13645 12600
rect 13679 12597 13691 12631
rect 13633 12591 13691 12597
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 13964 12600 14749 12628
rect 13964 12588 13970 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 15804 12600 15849 12628
rect 15804 12588 15810 12600
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 18693 12631 18751 12637
rect 18693 12628 18705 12631
rect 17828 12600 18705 12628
rect 17828 12588 17834 12600
rect 18693 12597 18705 12600
rect 18739 12597 18751 12631
rect 18693 12591 18751 12597
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 20254 12628 20260 12640
rect 18840 12600 18885 12628
rect 20215 12600 20260 12628
rect 18840 12588 18846 12600
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2590 12424 2596 12436
rect 2271 12396 2596 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 5902 12384 5908 12436
rect 5960 12424 5966 12436
rect 6270 12424 6276 12436
rect 5960 12396 6276 12424
rect 5960 12384 5966 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7248 12396 7573 12424
rect 7248 12384 7254 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 10962 12424 10968 12436
rect 7561 12387 7619 12393
rect 7944 12396 10968 12424
rect 2590 12288 2596 12300
rect 2551 12260 2596 12288
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5166 12288 5172 12300
rect 4764 12260 5172 12288
rect 4764 12248 4770 12260
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5307 12260 5764 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2556 12192 2697 12220
rect 2556 12180 2562 12192
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 2958 12220 2964 12232
rect 2915 12192 2964 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2958 12180 2964 12192
rect 3016 12220 3022 12232
rect 3694 12220 3700 12232
rect 3016 12192 3700 12220
rect 3016 12180 3022 12192
rect 3694 12180 3700 12192
rect 3752 12180 3758 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5626 12220 5632 12232
rect 5399 12192 5632 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 5368 12152 5396 12183
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 3108 12124 5396 12152
rect 5736 12152 5764 12260
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 5960 12260 6193 12288
rect 5960 12248 5966 12260
rect 6181 12257 6193 12260
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7944 12297 7972 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 11195 12396 12449 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 12437 12393 12449 12396
rect 12483 12393 12495 12427
rect 12437 12387 12495 12393
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15746 12424 15752 12436
rect 15335 12396 15752 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17770 12424 17776 12436
rect 17000 12396 17776 12424
rect 17000 12384 17006 12396
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 18012 12396 18153 12424
rect 18012 12384 18018 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18506 12424 18512 12436
rect 18419 12396 18512 12424
rect 18141 12387 18199 12393
rect 18506 12384 18512 12396
rect 18564 12424 18570 12436
rect 18564 12396 19104 12424
rect 18564 12384 18570 12396
rect 19076 12368 19104 12396
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 11238 12356 11244 12368
rect 8720 12328 11244 12356
rect 8720 12316 8726 12328
rect 11238 12316 11244 12328
rect 11296 12316 11302 12368
rect 12066 12356 12072 12368
rect 11440 12328 12072 12356
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 6972 12260 7941 12288
rect 6972 12248 6978 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 9677 12291 9735 12297
rect 9677 12288 9689 12291
rect 8628 12260 9689 12288
rect 8628 12248 8634 12260
rect 9677 12257 9689 12260
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 9933 12291 9991 12297
rect 9933 12288 9945 12291
rect 9824 12260 9945 12288
rect 9824 12248 9830 12260
rect 9933 12257 9945 12260
rect 9979 12288 9991 12291
rect 11440 12288 11468 12328
rect 9979 12260 11468 12288
rect 9979 12257 9991 12260
rect 9933 12251 9991 12257
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11572 12260 11617 12288
rect 11572 12248 11578 12260
rect 6270 12220 6276 12232
rect 6231 12192 6276 12220
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 7101 12223 7159 12229
rect 6420 12192 6465 12220
rect 6420 12180 6426 12192
rect 7101 12189 7113 12223
rect 7147 12220 7159 12223
rect 7466 12220 7472 12232
rect 7147 12192 7472 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7708 12192 8033 12220
rect 7708 12180 7714 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 8021 12183 8079 12189
rect 8036 12152 8064 12183
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11716 12229 11744 12328
rect 12066 12316 12072 12328
rect 12124 12356 12130 12368
rect 12124 12328 14596 12356
rect 12124 12316 12130 12328
rect 12342 12288 12348 12300
rect 12303 12260 12348 12288
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 12710 12288 12716 12300
rect 12492 12260 12716 12288
rect 12492 12248 12498 12260
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 13446 12297 13452 12300
rect 13440 12288 13452 12297
rect 13407 12260 13452 12288
rect 13440 12251 13452 12260
rect 13446 12248 13452 12251
rect 13504 12248 13510 12300
rect 14568 12288 14596 12328
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 18690 12356 18696 12368
rect 15252 12328 18696 12356
rect 15252 12316 15258 12328
rect 15286 12288 15292 12300
rect 14568 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11020 12192 11621 12220
rect 11020 12180 11026 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12189 11759 12223
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 11701 12183 11759 12189
rect 11808 12192 12541 12220
rect 8846 12152 8852 12164
rect 5736 12124 7420 12152
rect 8036 12124 8852 12152
rect 3108 12112 3114 12124
rect 4798 12084 4804 12096
rect 4759 12056 4804 12084
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5810 12084 5816 12096
rect 5771 12056 5816 12084
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7282 12084 7288 12096
rect 7064 12056 7288 12084
rect 7064 12044 7070 12056
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7392 12084 7420 12124
rect 8846 12112 8852 12124
rect 8904 12112 8910 12164
rect 11057 12155 11115 12161
rect 11057 12121 11069 12155
rect 11103 12152 11115 12155
rect 11808 12152 11836 12192
rect 12529 12189 12541 12192
rect 12575 12220 12587 12223
rect 12986 12220 12992 12232
rect 12575 12192 12992 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13170 12220 13176 12232
rect 13131 12192 13176 12220
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 15856 12229 15884 12328
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 19058 12316 19064 12368
rect 19116 12316 19122 12368
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 11103 12124 11836 12152
rect 11977 12155 12035 12161
rect 11103 12121 11115 12124
rect 11057 12115 11115 12121
rect 11977 12121 11989 12155
rect 12023 12152 12035 12155
rect 12802 12152 12808 12164
rect 12023 12124 12808 12152
rect 12023 12121 12035 12124
rect 11977 12115 12035 12121
rect 12802 12112 12808 12124
rect 12860 12112 12866 12164
rect 15764 12152 15792 12183
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 18708 12229 18736 12316
rect 19420 12291 19478 12297
rect 19420 12257 19432 12291
rect 19466 12288 19478 12291
rect 20346 12288 20352 12300
rect 19466 12260 20352 12288
rect 19466 12257 19478 12260
rect 19420 12251 19478 12257
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 17736 12192 18613 12220
rect 17736 12180 17742 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 19153 12223 19211 12229
rect 19153 12220 19165 12223
rect 18932 12192 19165 12220
rect 18932 12180 18938 12192
rect 19153 12189 19165 12192
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 16022 12152 16028 12164
rect 14384 12124 14780 12152
rect 15764 12124 16028 12152
rect 10962 12084 10968 12096
rect 7392 12056 10968 12084
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 14384 12084 14412 12124
rect 14550 12084 14556 12096
rect 11664 12056 14412 12084
rect 14511 12056 14556 12084
rect 11664 12044 11670 12056
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14752 12084 14780 12124
rect 16022 12112 16028 12124
rect 16080 12112 16086 12164
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18892 12152 18920 12180
rect 17920 12124 18920 12152
rect 17920 12112 17926 12124
rect 20162 12084 20168 12096
rect 14752 12056 20168 12084
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20530 12084 20536 12096
rect 20491 12056 20536 12084
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 4154 11880 4160 11892
rect 2332 11852 4160 11880
rect 2332 11753 2360 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4304 11852 4353 11880
rect 4304 11840 4310 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 5534 11880 5540 11892
rect 5495 11852 5540 11880
rect 4341 11843 4399 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 8754 11880 8760 11892
rect 7147 11852 8760 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 10778 11880 10784 11892
rect 8904 11852 10784 11880
rect 8904 11840 8910 11852
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 12342 11880 12348 11892
rect 11563 11852 12348 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12452 11852 13400 11880
rect 3694 11812 3700 11824
rect 3607 11784 3700 11812
rect 3694 11772 3700 11784
rect 3752 11812 3758 11824
rect 3752 11784 4936 11812
rect 3752 11772 3758 11784
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 4798 11744 4804 11756
rect 4759 11716 4804 11744
rect 2317 11707 2375 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 4908 11753 4936 11784
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 8481 11815 8539 11821
rect 5040 11784 7696 11812
rect 5040 11772 5046 11784
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5684 11716 6101 11744
rect 5684 11704 5690 11716
rect 6089 11713 6101 11716
rect 6135 11744 6147 11747
rect 6362 11744 6368 11756
rect 6135 11716 6368 11744
rect 6135 11713 6147 11716
rect 6089 11707 6147 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 2584 11679 2642 11685
rect 2584 11645 2596 11679
rect 2630 11676 2642 11679
rect 3050 11676 3056 11688
rect 2630 11648 3056 11676
rect 2630 11645 2642 11648
rect 2584 11639 2642 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 5810 11676 5816 11688
rect 4755 11648 5816 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 7006 11676 7012 11688
rect 5951 11648 7012 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7466 11676 7472 11688
rect 7427 11648 7472 11676
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7668 11676 7696 11784
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 9582 11812 9588 11824
rect 8527 11784 9588 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 9861 11815 9919 11821
rect 9861 11781 9873 11815
rect 9907 11812 9919 11815
rect 11146 11812 11152 11824
rect 9907 11784 11152 11812
rect 9907 11781 9919 11784
rect 9861 11775 9919 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11744 7803 11747
rect 8202 11744 8208 11756
rect 7791 11716 8208 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9766 11744 9772 11756
rect 9171 11716 9772 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 12066 11744 12072 11756
rect 12027 11716 12072 11744
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12452 11744 12480 11852
rect 13372 11812 13400 11852
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13504 11852 13829 11880
rect 13504 11840 13510 11852
rect 13817 11849 13829 11852
rect 13863 11849 13875 11883
rect 19242 11880 19248 11892
rect 13817 11843 13875 11849
rect 18800 11852 19248 11880
rect 18800 11812 18828 11852
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 13372 11784 18828 11812
rect 12360 11716 12480 11744
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 7668 11648 10333 11676
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 11882 11676 11888 11688
rect 11843 11648 11888 11676
rect 10321 11639 10379 11645
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 4120 11580 11345 11608
rect 4120 11568 4126 11580
rect 11333 11577 11345 11580
rect 11379 11608 11391 11611
rect 11977 11611 12035 11617
rect 11977 11608 11989 11611
rect 11379 11580 11989 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 11977 11577 11989 11580
rect 12023 11608 12035 11611
rect 12360 11608 12388 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15344 11716 15945 11744
rect 15344 11704 15350 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 12444 11679 12502 11685
rect 12444 11645 12456 11679
rect 12490 11645 12502 11679
rect 12444 11639 12502 11645
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 16942 11676 16948 11688
rect 15795 11648 16948 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 12023 11580 12388 11608
rect 12023 11577 12035 11580
rect 11977 11571 12035 11577
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 4856 11512 6009 11540
rect 4856 11500 4862 11512
rect 5997 11509 6009 11512
rect 6043 11540 6055 11543
rect 6730 11540 6736 11552
rect 6043 11512 6736 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 7248 11512 7573 11540
rect 7248 11500 7254 11512
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7561 11503 7619 11509
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 7800 11512 8861 11540
rect 7800 11500 7806 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8849 11503 8907 11509
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 10226 11540 10232 11552
rect 8996 11512 9041 11540
rect 10187 11512 10232 11540
rect 8996 11500 9002 11512
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12066 11540 12072 11552
rect 11756 11512 12072 11540
rect 11756 11500 11762 11512
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12452 11540 12480 11639
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 18800 11676 18828 11784
rect 18874 11704 18880 11756
rect 18932 11744 18938 11756
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 18932 11716 18981 11744
rect 18932 11704 18938 11716
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 18800 11648 18920 11676
rect 18892 11620 18920 11648
rect 12704 11611 12762 11617
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 12986 11608 12992 11620
rect 12750 11580 12992 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 16666 11568 16672 11620
rect 16724 11608 16730 11620
rect 17586 11608 17592 11620
rect 16724 11580 17592 11608
rect 16724 11568 16730 11580
rect 17586 11568 17592 11580
rect 17644 11608 17650 11620
rect 18690 11608 18696 11620
rect 17644 11580 18696 11608
rect 17644 11568 17650 11580
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 18874 11568 18880 11620
rect 18932 11568 18938 11620
rect 19242 11617 19248 11620
rect 19236 11608 19248 11617
rect 19203 11580 19248 11608
rect 19236 11571 19248 11580
rect 19242 11568 19248 11571
rect 19300 11568 19306 11620
rect 13170 11540 13176 11552
rect 12452 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 13320 11512 15393 11540
rect 13320 11500 13326 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 15841 11543 15899 11549
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 17034 11540 17040 11552
rect 15887 11512 17040 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 17954 11500 17960 11552
rect 18012 11540 18018 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 18012 11512 18061 11540
rect 18012 11500 18018 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2498 11336 2504 11348
rect 2459 11308 2504 11336
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5215 11308 6009 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 5997 11299 6055 11305
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7156 11308 8033 11336
rect 7156 11296 7162 11308
rect 8021 11305 8033 11308
rect 8067 11336 8079 11339
rect 8202 11336 8208 11348
rect 8067 11308 8208 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9306 11336 9312 11348
rect 8904 11308 9312 11336
rect 8904 11296 8910 11308
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11336 12955 11339
rect 13262 11336 13268 11348
rect 12943 11308 13268 11336
rect 12943 11305 12955 11308
rect 12897 11299 12955 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 13814 11336 13820 11348
rect 13495 11308 13820 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 17310 11336 17316 11348
rect 15335 11308 17316 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 18656 11308 18889 11336
rect 18656 11296 18662 11308
rect 18877 11305 18889 11308
rect 18923 11305 18935 11339
rect 18877 11299 18935 11305
rect 2869 11271 2927 11277
rect 2869 11237 2881 11271
rect 2915 11268 2927 11271
rect 2958 11268 2964 11280
rect 2915 11240 2964 11268
rect 2915 11237 2927 11240
rect 2869 11231 2927 11237
rect 2958 11228 2964 11240
rect 3016 11268 3022 11280
rect 3510 11268 3516 11280
rect 3016 11240 3516 11268
rect 3016 11228 3022 11240
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 7466 11268 7472 11280
rect 5500 11240 7472 11268
rect 5500 11228 5506 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 12805 11271 12863 11277
rect 12805 11268 12817 11271
rect 9640 11240 12817 11268
rect 9640 11228 9646 11240
rect 12805 11237 12817 11240
rect 12851 11237 12863 11271
rect 12805 11231 12863 11237
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 1946 11200 1952 11212
rect 1811 11172 1952 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5718 11200 5724 11212
rect 5307 11172 5724 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7742 11200 7748 11212
rect 7156 11172 7748 11200
rect 7156 11160 7162 11172
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8251 11172 9505 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10686 11200 10692 11212
rect 10643 11172 10692 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 13633 11163 13691 11169
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2774 11064 2780 11076
rect 1995 11036 2780 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 2976 11064 3004 11095
rect 3050 11092 3056 11144
rect 3108 11132 3114 11144
rect 5442 11132 5448 11144
rect 3108 11104 3153 11132
rect 5403 11104 5448 11132
rect 3108 11092 3114 11104
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 6454 11132 6460 11144
rect 6415 11104 6460 11132
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 6604 11104 6649 11132
rect 6604 11092 6610 11104
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 6788 11104 8156 11132
rect 6788 11092 6794 11104
rect 3234 11064 3240 11076
rect 2976 11036 3240 11064
rect 3234 11024 3240 11036
rect 3292 11064 3298 11076
rect 7282 11064 7288 11076
rect 3292 11036 7288 11064
rect 3292 11024 3298 11036
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 4801 10999 4859 11005
rect 4801 10996 4813 10999
rect 4212 10968 4813 10996
rect 4212 10956 4218 10968
rect 4801 10965 4813 10968
rect 4847 10965 4859 10999
rect 4801 10959 4859 10965
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7558 10996 7564 11008
rect 7156 10968 7564 10996
rect 7156 10956 7162 10968
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 8128 10996 8156 11104
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 8444 11104 10517 11132
rect 8444 11092 8450 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 10505 11095 10563 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 9539 11036 11897 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 11885 11033 11897 11036
rect 11931 11064 11943 11067
rect 13648 11064 13676 11163
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 17494 11209 17500 11212
rect 17488 11163 17500 11209
rect 17552 11200 17558 11212
rect 17552 11172 17588 11200
rect 17494 11160 17500 11163
rect 17552 11160 17558 11172
rect 18506 11160 18512 11212
rect 18564 11200 18570 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 18564 11172 19257 11200
rect 18564 11160 18570 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 15896 11104 15941 11132
rect 15896 11092 15902 11104
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 16908 11104 17233 11132
rect 16908 11092 16914 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19337 11135 19395 11141
rect 19337 11132 19349 11135
rect 18748 11104 19349 11132
rect 18748 11092 18754 11104
rect 19337 11101 19349 11104
rect 19383 11101 19395 11135
rect 19337 11095 19395 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 11931 11036 13676 11064
rect 18601 11067 18659 11073
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 18601 11033 18613 11067
rect 18647 11064 18659 11067
rect 19242 11064 19248 11076
rect 18647 11036 19248 11064
rect 18647 11033 18659 11036
rect 18601 11027 18659 11033
rect 19242 11024 19248 11036
rect 19300 11064 19306 11076
rect 19444 11064 19472 11095
rect 19300 11036 19472 11064
rect 19300 11024 19306 11036
rect 8938 10996 8944 11008
rect 8128 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 10505 10999 10563 11005
rect 10505 10965 10517 10999
rect 10551 10996 10563 10999
rect 15470 10996 15476 11008
rect 10551 10968 15476 10996
rect 10551 10965 10563 10968
rect 10505 10959 10563 10965
rect 15470 10956 15476 10968
rect 15528 10996 15534 11008
rect 19610 10996 19616 11008
rect 15528 10968 19616 10996
rect 15528 10956 15534 10968
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2590 10792 2596 10804
rect 2547 10764 2596 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4982 10792 4988 10804
rect 4120 10764 4988 10792
rect 4120 10752 4126 10764
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5684 10764 5733 10792
rect 5684 10752 5690 10764
rect 5721 10761 5733 10764
rect 5767 10761 5779 10795
rect 5721 10755 5779 10761
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6512 10764 6837 10792
rect 6512 10752 6518 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 13906 10792 13912 10804
rect 6825 10755 6883 10761
rect 7116 10764 13912 10792
rect 1946 10656 1952 10668
rect 1907 10628 1952 10656
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 3050 10656 3056 10668
rect 3011 10628 3056 10656
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4341 10659 4399 10665
rect 4341 10656 4353 10659
rect 3844 10628 4353 10656
rect 3844 10616 3850 10628
rect 4341 10625 4353 10628
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 4154 10588 4160 10600
rect 1811 10560 4160 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 7116 10588 7144 10764
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14001 10795 14059 10801
rect 14001 10761 14013 10795
rect 14047 10792 14059 10795
rect 15654 10792 15660 10804
rect 14047 10764 15660 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18506 10792 18512 10804
rect 18095 10764 18512 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 13170 10684 13176 10736
rect 13228 10724 13234 10736
rect 14458 10724 14464 10736
rect 13228 10696 14464 10724
rect 13228 10684 13234 10696
rect 14458 10684 14464 10696
rect 14516 10724 14522 10736
rect 16945 10727 17003 10733
rect 14516 10696 15608 10724
rect 14516 10684 14522 10696
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 14550 10656 14556 10668
rect 14511 10628 14556 10656
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 15470 10656 15476 10668
rect 15431 10628 15476 10656
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15580 10665 15608 10696
rect 16945 10693 16957 10727
rect 16991 10724 17003 10727
rect 18690 10724 18696 10736
rect 16991 10696 18696 10724
rect 16991 10693 17003 10696
rect 16945 10687 17003 10693
rect 18690 10684 18696 10696
rect 18748 10684 18754 10736
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 16206 10656 16212 10668
rect 15611 10628 16212 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 17494 10656 17500 10668
rect 17455 10628 17500 10656
rect 17494 10616 17500 10628
rect 17552 10656 17558 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 17552 10628 18613 10656
rect 17552 10616 17558 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 19668 10628 20177 10656
rect 19668 10616 19674 10628
rect 20165 10625 20177 10628
rect 20211 10625 20223 10659
rect 20165 10619 20223 10625
rect 20349 10659 20407 10665
rect 20349 10625 20361 10659
rect 20395 10656 20407 10659
rect 20530 10656 20536 10668
rect 20395 10628 20536 10656
rect 20395 10625 20407 10628
rect 20349 10619 20407 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 4448 10560 7144 10588
rect 2774 10480 2780 10532
rect 2832 10520 2838 10532
rect 2869 10523 2927 10529
rect 2869 10520 2881 10523
rect 2832 10492 2881 10520
rect 2832 10480 2838 10492
rect 2869 10489 2881 10492
rect 2915 10520 2927 10523
rect 3878 10520 3884 10532
rect 2915 10492 3884 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3878 10480 3884 10492
rect 3936 10480 3942 10532
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 4448 10520 4476 10560
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10502 10597 10508 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9916 10560 10241 10588
rect 9916 10548 9922 10560
rect 10229 10557 10241 10560
rect 10275 10557 10287 10591
rect 10496 10588 10508 10597
rect 10463 10560 10508 10588
rect 10229 10551 10287 10557
rect 10496 10551 10508 10560
rect 10502 10548 10508 10551
rect 10560 10548 10566 10600
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 17402 10588 17408 10600
rect 10836 10560 16252 10588
rect 17363 10560 17408 10588
rect 10836 10548 10842 10560
rect 4028 10492 4476 10520
rect 4608 10523 4666 10529
rect 4028 10480 4034 10492
rect 4608 10489 4620 10523
rect 4654 10520 4666 10523
rect 5442 10520 5448 10532
rect 4654 10492 5448 10520
rect 4654 10489 4666 10492
rect 4608 10483 4666 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 14369 10523 14427 10529
rect 14369 10489 14381 10523
rect 14415 10520 14427 10523
rect 15381 10523 15439 10529
rect 14415 10492 15056 10520
rect 14415 10489 14427 10492
rect 14369 10483 14427 10489
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3602 10452 3608 10464
rect 3007 10424 3608 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3602 10412 3608 10424
rect 3660 10452 3666 10464
rect 7190 10452 7196 10464
rect 3660 10424 7196 10452
rect 3660 10412 3666 10424
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7432 10424 7849 10452
rect 7432 10412 7438 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 11609 10455 11667 10461
rect 11609 10421 11621 10455
rect 11655 10452 11667 10455
rect 11698 10452 11704 10464
rect 11655 10424 11704 10452
rect 11655 10421 11667 10424
rect 11609 10415 11667 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 15028 10461 15056 10492
rect 15381 10489 15393 10523
rect 15427 10520 15439 10523
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 15427 10492 16037 10520
rect 15427 10489 15439 10492
rect 15381 10483 15439 10489
rect 16025 10489 16037 10492
rect 16071 10489 16083 10523
rect 16224 10520 16252 10560
rect 17402 10548 17408 10560
rect 17460 10548 17466 10600
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18012 10560 18429 10588
rect 18012 10548 18018 10560
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 18874 10588 18880 10600
rect 18555 10560 18880 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 19978 10520 19984 10532
rect 16224 10492 19984 10520
rect 16025 10483 16083 10489
rect 19978 10480 19984 10492
rect 20036 10480 20042 10532
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13964 10424 14473 10452
rect 13964 10412 13970 10424
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14461 10415 14519 10421
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 17313 10455 17371 10461
rect 17313 10452 17325 10455
rect 16724 10424 17325 10452
rect 16724 10412 16730 10424
rect 17313 10421 17325 10424
rect 17359 10421 17371 10455
rect 17313 10415 17371 10421
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19058 10452 19064 10464
rect 18748 10424 19064 10452
rect 18748 10412 18754 10424
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 19705 10455 19763 10461
rect 19705 10452 19717 10455
rect 19576 10424 19717 10452
rect 19576 10412 19582 10424
rect 19705 10421 19717 10424
rect 19751 10421 19763 10455
rect 20070 10452 20076 10464
rect 20031 10424 20076 10452
rect 19705 10415 19763 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2866 10248 2872 10260
rect 1995 10220 2872 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6362 10248 6368 10260
rect 6319 10220 6368 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10248 6699 10251
rect 7374 10248 7380 10260
rect 6687 10220 7380 10248
rect 6687 10217 6699 10220
rect 6641 10211 6699 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10134 10248 10140 10260
rect 9732 10220 10140 10248
rect 9732 10208 9738 10220
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10284 10220 10701 10248
rect 10284 10208 10290 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 10689 10211 10747 10217
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15746 10248 15752 10260
rect 15335 10220 15752 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 17552 10220 18245 10248
rect 17552 10208 17558 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 19978 10248 19984 10260
rect 19939 10220 19984 10248
rect 18233 10211 18291 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20128 10220 20913 10248
rect 20128 10208 20134 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 15194 10180 15200 10192
rect 4120 10152 15200 10180
rect 4120 10140 4126 10152
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 15378 10140 15384 10192
rect 15436 10180 15442 10192
rect 17954 10180 17960 10192
rect 15436 10152 17960 10180
rect 15436 10140 15442 10152
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 1946 10112 1952 10124
rect 1811 10084 1952 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 6546 10112 6552 10124
rect 4378 10084 6552 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7558 10121 7564 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6696 10084 6745 10112
rect 6696 10072 6702 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 7541 10115 7564 10121
rect 7541 10112 7553 10115
rect 6733 10075 6791 10081
rect 6932 10084 7553 10112
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 4062 10044 4068 10056
rect 3844 10016 4068 10044
rect 3844 10004 3850 10016
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 6656 10044 6684 10072
rect 6932 10053 6960 10084
rect 7541 10081 7553 10084
rect 7541 10075 7564 10081
rect 7558 10072 7564 10075
rect 7616 10072 7622 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9824 10084 10057 10112
rect 9824 10072 9830 10084
rect 10045 10081 10057 10084
rect 10091 10112 10103 10115
rect 10778 10112 10784 10124
rect 10091 10084 10784 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 11698 10121 11704 10124
rect 11692 10112 11704 10121
rect 11659 10084 11704 10112
rect 11692 10075 11704 10084
rect 11698 10072 11704 10075
rect 11756 10072 11762 10124
rect 13170 10072 13176 10124
rect 13228 10112 13234 10124
rect 13337 10115 13395 10121
rect 13337 10112 13349 10115
rect 13228 10084 13349 10112
rect 13228 10072 13234 10084
rect 13337 10081 13349 10084
rect 13383 10081 13395 10115
rect 13337 10075 13395 10081
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 14148 10084 15669 10112
rect 14148 10072 14154 10084
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 17120 10115 17178 10121
rect 17120 10081 17132 10115
rect 17166 10112 17178 10115
rect 17494 10112 17500 10124
rect 17166 10084 17500 10112
rect 17166 10081 17178 10084
rect 17120 10075 17178 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 20073 10115 20131 10121
rect 20073 10081 20085 10115
rect 20119 10112 20131 10115
rect 20254 10112 20260 10124
rect 20119 10084 20260 10112
rect 20119 10081 20131 10084
rect 20073 10075 20131 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 5132 10016 6684 10044
rect 6917 10047 6975 10053
rect 5132 10004 5138 10016
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 7282 10044 7288 10056
rect 7243 10016 7288 10044
rect 6917 10007 6975 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 11425 10047 11483 10053
rect 10284 10016 10329 10044
rect 10284 10004 10290 10016
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 11425 10007 11483 10013
rect 12544 10016 13093 10044
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10778 9976 10784 9988
rect 10192 9948 10784 9976
rect 10192 9936 10198 9948
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6546 9908 6552 9920
rect 6420 9880 6552 9908
rect 6420 9868 6426 9880
rect 6546 9868 6552 9880
rect 6604 9908 6610 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 6604 9880 8677 9908
rect 6604 9868 6610 9880
rect 8665 9877 8677 9880
rect 8711 9877 8723 9911
rect 8665 9871 8723 9877
rect 9677 9911 9735 9917
rect 9677 9877 9689 9911
rect 9723 9908 9735 9911
rect 10962 9908 10968 9920
rect 9723 9880 10968 9908
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 11440 9908 11468 10007
rect 12544 9920 12572 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 13081 10007 13139 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 16850 10044 16856 10056
rect 16811 10016 16856 10044
rect 15841 10007 15899 10013
rect 14461 9979 14519 9985
rect 14461 9945 14473 9979
rect 14507 9976 14519 9979
rect 14550 9976 14556 9988
rect 14507 9948 14556 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 14550 9936 14556 9948
rect 14608 9976 14614 9988
rect 15856 9976 15884 10007
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 20162 10044 20168 10056
rect 20075 10016 20168 10044
rect 20162 10004 20168 10016
rect 20220 10044 20226 10056
rect 20530 10044 20536 10056
rect 20220 10016 20536 10044
rect 20220 10004 20226 10016
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 14608 9948 15884 9976
rect 14608 9936 14614 9948
rect 12526 9908 12532 9920
rect 11440 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12768 9880 12817 9908
rect 12768 9868 12774 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 15194 9908 15200 9920
rect 14056 9880 15200 9908
rect 14056 9868 14062 9880
rect 15194 9868 15200 9880
rect 15252 9868 15258 9920
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 16574 9908 16580 9920
rect 15344 9880 16580 9908
rect 15344 9868 15350 9880
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 19610 9908 19616 9920
rect 19571 9880 19616 9908
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 8294 9704 8300 9716
rect 7708 9676 8300 9704
rect 7708 9664 7714 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9858 9704 9864 9716
rect 8956 9676 9864 9704
rect 5718 9636 5724 9648
rect 5679 9608 5724 9636
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6328 9608 7236 9636
rect 6328 9596 6334 9608
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 6362 9568 6368 9580
rect 6323 9540 6368 9568
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3326 9500 3332 9512
rect 2823 9472 3332 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 7208 9500 7236 9608
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7742 9636 7748 9648
rect 7340 9608 7748 9636
rect 7340 9596 7346 9608
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 8956 9636 8984 9676
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10321 9707 10379 9713
rect 10321 9673 10333 9707
rect 10367 9704 10379 9707
rect 10502 9704 10508 9716
rect 10367 9676 10508 9704
rect 10367 9673 10379 9676
rect 10321 9667 10379 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 12434 9704 12440 9716
rect 10836 9676 12440 9704
rect 10836 9664 10842 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 15657 9707 15715 9713
rect 15657 9673 15669 9707
rect 15703 9704 15715 9707
rect 15746 9704 15752 9716
rect 15703 9676 15752 9704
rect 15703 9673 15715 9676
rect 15657 9667 15715 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16942 9704 16948 9716
rect 16632 9676 16948 9704
rect 16632 9664 16638 9676
rect 16942 9664 16948 9676
rect 17000 9704 17006 9716
rect 19242 9704 19248 9716
rect 17000 9676 19248 9704
rect 17000 9664 17006 9676
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 7800 9608 8984 9636
rect 10520 9636 10548 9664
rect 12529 9639 12587 9645
rect 10520 9608 11192 9636
rect 7800 9596 7806 9608
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8956 9577 8984 9608
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8036 9540 8861 9568
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 4120 9472 7144 9500
rect 7208 9472 7389 9500
rect 4120 9460 4126 9472
rect 3050 9441 3056 9444
rect 3044 9432 3056 9441
rect 3011 9404 3056 9432
rect 3044 9395 3056 9404
rect 3050 9392 3056 9395
rect 3108 9392 3114 9444
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9432 6147 9435
rect 7116 9432 7144 9472
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8036 9500 8064 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11164 9577 11192 9608
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 13906 9636 13912 9648
rect 12575 9608 13912 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 15838 9636 15844 9648
rect 15427 9608 15844 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 11020 9540 11069 9568
rect 11020 9528 11026 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 13170 9568 13176 9580
rect 13131 9540 13176 9568
rect 11149 9531 11207 9537
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 14008 9571 14066 9577
rect 14008 9568 14020 9571
rect 13412 9540 14020 9568
rect 13412 9528 13418 9540
rect 14008 9537 14020 9540
rect 14054 9537 14066 9571
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 14008 9531 14066 9537
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 8202 9500 8208 9512
rect 7515 9472 8064 9500
rect 8163 9472 8208 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 9208 9503 9266 9509
rect 8312 9472 8892 9500
rect 8312 9432 8340 9472
rect 6135 9404 7052 9432
rect 7116 9404 8340 9432
rect 8864 9432 8892 9472
rect 9208 9469 9220 9503
rect 9254 9500 9266 9503
rect 9674 9500 9680 9512
rect 9254 9472 9680 9500
rect 9254 9469 9266 9472
rect 9208 9463 9266 9469
rect 9674 9460 9680 9472
rect 9732 9500 9738 9512
rect 10226 9500 10232 9512
rect 9732 9472 10232 9500
rect 9732 9460 9738 9472
rect 10226 9460 10232 9472
rect 10284 9460 10290 9512
rect 12986 9500 12992 9512
rect 12947 9472 12992 9500
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13872 9472 13921 9500
rect 13872 9460 13878 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14268 9503 14326 9509
rect 14268 9469 14280 9503
rect 14314 9500 14326 9503
rect 14550 9500 14556 9512
rect 14314 9472 14556 9500
rect 14314 9469 14326 9472
rect 14268 9463 14326 9469
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14660 9472 17816 9500
rect 12250 9432 12256 9444
rect 8864 9404 12256 9432
rect 6135 9401 6147 9404
rect 6089 9395 6147 9401
rect 4154 9364 4160 9376
rect 4115 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 7024 9373 7052 9404
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12360 9404 12909 9432
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8202 9364 8208 9376
rect 8067 9336 8208 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9858 9364 9864 9376
rect 8895 9336 9864 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10928 9336 10977 9364
rect 10928 9324 10934 9336
rect 10965 9333 10977 9336
rect 11011 9364 11023 9367
rect 11606 9364 11612 9376
rect 11011 9336 11612 9364
rect 11011 9333 11023 9336
rect 10965 9327 11023 9333
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12360 9364 12388 9404
rect 12897 9401 12909 9404
rect 12943 9432 12955 9435
rect 13998 9432 14004 9444
rect 12943 9404 14004 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 13998 9392 14004 9404
rect 14056 9432 14062 9444
rect 14660 9432 14688 9472
rect 14056 9404 14688 9432
rect 16025 9435 16083 9441
rect 14056 9392 14062 9404
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 17678 9432 17684 9444
rect 16071 9404 17684 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 17678 9392 17684 9404
rect 17736 9392 17742 9444
rect 17788 9432 17816 9472
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19392 9472 19625 9500
rect 19392 9460 19398 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19880 9503 19938 9509
rect 19880 9469 19892 9503
rect 19926 9500 19938 9503
rect 20162 9500 20168 9512
rect 19926 9472 20168 9500
rect 19926 9469 19938 9472
rect 19880 9463 19938 9469
rect 20162 9460 20168 9472
rect 20220 9460 20226 9512
rect 19794 9432 19800 9444
rect 17788 9404 19800 9432
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 11940 9336 12388 9364
rect 11940 9324 11946 9336
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 13354 9364 13360 9376
rect 12584 9336 13360 9364
rect 12584 9324 12590 9336
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13722 9364 13728 9376
rect 13683 9336 13728 9364
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 16117 9367 16175 9373
rect 16117 9333 16129 9367
rect 16163 9364 16175 9367
rect 16574 9364 16580 9376
rect 16163 9336 16580 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16574 9324 16580 9336
rect 16632 9364 16638 9376
rect 17218 9364 17224 9376
rect 16632 9336 17224 9364
rect 16632 9324 16638 9336
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 19058 9364 19064 9376
rect 18840 9336 19064 9364
rect 18840 9324 18846 9336
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 20990 9364 20996 9376
rect 20951 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5166 9160 5172 9172
rect 4571 9132 5172 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 7193 9163 7251 9169
rect 7193 9160 7205 9163
rect 6236 9132 7205 9160
rect 6236 9120 6242 9132
rect 7193 9129 7205 9132
rect 7239 9129 7251 9163
rect 7193 9123 7251 9129
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 7432 9132 8677 9160
rect 7432 9120 7438 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 10652 9132 11253 9160
rect 10652 9120 10658 9132
rect 11241 9129 11253 9132
rect 11287 9129 11299 9163
rect 11241 9123 11299 9129
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12860 9132 13093 9160
rect 12860 9120 12866 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 17552 9132 18245 9160
rect 17552 9120 17558 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 18874 9120 18880 9172
rect 18932 9160 18938 9172
rect 19150 9160 19156 9172
rect 18932 9132 19156 9160
rect 18932 9120 18938 9132
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19610 9160 19616 9172
rect 19571 9132 19616 9160
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 3326 9092 3332 9104
rect 1688 9064 3332 9092
rect 1688 9033 1716 9064
rect 3326 9052 3332 9064
rect 3384 9092 3390 9104
rect 3970 9092 3976 9104
rect 3384 9064 3976 9092
rect 3384 9052 3390 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 5534 9092 5540 9104
rect 4120 9064 5540 9092
rect 4120 9052 4126 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 6788 9064 8585 9092
rect 6788 9052 6794 9064
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8573 9055 8631 9061
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 18506 9092 18512 9104
rect 11664 9064 18512 9092
rect 11664 9052 11670 9064
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 19518 9092 19524 9104
rect 19479 9064 19524 9092
rect 19518 9052 19524 9064
rect 19576 9052 19582 9104
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 1940 9027 1998 9033
rect 1940 8993 1952 9027
rect 1986 9024 1998 9027
rect 2958 9024 2964 9036
rect 1986 8996 2964 9024
rect 1986 8993 1998 8996
rect 1940 8987 1998 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4433 8987 4491 8993
rect 3050 8820 3056 8832
rect 3011 8792 3056 8820
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4246 8820 4252 8832
rect 4111 8792 4252 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4448 8820 4476 8987
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 5793 9027 5851 9033
rect 5793 9024 5805 9027
rect 5684 8996 5805 9024
rect 5684 8984 5690 8996
rect 5793 8993 5805 8996
rect 5839 8993 5851 9027
rect 5793 8987 5851 8993
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 6880 8996 7573 9024
rect 6880 8984 6886 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 11146 9024 11152 9036
rect 11107 8996 11152 9024
rect 7561 8987 7619 8993
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 12986 9024 12992 9036
rect 11348 8996 12848 9024
rect 12947 8996 12992 9024
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5500 8928 5549 8956
rect 5500 8916 5506 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7156 8928 7665 8956
rect 7156 8916 7162 8928
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8849 8959 8907 8965
rect 8849 8925 8861 8959
rect 8895 8956 8907 8959
rect 11348 8956 11376 8996
rect 8895 8928 11376 8956
rect 11425 8959 11483 8965
rect 8895 8925 8907 8928
rect 8849 8919 8907 8925
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 11698 8956 11704 8968
rect 11471 8928 11704 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 6917 8891 6975 8897
rect 6917 8857 6929 8891
rect 6963 8888 6975 8891
rect 7558 8888 7564 8900
rect 6963 8860 7564 8888
rect 6963 8857 6975 8860
rect 6917 8851 6975 8857
rect 7558 8848 7564 8860
rect 7616 8888 7622 8900
rect 7760 8888 7788 8919
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12820 8956 12848 8996
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 17120 9027 17178 9033
rect 17120 8993 17132 9027
rect 17166 9024 17178 9027
rect 17586 9024 17592 9036
rect 17166 8996 17592 9024
rect 17166 8993 17178 8996
rect 17120 8987 17178 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 13170 8956 13176 8968
rect 12820 8928 13176 8956
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8956 13323 8959
rect 13814 8956 13820 8968
rect 13311 8928 13820 8956
rect 13311 8925 13323 8928
rect 13265 8919 13323 8925
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 19794 8956 19800 8968
rect 19707 8928 19800 8956
rect 19794 8916 19800 8928
rect 19852 8956 19858 8968
rect 20990 8956 20996 8968
rect 19852 8928 20996 8956
rect 19852 8916 19858 8928
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 7616 8860 7788 8888
rect 8205 8891 8263 8897
rect 7616 8848 7622 8860
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 14090 8888 14096 8900
rect 8251 8860 14096 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 14090 8848 14096 8860
rect 14148 8848 14154 8900
rect 5718 8820 5724 8832
rect 4448 8792 5724 8820
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7190 8820 7196 8832
rect 6696 8792 7196 8820
rect 6696 8780 6702 8792
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 10781 8823 10839 8829
rect 10781 8789 10793 8823
rect 10827 8820 10839 8823
rect 11698 8820 11704 8832
rect 10827 8792 11704 8820
rect 10827 8789 10839 8792
rect 10781 8783 10839 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12618 8820 12624 8832
rect 12579 8792 12624 8820
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19153 8823 19211 8829
rect 19153 8820 19165 8823
rect 18840 8792 19165 8820
rect 18840 8780 18846 8792
rect 19153 8789 19165 8792
rect 19199 8789 19211 8823
rect 19153 8783 19211 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 5626 8616 5632 8628
rect 5587 8588 5632 8616
rect 5626 8576 5632 8588
rect 5684 8616 5690 8628
rect 6822 8616 6828 8628
rect 5684 8588 6500 8616
rect 6783 8588 6828 8616
rect 5684 8576 5690 8588
rect 2958 8480 2964 8492
rect 2919 8452 2964 8480
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 6472 8480 6500 8588
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9674 8616 9680 8628
rect 9539 8588 9680 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10226 8508 10232 8560
rect 10284 8548 10290 8560
rect 10778 8548 10784 8560
rect 10284 8520 10784 8548
rect 10284 8508 10290 8520
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 13814 8548 13820 8560
rect 13775 8520 13820 8548
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 17218 8548 17224 8560
rect 16991 8520 17224 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 17328 8520 18061 8548
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6472 8452 7389 8480
rect 7377 8449 7389 8452
rect 7423 8480 7435 8483
rect 7558 8480 7564 8492
rect 7423 8452 7564 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 7800 8452 8125 8480
rect 7800 8440 7806 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3142 8412 3148 8424
rect 2832 8384 3148 8412
rect 2832 8372 2838 8384
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 4028 8384 4261 8412
rect 4028 8372 4034 8384
rect 4249 8381 4261 8384
rect 4295 8412 4307 8415
rect 5442 8412 5448 8424
rect 4295 8384 5448 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 5442 8372 5448 8384
rect 5500 8412 5506 8424
rect 5626 8412 5632 8424
rect 5500 8384 5632 8412
rect 5500 8372 5506 8384
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 7116 8384 7205 8412
rect 2685 8347 2743 8353
rect 2685 8313 2697 8347
rect 2731 8344 2743 8347
rect 3234 8344 3240 8356
rect 2731 8316 3240 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 4494 8347 4552 8353
rect 4494 8313 4506 8347
rect 4540 8313 4552 8347
rect 4494 8307 4552 8313
rect 2314 8276 2320 8288
rect 2275 8248 2320 8276
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 4154 8276 4160 8288
rect 2648 8248 4160 8276
rect 2648 8236 2654 8248
rect 4154 8236 4160 8248
rect 4212 8276 4218 8288
rect 4509 8276 4537 8307
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7116 8344 7144 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7340 8384 7385 8412
rect 7340 8372 7346 8384
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 10962 8412 10968 8424
rect 7984 8384 10968 8412
rect 7984 8372 7990 8384
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12400 8384 12449 8412
rect 12400 8372 12406 8384
rect 12437 8381 12449 8384
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12710 8421 12716 8424
rect 12704 8412 12716 8421
rect 12671 8384 12716 8412
rect 12704 8375 12716 8384
rect 12710 8372 12716 8375
rect 12768 8372 12774 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 15841 8415 15899 8421
rect 15841 8412 15853 8415
rect 13780 8384 15853 8412
rect 13780 8372 13786 8384
rect 15841 8381 15853 8384
rect 15887 8381 15899 8415
rect 16666 8412 16672 8424
rect 15841 8375 15899 8381
rect 15939 8384 16672 8412
rect 6880 8316 7144 8344
rect 8380 8347 8438 8353
rect 6880 8304 6886 8316
rect 8380 8313 8392 8347
rect 8426 8344 8438 8347
rect 8478 8344 8484 8356
rect 8426 8316 8484 8344
rect 8426 8313 8438 8316
rect 8380 8307 8438 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 11882 8344 11888 8356
rect 10704 8316 11888 8344
rect 4212 8248 4537 8276
rect 4212 8236 4218 8248
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 10704 8276 10732 8316
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 15939 8344 15967 8384
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 17328 8421 17356 8520
rect 18049 8517 18061 8520
rect 18095 8517 18107 8551
rect 18049 8511 18107 8517
rect 17494 8480 17500 8492
rect 17455 8452 17500 8480
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 17644 8452 18613 8480
rect 17644 8440 17650 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18966 8440 18972 8492
rect 19024 8440 19030 8492
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18984 8412 19012 8440
rect 18555 8384 19012 8412
rect 19245 8415 19303 8421
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 19334 8412 19340 8424
rect 19291 8384 19340 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19512 8415 19570 8421
rect 19512 8381 19524 8415
rect 19558 8412 19570 8415
rect 19794 8412 19800 8424
rect 19558 8384 19800 8412
rect 19558 8381 19570 8384
rect 19512 8375 19570 8381
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 12452 8316 15967 8344
rect 4764 8248 10732 8276
rect 4764 8236 4770 8248
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 12452 8276 12480 8316
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 18966 8344 18972 8356
rect 16632 8316 18972 8344
rect 16632 8304 16638 8316
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 10836 8248 12480 8276
rect 10836 8236 10842 8248
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13170 8276 13176 8288
rect 12952 8248 13176 8276
rect 12952 8236 12958 8248
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 15657 8279 15715 8285
rect 15657 8245 15669 8279
rect 15703 8276 15715 8279
rect 16206 8276 16212 8288
rect 15703 8248 16212 8276
rect 15703 8245 15715 8248
rect 15657 8239 15715 8245
rect 16206 8236 16212 8248
rect 16264 8276 16270 8288
rect 16850 8276 16856 8288
rect 16264 8248 16856 8276
rect 16264 8236 16270 8248
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 20622 8276 20628 8288
rect 20583 8248 20628 8276
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1762 8072 1768 8084
rect 1443 8044 1768 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 1857 8075 1915 8081
rect 1857 8041 1869 8075
rect 1903 8072 1915 8075
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 1903 8044 4077 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4304 8044 4445 8072
rect 4304 8032 4310 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 6641 8075 6699 8081
rect 6641 8041 6653 8075
rect 6687 8072 6699 8075
rect 7098 8072 7104 8084
rect 6687 8044 7104 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7742 8072 7748 8084
rect 7340 8044 7748 8072
rect 7340 8032 7346 8044
rect 7742 8032 7748 8044
rect 7800 8072 7806 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7800 8044 8125 8072
rect 7800 8032 7806 8044
rect 8113 8041 8125 8044
rect 8159 8072 8171 8075
rect 9674 8072 9680 8084
rect 8159 8044 9680 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 12342 8072 12348 8084
rect 12303 8044 12348 8072
rect 10137 8035 10195 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12621 8075 12679 8081
rect 12621 8041 12633 8075
rect 12667 8072 12679 8075
rect 17037 8075 17095 8081
rect 12667 8044 14136 8072
rect 12667 8041 12679 8044
rect 12621 8035 12679 8041
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 2777 8007 2835 8013
rect 2777 8004 2789 8007
rect 2740 7976 2789 8004
rect 2740 7964 2746 7976
rect 2777 7973 2789 7976
rect 2823 8004 2835 8007
rect 3142 8004 3148 8016
rect 2823 7976 3148 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 8202 8004 8208 8016
rect 5828 7976 8208 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2222 7936 2228 7948
rect 1811 7908 2228 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 3050 7896 3056 7948
rect 3108 7936 3114 7948
rect 5828 7945 5856 7976
rect 8202 7964 8208 7976
rect 8260 8004 8266 8016
rect 8260 7976 8340 8004
rect 8260 7964 8266 7976
rect 5813 7939 5871 7945
rect 3108 7908 4660 7936
rect 3108 7896 3114 7908
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2590 7868 2596 7880
rect 2087 7840 2596 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 4632 7877 4660 7908
rect 5813 7905 5825 7939
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 8312 7945 8340 7976
rect 8570 7964 8576 8016
rect 8628 8004 8634 8016
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 8628 7976 13001 8004
rect 8628 7964 8634 7976
rect 12989 7973 13001 7976
rect 13035 8004 13047 8007
rect 13262 8004 13268 8016
rect 13035 7976 13268 8004
rect 13035 7973 13047 7976
rect 12989 7967 13047 7973
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 13998 8004 14004 8016
rect 13959 7976 14004 8004
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 14108 8013 14136 8044
rect 17037 8041 17049 8075
rect 17083 8072 17095 8075
rect 17402 8072 17408 8084
rect 17083 8044 17408 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17678 8072 17684 8084
rect 17543 8044 17684 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 18414 8072 18420 8084
rect 18095 8044 18420 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 20346 8072 20352 8084
rect 20211 8044 20352 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 14093 8007 14151 8013
rect 14093 7973 14105 8007
rect 14139 7973 14151 8007
rect 14093 7967 14151 7973
rect 15556 8007 15614 8013
rect 15556 7973 15568 8007
rect 15602 8004 15614 8007
rect 15838 8004 15844 8016
rect 15602 7976 15844 8004
rect 15602 7973 15614 7976
rect 15556 7967 15614 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 15930 7964 15936 8016
rect 15988 8004 15994 8016
rect 20073 8007 20131 8013
rect 20073 8004 20085 8007
rect 15988 7976 20085 8004
rect 15988 7964 15994 7976
rect 20073 7973 20085 7976
rect 20119 7973 20131 8007
rect 20073 7967 20131 7973
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6052 7908 6561 7936
rect 6052 7896 6058 7908
rect 6549 7905 6561 7908
rect 6595 7936 6607 7939
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6595 7908 7021 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 7009 7905 7021 7908
rect 7055 7936 7067 7939
rect 8297 7939 8355 7945
rect 7055 7908 7972 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 4525 7871 4583 7877
rect 3016 7840 3061 7868
rect 3016 7828 3022 7840
rect 4525 7837 4537 7871
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4540 7800 4568 7831
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6788 7840 7113 7868
rect 6788 7828 6794 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7868 7343 7871
rect 7558 7868 7564 7880
rect 7331 7840 7564 7868
rect 7331 7837 7343 7840
rect 7285 7831 7343 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7944 7868 7972 7908
rect 8297 7905 8309 7939
rect 8343 7905 8355 7939
rect 8297 7899 8355 7905
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 8444 7908 10057 7936
rect 8444 7896 8450 7908
rect 10045 7905 10057 7908
rect 10091 7936 10103 7939
rect 12529 7939 12587 7945
rect 10091 7908 10640 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10612 7877 10640 7908
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 13722 7936 13728 7948
rect 12575 7908 13728 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 17402 7936 17408 7948
rect 13832 7908 16344 7936
rect 17363 7908 17408 7936
rect 10229 7871 10287 7877
rect 7944 7840 9996 7868
rect 8662 7800 8668 7812
rect 4540 7772 8668 7800
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 9766 7800 9772 7812
rect 8772 7772 9772 7800
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 2682 7732 2688 7744
rect 2455 7704 2688 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 5626 7732 5632 7744
rect 5587 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 8772 7732 8800 7772
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 6236 7704 8800 7732
rect 6236 7692 6242 7704
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9180 7704 9689 7732
rect 9180 7692 9186 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9968 7732 9996 7840
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 13081 7871 13139 7877
rect 10643 7840 12572 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10042 7760 10048 7812
rect 10100 7800 10106 7812
rect 10244 7800 10272 7831
rect 10100 7772 10272 7800
rect 10100 7760 10106 7772
rect 11974 7732 11980 7744
rect 9968 7704 11980 7732
rect 9677 7695 9735 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 12544 7732 12572 7840
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13170 7868 13176 7880
rect 13127 7840 13176 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13832 7868 13860 7908
rect 13265 7831 13323 7837
rect 13372 7840 13860 7868
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 13280 7800 13308 7831
rect 13372 7812 13400 7840
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13964 7840 14197 7868
rect 13964 7828 13970 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 14185 7831 14243 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 16316 7868 16344 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 18046 7936 18052 7948
rect 17512 7908 18052 7936
rect 17512 7868 17540 7908
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 16316 7840 17540 7868
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 20349 7871 20407 7877
rect 17644 7840 17689 7868
rect 17644 7828 17650 7840
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20622 7868 20628 7880
rect 20395 7840 20628 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 12768 7772 13308 7800
rect 12768 7760 12774 7772
rect 13354 7760 13360 7812
rect 13412 7760 13418 7812
rect 13464 7772 13768 7800
rect 13464 7732 13492 7772
rect 13630 7732 13636 7744
rect 12544 7704 13492 7732
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13740 7732 13768 7772
rect 14274 7732 14280 7744
rect 13740 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 17126 7732 17132 7744
rect 16715 7704 17132 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 19668 7704 19717 7732
rect 19668 7692 19674 7704
rect 19705 7701 19717 7704
rect 19751 7701 19763 7735
rect 19705 7695 19763 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 10870 7528 10876 7540
rect 8812 7500 10876 7528
rect 8812 7488 8818 7500
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12250 7528 12256 7540
rect 11112 7500 12256 7528
rect 11112 7488 11118 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 17586 7528 17592 7540
rect 12492 7500 17172 7528
rect 17547 7500 17592 7528
rect 12492 7488 12498 7500
rect 5721 7463 5779 7469
rect 5721 7429 5733 7463
rect 5767 7460 5779 7463
rect 8202 7460 8208 7472
rect 5767 7432 8208 7460
rect 5767 7429 5779 7432
rect 5721 7423 5779 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 17144 7460 17172 7500
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 18506 7460 18512 7472
rect 17144 7432 18512 7460
rect 18506 7420 18512 7432
rect 18564 7420 18570 7472
rect 2682 7392 2688 7404
rect 2643 7364 2688 7392
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3050 7392 3056 7404
rect 2915 7364 3056 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 7190 7392 7196 7404
rect 6411 7364 7196 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 9306 7392 9312 7404
rect 9219 7364 9312 7392
rect 9306 7352 9312 7364
rect 9364 7392 9370 7404
rect 12805 7395 12863 7401
rect 9364 7364 9812 7392
rect 9364 7352 9370 7364
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 2593 7327 2651 7333
rect 2593 7324 2605 7327
rect 2372 7296 2605 7324
rect 2372 7284 2378 7296
rect 2593 7293 2605 7296
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9674 7324 9680 7336
rect 9180 7296 9225 7324
rect 9635 7296 9680 7324
rect 9180 7284 9186 7296
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 9784 7324 9812 7364
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 12986 7392 12992 7404
rect 12851 7364 12992 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 9784 7296 11100 7324
rect 5994 7216 6000 7268
rect 6052 7256 6058 7268
rect 6089 7259 6147 7265
rect 6089 7256 6101 7259
rect 6052 7228 6101 7256
rect 6052 7216 6058 7228
rect 6089 7225 6101 7228
rect 6135 7225 6147 7259
rect 6089 7219 6147 7225
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 9944 7259 10002 7265
rect 6420 7228 9168 7256
rect 6420 7216 6426 7228
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5868 7160 6193 7188
rect 5868 7148 5874 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 9030 7188 9036 7200
rect 8991 7160 9036 7188
rect 6181 7151 6239 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9140 7188 9168 7228
rect 9944 7225 9956 7259
rect 9990 7256 10002 7259
rect 10042 7256 10048 7268
rect 9990 7228 10048 7256
rect 9990 7225 10002 7228
rect 9944 7219 10002 7225
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 9766 7188 9772 7200
rect 9140 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 10870 7188 10876 7200
rect 10652 7160 10876 7188
rect 10652 7148 10658 7160
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 11072 7197 11100 7296
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 13265 7327 13323 7333
rect 13265 7324 13277 7327
rect 12400 7296 13277 7324
rect 12400 7284 12406 7296
rect 13265 7293 13277 7296
rect 13311 7293 13323 7327
rect 13265 7287 13323 7293
rect 13532 7327 13590 7333
rect 13532 7293 13544 7327
rect 13578 7324 13590 7327
rect 13814 7324 13820 7336
rect 13578 7296 13820 7324
rect 13578 7293 13590 7296
rect 13532 7287 13590 7293
rect 13280 7256 13308 7287
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 13964 7296 16160 7324
rect 13964 7284 13970 7296
rect 13446 7256 13452 7268
rect 13280 7228 13452 7256
rect 13446 7216 13452 7228
rect 13504 7256 13510 7268
rect 15286 7256 15292 7268
rect 13504 7228 15292 7256
rect 13504 7216 13510 7228
rect 15286 7216 15292 7228
rect 15344 7216 15350 7268
rect 16132 7256 16160 7296
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 16482 7333 16488 7336
rect 16264 7296 16309 7324
rect 16264 7284 16270 7296
rect 16476 7287 16488 7333
rect 16540 7324 16546 7336
rect 19334 7324 19340 7336
rect 16540 7296 16576 7324
rect 19295 7296 19340 7324
rect 16482 7284 16488 7287
rect 16540 7284 16546 7296
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 19426 7284 19432 7336
rect 19484 7284 19490 7336
rect 19604 7327 19662 7333
rect 19604 7293 19616 7327
rect 19650 7324 19662 7327
rect 20622 7324 20628 7336
rect 19650 7296 20628 7324
rect 19650 7293 19662 7296
rect 19604 7287 19662 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 19444 7256 19472 7284
rect 20530 7256 20536 7268
rect 16132 7228 20536 7256
rect 20530 7216 20536 7228
rect 20588 7216 20594 7268
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 12710 7188 12716 7200
rect 11204 7160 12716 7188
rect 11204 7148 11210 7160
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 13780 7160 14657 7188
rect 13780 7148 13786 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 14645 7151 14703 7157
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 17954 7188 17960 7200
rect 15528 7160 17960 7188
rect 15528 7148 15534 7160
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 19426 7148 19432 7200
rect 19484 7188 19490 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 19484 7160 20729 7188
rect 19484 7148 19490 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 5810 6984 5816 6996
rect 5771 6956 5816 6984
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 6178 6984 6184 6996
rect 6139 6956 6184 6984
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 6696 6956 8217 6984
rect 6696 6944 6702 6956
rect 8205 6953 8217 6956
rect 8251 6984 8263 6987
rect 8570 6984 8576 6996
rect 8251 6956 8576 6984
rect 8251 6953 8263 6956
rect 8205 6947 8263 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 11606 6984 11612 6996
rect 10520 6956 11612 6984
rect 1302 6876 1308 6928
rect 1360 6916 1366 6928
rect 2501 6919 2559 6925
rect 2501 6916 2513 6919
rect 1360 6888 2513 6916
rect 1360 6876 1366 6888
rect 2501 6885 2513 6888
rect 2547 6916 2559 6919
rect 2961 6919 3019 6925
rect 2961 6916 2973 6919
rect 2547 6888 2973 6916
rect 2547 6885 2559 6888
rect 2501 6879 2559 6885
rect 2961 6885 2973 6888
rect 3007 6916 3019 6919
rect 6362 6916 6368 6928
rect 3007 6888 6368 6916
rect 3007 6885 3019 6888
rect 2961 6879 3019 6885
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 6914 6876 6920 6928
rect 6972 6916 6978 6928
rect 8386 6916 8392 6928
rect 6972 6888 8392 6916
rect 6972 6876 6978 6888
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 6178 6848 6184 6860
rect 4120 6820 6184 6848
rect 4120 6808 4126 6820
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6848 6331 6851
rect 7926 6848 7932 6860
rect 6319 6820 7932 6848
rect 6319 6817 6331 6820
rect 6273 6811 6331 6817
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 1946 6780 1952 6792
rect 1903 6752 1952 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 2222 6672 2228 6724
rect 2280 6712 2286 6724
rect 3160 6712 3188 6743
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 6288 6780 6316 6811
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 10520 6848 10548 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12676 6956 12909 6984
rect 12676 6944 12682 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13630 6984 13636 6996
rect 13035 6956 13636 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 12342 6916 12348 6928
rect 10612 6888 12348 6916
rect 10612 6857 10640 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 16206 6916 16212 6928
rect 15304 6888 16212 6916
rect 15304 6857 15332 6888
rect 16206 6876 16212 6888
rect 16264 6916 16270 6928
rect 16758 6916 16764 6928
rect 16264 6888 16764 6916
rect 16264 6876 16270 6888
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 19334 6916 19340 6928
rect 19260 6888 19340 6916
rect 8312 6820 10548 6848
rect 10597 6851 10655 6857
rect 5960 6752 6316 6780
rect 6457 6783 6515 6789
rect 5960 6740 5966 6752
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 2280 6684 3188 6712
rect 6472 6712 6500 6743
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 8312 6789 8340 6820
rect 10597 6817 10609 6851
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10864 6851 10922 6857
rect 10864 6817 10876 6851
rect 10910 6848 10922 6851
rect 15289 6851 15347 6857
rect 10910 6820 13216 6848
rect 10910 6817 10922 6820
rect 10864 6811 10922 6817
rect 13188 6789 13216 6820
rect 15289 6817 15301 6851
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15556 6851 15614 6857
rect 15556 6817 15568 6851
rect 15602 6848 15614 6851
rect 16574 6848 16580 6860
rect 15602 6820 16580 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16776 6848 16804 6876
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 16776 6820 19165 6848
rect 19153 6817 19165 6820
rect 19199 6848 19211 6851
rect 19260 6848 19288 6888
rect 19334 6876 19340 6888
rect 19392 6876 19398 6928
rect 19426 6857 19432 6860
rect 19420 6848 19432 6857
rect 19199 6820 19288 6848
rect 19387 6820 19432 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 19420 6811 19432 6820
rect 19426 6808 19432 6811
rect 19484 6808 19490 6860
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7524 6752 8309 6780
rect 7524 6740 7530 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13722 6780 13728 6792
rect 13219 6752 13728 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 6914 6712 6920 6724
rect 6472 6684 6920 6712
rect 2280 6672 2286 6684
rect 6914 6672 6920 6684
rect 6972 6712 6978 6724
rect 7558 6712 7564 6724
rect 6972 6684 7564 6712
rect 6972 6672 6978 6684
rect 7558 6672 7564 6684
rect 7616 6712 7622 6724
rect 8404 6712 8432 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 17000 6752 17049 6780
rect 17000 6740 17006 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 18690 6780 18696 6792
rect 18651 6752 18696 6780
rect 17037 6743 17095 6749
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 7616 6684 8432 6712
rect 7616 6672 7622 6684
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 13906 6712 13912 6724
rect 12492 6684 13912 6712
rect 12492 6672 12498 6684
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 16224 6684 16804 6712
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 1912 6616 2605 6644
rect 1912 6604 1918 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7800 6616 7849 6644
rect 7800 6604 7806 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 10778 6644 10784 6656
rect 7984 6616 10784 6644
rect 7984 6604 7990 6616
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11977 6647 12035 6653
rect 11977 6644 11989 6647
rect 11020 6616 11989 6644
rect 11020 6604 11026 6616
rect 11977 6613 11989 6616
rect 12023 6613 12035 6647
rect 11977 6607 12035 6613
rect 12529 6647 12587 6653
rect 12529 6613 12541 6647
rect 12575 6644 12587 6647
rect 13078 6644 13084 6656
rect 12575 6616 13084 6644
rect 12575 6613 12587 6616
rect 12529 6607 12587 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 16224 6644 16252 6684
rect 13320 6616 16252 6644
rect 13320 6604 13326 6616
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16540 6616 16681 6644
rect 16540 6604 16546 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16776 6644 16804 6684
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 16776 6616 20545 6644
rect 16669 6607 16727 6613
rect 20533 6613 20545 6616
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5994 6440 6000 6452
rect 5307 6412 6000 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 7282 6440 7288 6452
rect 7116 6412 7288 6440
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2222 6304 2228 6316
rect 2183 6276 2228 6304
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5592 6276 5733 6304
rect 5592 6264 5598 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 5994 6304 6000 6316
rect 5951 6276 6000 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 5994 6264 6000 6276
rect 6052 6304 6058 6316
rect 6914 6304 6920 6316
rect 6052 6276 6920 6304
rect 6052 6264 6058 6276
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7116 6313 7144 6412
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8478 6440 8484 6452
rect 7524 6412 8064 6440
rect 8439 6412 8484 6440
rect 7524 6400 7530 6412
rect 8036 6372 8064 6412
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9088 6412 9413 6440
rect 9088 6400 9094 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 12434 6440 12440 6452
rect 10459 6412 12440 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 18506 6440 18512 6452
rect 12584 6412 18512 6440
rect 12584 6400 12590 6412
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 11882 6372 11888 6384
rect 8036 6344 11888 6372
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 17954 6372 17960 6384
rect 11992 6344 17960 6372
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 10042 6304 10048 6316
rect 9955 6276 10048 6304
rect 7101 6267 7159 6273
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 11330 6304 11336 6316
rect 11103 6276 11336 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11992 6304 12020 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 19426 6332 19432 6384
rect 19484 6372 19490 6384
rect 19484 6344 19748 6372
rect 19484 6332 19490 6344
rect 11664 6276 12020 6304
rect 11664 6264 11670 6276
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13541 6307 13599 6313
rect 13228 6276 13492 6304
rect 13228 6264 13234 6276
rect 1946 6236 1952 6248
rect 1907 6208 1952 6236
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 3786 6236 3792 6248
rect 2731 6208 3792 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7357 6239 7415 6245
rect 7357 6236 7369 6239
rect 7248 6208 7369 6236
rect 7248 6196 7254 6208
rect 7357 6205 7369 6208
rect 7403 6205 7415 6239
rect 7357 6199 7415 6205
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 9214 6236 9220 6248
rect 8720 6208 9220 6236
rect 8720 6196 8726 6208
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9858 6236 9864 6248
rect 9692 6208 9864 6236
rect 2498 6128 2504 6180
rect 2556 6168 2562 6180
rect 2930 6171 2988 6177
rect 2930 6168 2942 6171
rect 2556 6140 2942 6168
rect 2556 6128 2562 6140
rect 2930 6137 2942 6140
rect 2976 6137 2988 6171
rect 2930 6131 2988 6137
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 6273 6171 6331 6177
rect 6273 6168 6285 6171
rect 5675 6140 6285 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 6273 6137 6285 6140
rect 6319 6137 6331 6171
rect 6273 6131 6331 6137
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 9692 6168 9720 6208
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 10060 6236 10088 6264
rect 13262 6236 13268 6248
rect 10060 6208 13268 6236
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13464 6245 13492 6276
rect 13541 6273 13553 6307
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 13449 6239 13507 6245
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 13556 6180 13584 6267
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15436 6276 15577 6304
rect 15436 6264 15442 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 16574 6304 16580 6316
rect 15795 6276 16580 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 16574 6264 16580 6276
rect 16632 6304 16638 6316
rect 17221 6307 17279 6313
rect 17221 6304 17233 6307
rect 16632 6276 17233 6304
rect 16632 6264 16638 6276
rect 17221 6273 17233 6276
rect 17267 6304 17279 6307
rect 17310 6304 17316 6316
rect 17267 6276 17316 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 17920 6276 18613 6304
rect 17920 6264 17926 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 19610 6304 19616 6316
rect 19571 6276 19616 6304
rect 18601 6267 18659 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 19720 6313 19748 6344
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20717 6307 20775 6313
rect 20717 6304 20729 6307
rect 19852 6276 20729 6304
rect 19852 6264 19858 6276
rect 20717 6273 20729 6276
rect 20763 6273 20775 6307
rect 20717 6267 20775 6273
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 17092 6208 17137 6236
rect 17092 6196 17098 6208
rect 18690 6196 18696 6248
rect 18748 6236 18754 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 18748 6208 19533 6236
rect 18748 6196 18754 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 20530 6196 20536 6248
rect 20588 6236 20594 6248
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 20588 6208 20637 6236
rect 20588 6196 20594 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 6788 6140 9720 6168
rect 13357 6171 13415 6177
rect 6788 6128 6794 6140
rect 13357 6137 13369 6171
rect 13403 6168 13415 6171
rect 13403 6140 13492 6168
rect 13403 6137 13415 6140
rect 13357 6131 13415 6137
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 5258 6100 5264 6112
rect 4212 6072 5264 6100
rect 4212 6060 4218 6072
rect 5258 6060 5264 6072
rect 5316 6100 5322 6112
rect 9122 6100 9128 6112
rect 5316 6072 9128 6100
rect 5316 6060 5322 6072
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9272 6072 9781 6100
rect 9272 6060 9278 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 9769 6063 9827 6069
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10778 6100 10784 6112
rect 9916 6072 9961 6100
rect 10739 6072 10784 6100
rect 9916 6060 9922 6072
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 12989 6103 13047 6109
rect 10928 6072 10973 6100
rect 10928 6060 10934 6072
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 13262 6100 13268 6112
rect 13035 6072 13268 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13262 6060 13268 6072
rect 13320 6060 13326 6112
rect 13464 6100 13492 6140
rect 13538 6128 13544 6180
rect 13596 6128 13602 6180
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 13780 6140 15485 6168
rect 13780 6128 13786 6140
rect 15473 6137 15485 6140
rect 15519 6137 15531 6171
rect 15473 6131 15531 6137
rect 18509 6171 18567 6177
rect 18509 6137 18521 6171
rect 18555 6168 18567 6171
rect 18874 6168 18880 6180
rect 18555 6140 18880 6168
rect 18555 6137 18567 6140
rect 18509 6131 18567 6137
rect 18708 6112 18736 6140
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 18966 6128 18972 6180
rect 19024 6168 19030 6180
rect 19334 6168 19340 6180
rect 19024 6140 19340 6168
rect 19024 6128 19030 6140
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13464 6072 14013 6100
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 15102 6100 15108 6112
rect 15063 6072 15108 6100
rect 14001 6063 14059 6069
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16577 6103 16635 6109
rect 16577 6100 16589 6103
rect 16264 6072 16589 6100
rect 16264 6060 16270 6072
rect 16577 6069 16589 6072
rect 16623 6069 16635 6103
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 16577 6063 16635 6069
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 18414 6100 18420 6112
rect 18375 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 18690 6060 18696 6112
rect 18748 6060 18754 6112
rect 19153 6103 19211 6109
rect 19153 6069 19165 6103
rect 19199 6100 19211 6103
rect 19242 6100 19248 6112
rect 19199 6072 19248 6100
rect 19199 6069 19211 6072
rect 19153 6063 19211 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 19944 6072 20177 6100
rect 19944 6060 19950 6072
rect 20165 6069 20177 6072
rect 20211 6069 20223 6103
rect 20530 6100 20536 6112
rect 20491 6072 20536 6100
rect 20165 6063 20223 6069
rect 20530 6060 20536 6072
rect 20588 6060 20594 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 5445 5899 5503 5905
rect 4028 5868 4476 5896
rect 4028 5856 4034 5868
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 4310 5831 4368 5837
rect 4310 5828 4322 5831
rect 4120 5800 4322 5828
rect 4120 5788 4126 5800
rect 4310 5797 4322 5800
rect 4356 5797 4368 5831
rect 4448 5828 4476 5868
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5994 5896 6000 5908
rect 5491 5868 6000 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 7101 5899 7159 5905
rect 7101 5865 7113 5899
rect 7147 5896 7159 5899
rect 7190 5896 7196 5908
rect 7147 5868 7196 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 7484 5828 7512 5859
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7800 5868 7941 5896
rect 7800 5856 7806 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8260 5868 8861 5896
rect 8260 5856 8266 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 10870 5896 10876 5908
rect 10183 5868 10876 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11164 5868 11836 5896
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 4448 5800 6776 5828
rect 7484 5800 8953 5828
rect 4310 5791 4368 5797
rect 5460 5772 5488 5800
rect 2590 5760 2596 5772
rect 2551 5732 2596 5760
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 4080 5732 5120 5760
rect 2682 5692 2688 5704
rect 2643 5664 2688 5692
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 2792 5624 2820 5655
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4080 5701 4108 5732
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3844 5664 4077 5692
rect 3844 5652 3850 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 5092 5692 5120 5732
rect 5442 5720 5448 5772
rect 5500 5720 5506 5772
rect 5994 5769 6000 5772
rect 5988 5760 6000 5769
rect 5955 5732 6000 5760
rect 5988 5723 6000 5732
rect 5994 5720 6000 5723
rect 6052 5720 6058 5772
rect 5626 5692 5632 5704
rect 5092 5664 5632 5692
rect 4065 5655 4123 5661
rect 5626 5652 5632 5664
rect 5684 5692 5690 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5684 5664 5733 5692
rect 5684 5652 5690 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 2556 5596 2820 5624
rect 2556 5584 2562 5596
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 3878 5556 3884 5568
rect 2271 5528 3884 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5902 5556 5908 5568
rect 5592 5528 5908 5556
rect 5592 5516 5598 5528
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 6748 5556 6776 5800
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 11164 5828 11192 5868
rect 11606 5828 11612 5840
rect 9272 5800 11192 5828
rect 11256 5800 11612 5828
rect 9272 5788 9278 5800
rect 7834 5760 7840 5772
rect 7795 5732 7840 5760
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8478 5720 8484 5772
rect 8536 5720 8542 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 11256 5769 11284 5800
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 11808 5828 11836 5868
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 13265 5899 13323 5905
rect 13265 5896 13277 5899
rect 11940 5868 13277 5896
rect 11940 5856 11946 5868
rect 13265 5865 13277 5868
rect 13311 5865 13323 5899
rect 13265 5859 13323 5865
rect 13357 5899 13415 5905
rect 13357 5865 13369 5899
rect 13403 5896 13415 5899
rect 14274 5896 14280 5908
rect 13403 5868 14280 5896
rect 13403 5865 13415 5868
rect 13357 5859 13415 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14424 5868 14657 5896
rect 14424 5856 14430 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 16206 5896 16212 5908
rect 16167 5868 16212 5896
rect 14645 5859 14703 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 17126 5896 17132 5908
rect 16684 5868 17132 5896
rect 14553 5831 14611 5837
rect 14553 5828 14565 5831
rect 11808 5800 14565 5828
rect 14553 5797 14565 5800
rect 14599 5797 14611 5831
rect 14553 5791 14611 5797
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15160 5800 16313 5828
rect 15160 5788 15166 5800
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10192 5732 10517 5760
rect 10192 5720 10198 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11497 5763 11555 5769
rect 11497 5760 11509 5763
rect 11388 5732 11509 5760
rect 11388 5720 11394 5732
rect 11497 5729 11509 5732
rect 11543 5729 11555 5763
rect 16684 5760 16712 5868
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 18104 5868 19349 5896
rect 18104 5856 18110 5868
rect 19337 5865 19349 5868
rect 19383 5865 19395 5899
rect 19337 5859 19395 5865
rect 20073 5899 20131 5905
rect 20073 5865 20085 5899
rect 20119 5896 20131 5899
rect 20530 5896 20536 5908
rect 20119 5868 20536 5896
rect 20119 5865 20131 5868
rect 20073 5859 20131 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 19245 5831 19303 5837
rect 19245 5828 19257 5831
rect 11497 5723 11555 5729
rect 14844 5732 16712 5760
rect 16776 5800 19257 5828
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7248 5664 8033 5692
rect 7248 5652 7254 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8496 5692 8524 5720
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8496 5664 9045 5692
rect 8021 5655 8079 5661
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 10376 5664 10609 5692
rect 10376 5652 10382 5664
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 10962 5692 10968 5704
rect 10827 5664 10968 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 12802 5692 12808 5704
rect 12636 5664 12808 5692
rect 12636 5633 12664 5664
rect 12802 5652 12808 5664
rect 12860 5692 12866 5704
rect 13538 5692 13544 5704
rect 12860 5664 13544 5692
rect 12860 5652 12866 5664
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 14844 5701 14872 5732
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 14829 5655 14887 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 8481 5627 8539 5633
rect 8481 5593 8493 5627
rect 8527 5624 8539 5627
rect 12621 5627 12679 5633
rect 8527 5596 11100 5624
rect 8527 5593 8539 5596
rect 8481 5587 8539 5593
rect 9766 5556 9772 5568
rect 6748 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 11072 5556 11100 5596
rect 12621 5593 12633 5627
rect 12667 5593 12679 5627
rect 12621 5587 12679 5593
rect 14185 5627 14243 5633
rect 14185 5593 14197 5627
rect 14231 5624 14243 5627
rect 16776 5624 16804 5800
rect 19245 5797 19257 5800
rect 19291 5797 19303 5831
rect 19245 5791 19303 5797
rect 17126 5720 17132 5772
rect 17184 5760 17190 5772
rect 17477 5763 17535 5769
rect 17477 5760 17489 5763
rect 17184 5732 17489 5760
rect 17184 5720 17190 5732
rect 17477 5729 17489 5732
rect 17523 5760 17535 5763
rect 17862 5760 17868 5772
rect 17523 5732 17868 5760
rect 17523 5729 17535 5732
rect 17477 5723 17535 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 18966 5692 18972 5704
rect 17221 5655 17279 5661
rect 18616 5664 18972 5692
rect 14231 5596 16804 5624
rect 14231 5593 14243 5596
rect 14185 5587 14243 5593
rect 12434 5556 12440 5568
rect 11072 5528 12440 5556
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12894 5556 12900 5568
rect 12855 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16114 5556 16120 5568
rect 15887 5528 16120 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 17236 5556 17264 5655
rect 18616 5633 18644 5664
rect 18966 5652 18972 5664
rect 19024 5692 19030 5704
rect 19521 5695 19579 5701
rect 19521 5692 19533 5695
rect 19024 5664 19533 5692
rect 19024 5652 19030 5664
rect 19521 5661 19533 5664
rect 19567 5692 19579 5695
rect 19794 5692 19800 5704
rect 19567 5664 19800 5692
rect 19567 5661 19579 5664
rect 19521 5655 19579 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 18601 5627 18659 5633
rect 18601 5593 18613 5627
rect 18647 5593 18659 5627
rect 18601 5587 18659 5593
rect 18874 5556 18880 5568
rect 16724 5528 17264 5556
rect 18835 5528 18880 5556
rect 16724 5516 16730 5528
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2682 5352 2688 5364
rect 2455 5324 2688 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 7834 5352 7840 5364
rect 7795 5324 7840 5352
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11241 5355 11299 5361
rect 11241 5352 11253 5355
rect 11204 5324 11253 5352
rect 11204 5312 11210 5324
rect 11241 5321 11253 5324
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 2222 5244 2228 5296
rect 2280 5284 2286 5296
rect 3421 5287 3479 5293
rect 2280 5256 2728 5284
rect 2280 5244 2286 5256
rect 2700 5228 2728 5256
rect 3421 5253 3433 5287
rect 3467 5284 3479 5287
rect 8478 5284 8484 5296
rect 3467 5256 8484 5284
rect 3467 5253 3479 5256
rect 3421 5247 3479 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2498 5216 2504 5228
rect 2087 5188 2504 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2740 5188 2973 5216
rect 2740 5176 2746 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 2961 5179 3019 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 7616 5188 8401 5216
rect 7616 5176 7622 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 16724 5188 18797 5216
rect 16724 5176 16730 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1636 5120 1777 5148
rect 1636 5108 1642 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3326 5148 3332 5160
rect 2823 5120 3332 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 9861 5151 9919 5157
rect 9861 5148 9873 5151
rect 7340 5120 9873 5148
rect 7340 5108 7346 5120
rect 9861 5117 9873 5120
rect 9907 5117 9919 5151
rect 9861 5111 9919 5117
rect 10128 5151 10186 5157
rect 10128 5117 10140 5151
rect 10174 5148 10186 5151
rect 10962 5148 10968 5160
rect 10174 5120 10968 5148
rect 10174 5117 10186 5120
rect 10128 5111 10186 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 12802 5157 12808 5160
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 11664 5120 12541 5148
rect 11664 5108 11670 5120
rect 12529 5117 12541 5120
rect 12575 5117 12587 5151
rect 12796 5148 12808 5157
rect 12763 5120 12808 5148
rect 12529 5111 12587 5117
rect 12796 5111 12808 5120
rect 3789 5083 3847 5089
rect 3789 5080 3801 5083
rect 1412 5052 3801 5080
rect 1412 5021 1440 5052
rect 3789 5049 3801 5052
rect 3835 5049 3847 5083
rect 3789 5043 3847 5049
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 8205 5083 8263 5089
rect 8205 5080 8217 5083
rect 6972 5052 8217 5080
rect 6972 5040 6978 5052
rect 8205 5049 8217 5052
rect 8251 5080 8263 5083
rect 12544 5080 12572 5111
rect 12802 5108 12808 5111
rect 12860 5108 12866 5160
rect 13538 5148 13544 5160
rect 12912 5120 13544 5148
rect 12912 5080 12940 5120
rect 13538 5108 13544 5120
rect 13596 5148 13602 5160
rect 14185 5151 14243 5157
rect 14185 5148 14197 5151
rect 13596 5120 14197 5148
rect 13596 5108 13602 5120
rect 14185 5117 14197 5120
rect 14231 5117 14243 5151
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 14185 5111 14243 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 13722 5080 13728 5092
rect 8251 5052 12480 5080
rect 12544 5052 12940 5080
rect 13004 5052 13728 5080
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 1397 5015 1455 5021
rect 1397 4981 1409 5015
rect 1443 4981 1455 5015
rect 1397 4975 1455 4981
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 4154 5012 4160 5024
rect 2915 4984 4160 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 7524 4984 8309 5012
rect 7524 4972 7530 4984
rect 8297 4981 8309 4984
rect 8343 4981 8355 5015
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 8297 4975 8355 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 12452 5012 12480 5052
rect 13004 5012 13032 5052
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 14430 5083 14488 5089
rect 14430 5080 14442 5083
rect 13924 5052 14442 5080
rect 12452 4984 13032 5012
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 13924 5021 13952 5052
rect 14430 5049 14442 5052
rect 14476 5049 14488 5083
rect 14430 5043 14488 5049
rect 18966 5040 18972 5092
rect 19024 5089 19030 5092
rect 19024 5083 19088 5089
rect 19024 5049 19042 5083
rect 19076 5049 19088 5083
rect 19024 5043 19088 5049
rect 19024 5040 19030 5043
rect 13909 5015 13967 5021
rect 13909 5012 13921 5015
rect 13688 4984 13921 5012
rect 13688 4972 13694 4984
rect 13909 4981 13921 4984
rect 13955 4981 13967 5015
rect 13909 4975 13967 4981
rect 15565 5015 15623 5021
rect 15565 4981 15577 5015
rect 15611 5012 15623 5015
rect 15930 5012 15936 5024
rect 15611 4984 15936 5012
rect 15611 4981 15623 4984
rect 15565 4975 15623 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 20717 5015 20775 5021
rect 20717 5012 20729 5015
rect 20312 4984 20729 5012
rect 20312 4972 20318 4984
rect 20717 4981 20729 4984
rect 20763 4981 20775 5015
rect 20717 4975 20775 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2590 4808 2596 4820
rect 2363 4780 2596 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 10134 4808 10140 4820
rect 2823 4780 10140 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2004 4644 2697 4672
rect 2004 4632 2010 4644
rect 2685 4641 2697 4644
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 1026 4564 1032 4616
rect 1084 4604 1090 4616
rect 2792 4604 2820 4771
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10778 4808 10784 4820
rect 10643 4780 10784 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11514 4808 11520 4820
rect 11011 4780 11520 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 12952 4780 13461 4808
rect 12952 4768 12958 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13449 4771 13507 4777
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15252 4780 15853 4808
rect 15252 4768 15258 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 18049 4811 18107 4817
rect 18049 4808 18061 4811
rect 17368 4780 18061 4808
rect 17368 4768 17374 4780
rect 18049 4777 18061 4780
rect 18095 4777 18107 4811
rect 18049 4771 18107 4777
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 8849 4743 8907 4749
rect 8849 4740 8861 4743
rect 6236 4712 8861 4740
rect 6236 4700 6242 4712
rect 8849 4709 8861 4712
rect 8895 4740 8907 4743
rect 12986 4740 12992 4752
rect 8895 4712 12992 4740
rect 8895 4709 8907 4712
rect 8849 4703 8907 4709
rect 12986 4700 12992 4712
rect 13044 4700 13050 4752
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 13357 4743 13415 4749
rect 13357 4740 13369 4743
rect 13320 4712 13369 4740
rect 13320 4700 13326 4712
rect 13357 4709 13369 4712
rect 13403 4709 13415 4743
rect 13357 4703 13415 4709
rect 16936 4743 16994 4749
rect 16936 4709 16948 4743
rect 16982 4740 16994 4743
rect 17034 4740 17040 4752
rect 16982 4712 17040 4740
rect 16982 4709 16994 4712
rect 16936 4703 16994 4709
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 5350 4672 5356 4684
rect 5311 4644 5356 4672
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5442 4632 5448 4684
rect 5500 4672 5506 4684
rect 8294 4672 8300 4684
rect 5500 4644 5545 4672
rect 8255 4644 8300 4672
rect 5500 4632 5506 4644
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 9674 4672 9680 4684
rect 8496 4644 9680 4672
rect 1084 4576 2820 4604
rect 2869 4607 2927 4613
rect 1084 4564 1090 4576
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 5810 4604 5816 4616
rect 5675 4576 5816 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 2682 4496 2688 4548
rect 2740 4536 2746 4548
rect 2884 4536 2912 4567
rect 5810 4564 5816 4576
rect 5868 4604 5874 4616
rect 6178 4604 6184 4616
rect 5868 4576 6184 4604
rect 5868 4564 5874 4576
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 7616 4576 8401 4604
rect 7616 4564 7622 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 2740 4508 2912 4536
rect 2740 4496 2746 4508
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3326 4536 3332 4548
rect 3016 4508 3332 4536
rect 3016 4496 3022 4508
rect 3326 4496 3332 4508
rect 3384 4536 3390 4548
rect 8496 4536 8524 4644
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 10778 4672 10784 4684
rect 9732 4644 10784 4672
rect 9732 4632 9738 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 15749 4675 15807 4681
rect 11020 4644 11192 4672
rect 11020 4632 11026 4644
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8938 4604 8944 4616
rect 8899 4576 8944 4604
rect 8573 4567 8631 4573
rect 3384 4508 8524 4536
rect 8588 4536 8616 4567
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 11164 4613 11192 4644
rect 15749 4641 15761 4675
rect 15795 4672 15807 4675
rect 16298 4672 16304 4684
rect 15795 4644 16304 4672
rect 15795 4641 15807 4644
rect 15749 4635 15807 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 19153 4675 19211 4681
rect 19153 4672 19165 4675
rect 16684 4644 19165 4672
rect 16684 4616 16712 4644
rect 19153 4641 19165 4644
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 19420 4675 19478 4681
rect 19420 4641 19432 4675
rect 19466 4672 19478 4675
rect 20162 4672 20168 4684
rect 19466 4644 20168 4672
rect 19466 4641 19478 4644
rect 19420 4635 19478 4641
rect 20162 4632 20168 4644
rect 20220 4632 20226 4684
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10652 4576 11069 4604
rect 10652 4564 10658 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4573 11207 4607
rect 13630 4604 13636 4616
rect 13591 4576 13636 4604
rect 11149 4567 11207 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 15930 4564 15936 4616
rect 15988 4604 15994 4616
rect 16666 4604 16672 4616
rect 15988 4576 16033 4604
rect 16627 4576 16672 4604
rect 15988 4564 15994 4576
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 9674 4536 9680 4548
rect 8588 4508 9680 4536
rect 3384 4496 3390 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4212 4440 4997 4468
rect 4212 4428 4218 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 4985 4431 5043 4437
rect 7929 4471 7987 4477
rect 7929 4437 7941 4471
rect 7975 4468 7987 4471
rect 8754 4468 8760 4480
rect 7975 4440 8760 4468
rect 7975 4437 7987 4440
rect 7929 4431 7987 4437
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 8849 4471 8907 4477
rect 8849 4437 8861 4471
rect 8895 4468 8907 4471
rect 9030 4468 9036 4480
rect 8895 4440 9036 4468
rect 8895 4437 8907 4440
rect 8849 4431 8907 4437
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4468 13047 4471
rect 13630 4468 13636 4480
rect 13035 4440 13636 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 18506 4428 18512 4480
rect 18564 4468 18570 4480
rect 20533 4471 20591 4477
rect 20533 4468 20545 4471
rect 18564 4440 20545 4468
rect 18564 4428 18570 4440
rect 20533 4437 20545 4440
rect 20579 4437 20591 4471
rect 20533 4431 20591 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 7558 4264 7564 4276
rect 3108 4236 6868 4264
rect 7519 4236 7564 4264
rect 3108 4224 3114 4236
rect 3970 4156 3976 4208
rect 4028 4156 4034 4208
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 5902 4196 5908 4208
rect 4120 4168 5908 4196
rect 4120 4156 4126 4168
rect 5902 4156 5908 4168
rect 5960 4156 5966 4208
rect 6730 4196 6736 4208
rect 6012 4168 6736 4196
rect 3988 4128 4016 4156
rect 4617 4131 4675 4137
rect 3988 4100 4384 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1578 4060 1584 4072
rect 1535 4032 1584 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 1756 4063 1814 4069
rect 1756 4029 1768 4063
rect 1802 4060 1814 4063
rect 2682 4060 2688 4072
rect 1802 4032 2688 4060
rect 1802 4029 1814 4032
rect 1756 4023 1814 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 4356 4069 4384 4100
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5350 4128 5356 4140
rect 5123 4100 5356 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 4632 3992 4660 4091
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 6012 4137 6040 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 6178 4128 6184 4140
rect 6139 4100 6184 4128
rect 5997 4091 6055 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6840 4128 6868 4236
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8573 4267 8631 4273
rect 8573 4264 8585 4267
rect 8352 4236 8585 4264
rect 8352 4224 8358 4236
rect 8573 4233 8585 4236
rect 8619 4233 8631 4267
rect 9401 4267 9459 4273
rect 9401 4264 9413 4267
rect 8573 4227 8631 4233
rect 9140 4236 9413 4264
rect 9140 4196 9168 4236
rect 9401 4233 9413 4236
rect 9447 4233 9459 4267
rect 9401 4227 9459 4233
rect 9493 4267 9551 4273
rect 9493 4233 9505 4267
rect 9539 4264 9551 4267
rect 10870 4264 10876 4276
rect 9539 4236 10876 4264
rect 9539 4233 9551 4236
rect 9493 4227 9551 4233
rect 10870 4224 10876 4236
rect 10928 4264 10934 4276
rect 18506 4264 18512 4276
rect 10928 4236 18512 4264
rect 10928 4224 10934 4236
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 8220 4168 9168 4196
rect 8220 4140 8248 4168
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 6840 4100 8033 4128
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8202 4128 8208 4140
rect 8115 4100 8208 4128
rect 8021 4091 8079 4097
rect 4982 4020 4988 4072
rect 5040 4060 5046 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5040 4032 5917 4060
rect 5040 4020 5046 4032
rect 5905 4029 5917 4032
rect 5951 4060 5963 4063
rect 6638 4060 6644 4072
rect 5951 4032 6644 4060
rect 5951 4029 5963 4032
rect 5905 4023 5963 4029
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 5810 3992 5816 4004
rect 3384 3964 4476 3992
rect 4632 3964 5816 3992
rect 3384 3952 3390 3964
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2556 3896 2881 3924
rect 2556 3884 2562 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 2869 3887 2927 3893
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4448 3933 4476 3964
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 8036 3992 8064 4091
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 9030 4128 9036 4140
rect 8991 4100 9036 4128
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 9140 4137 9168 4168
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 9585 4199 9643 4205
rect 9585 4196 9597 4199
rect 9364 4168 9597 4196
rect 9364 4156 9370 4168
rect 9585 4165 9597 4168
rect 9631 4165 9643 4199
rect 9585 4159 9643 4165
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 9732 4168 10272 4196
rect 9732 4156 9738 4168
rect 10244 4137 10272 4168
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 15289 4131 15347 4137
rect 15289 4097 15301 4131
rect 15335 4128 15347 4131
rect 15335 4100 15792 4128
rect 15335 4097 15347 4100
rect 15289 4091 15347 4097
rect 8938 4060 8944 4072
rect 8899 4032 8944 4060
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 15105 4063 15163 4069
rect 9048 4032 13575 4060
rect 9048 3992 9076 4032
rect 8036 3964 9076 3992
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 10410 3992 10416 4004
rect 9180 3964 10416 3992
rect 9180 3952 9186 3964
rect 10410 3952 10416 3964
rect 10468 3952 10474 4004
rect 13547 3992 13575 4032
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15470 4060 15476 4072
rect 15151 4032 15476 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15611 4032 15669 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15764 4060 15792 4100
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 18932 4100 19993 4128
rect 18932 4088 18938 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 20162 4128 20168 4140
rect 20123 4100 20168 4128
rect 19981 4091 20039 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 15930 4069 15936 4072
rect 15924 4060 15936 4069
rect 15764 4032 15936 4060
rect 15657 4023 15715 4029
rect 15924 4023 15936 4032
rect 15930 4020 15936 4023
rect 15988 4020 15994 4072
rect 18966 4060 18972 4072
rect 18927 4032 18972 4060
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19886 4060 19892 4072
rect 19847 4032 19892 4060
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 20533 4063 20591 4069
rect 20533 4029 20545 4063
rect 20579 4060 20591 4063
rect 20622 4060 20628 4072
rect 20579 4032 20628 4060
rect 20579 4029 20591 4032
rect 20533 4023 20591 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 20714 4020 20720 4072
rect 20772 4020 20778 4072
rect 17402 3992 17408 4004
rect 13547 3964 17408 3992
rect 17402 3952 17408 3964
rect 17460 3952 17466 4004
rect 20732 3992 20760 4020
rect 19168 3964 20760 3992
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3752 3896 3985 3924
rect 3752 3884 3758 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 5258 3924 5264 3936
rect 4479 3896 5264 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3924 5595 3927
rect 5626 3924 5632 3936
rect 5583 3896 5632 3924
rect 5583 3893 5595 3896
rect 5537 3887 5595 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 6052 3896 7941 3924
rect 6052 3884 6058 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 8812 3896 9413 3924
rect 8812 3884 8818 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 9493 3927 9551 3933
rect 9493 3893 9505 3927
rect 9539 3924 9551 3927
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 9539 3896 9965 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10318 3924 10324 3936
rect 10091 3896 10324 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14608 3896 14657 3924
rect 14608 3884 14614 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 15010 3924 15016 3936
rect 14971 3896 15016 3924
rect 14645 3887 14703 3893
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 15565 3927 15623 3933
rect 15565 3893 15577 3927
rect 15611 3924 15623 3927
rect 16666 3924 16672 3936
rect 15611 3896 16672 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 17034 3924 17040 3936
rect 16995 3896 17040 3924
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 18874 3924 18880 3936
rect 18748 3896 18880 3924
rect 18748 3884 18754 3896
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19168 3933 19196 3964
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3893 19211 3927
rect 19153 3887 19211 3893
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3924 19579 3927
rect 19702 3924 19708 3936
rect 19567 3896 19708 3924
rect 19567 3893 19579 3896
rect 19521 3887 19579 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 20717 3927 20775 3933
rect 20717 3924 20729 3927
rect 19852 3896 20729 3924
rect 19852 3884 19858 3896
rect 20717 3893 20729 3896
rect 20763 3893 20775 3927
rect 20717 3887 20775 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 198 3680 204 3732
rect 256 3720 262 3732
rect 2958 3720 2964 3732
rect 256 3692 2964 3720
rect 256 3680 262 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 4939 3692 5549 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 9858 3720 9864 3732
rect 6512 3692 9864 3720
rect 6512 3680 6518 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10008 3692 10701 3720
rect 10008 3680 10014 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 15102 3720 15108 3732
rect 10735 3692 15108 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 15436 3692 15669 3720
rect 15436 3680 15442 3692
rect 15657 3689 15669 3692
rect 15703 3689 15715 3723
rect 16298 3720 16304 3732
rect 16259 3692 16304 3720
rect 15657 3683 15715 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 4154 3652 4160 3664
rect 3375 3624 4160 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 4985 3655 5043 3661
rect 4985 3621 4997 3655
rect 5031 3652 5043 3655
rect 5626 3652 5632 3664
rect 5031 3624 5632 3652
rect 5031 3621 5043 3624
rect 4985 3615 5043 3621
rect 5626 3612 5632 3624
rect 5684 3612 5690 3664
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 6914 3652 6920 3664
rect 5951 3624 6920 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 5920 3584 5948 3615
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7466 3652 7472 3664
rect 7208 3624 7472 3652
rect 2884 3556 5948 3584
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2884 3380 2912 3556
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 7208 3584 7236 3624
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7828 3655 7886 3661
rect 7828 3621 7840 3655
rect 7874 3652 7886 3655
rect 8202 3652 8208 3664
rect 7874 3624 8208 3652
rect 7874 3621 7886 3624
rect 7828 3615 7886 3621
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 11977 3655 12035 3661
rect 8536 3624 11744 3652
rect 8536 3612 8542 3624
rect 6052 3556 7236 3584
rect 6052 3544 6058 3556
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7340 3556 7573 3584
rect 7340 3544 7346 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10410 3584 10416 3596
rect 10284 3556 10416 3584
rect 10284 3544 10290 3556
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 10778 3584 10784 3596
rect 10643 3556 10784 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11716 3593 11744 3624
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 12986 3652 12992 3664
rect 12023 3624 12992 3652
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 15749 3655 15807 3661
rect 15749 3652 15761 3655
rect 14608 3624 15761 3652
rect 14608 3612 14614 3624
rect 15749 3621 15761 3624
rect 15795 3621 15807 3655
rect 15749 3615 15807 3621
rect 11701 3587 11759 3593
rect 11701 3553 11713 3587
rect 11747 3553 11759 3587
rect 12434 3584 12440 3596
rect 12395 3556 12440 3584
rect 11701 3547 11759 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 13630 3584 13636 3596
rect 13591 3556 13636 3584
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 15252 3556 18061 3584
rect 15252 3544 15258 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18598 3584 18604 3596
rect 18559 3556 18604 3584
rect 18049 3547 18107 3553
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 19208 3556 19257 3584
rect 19208 3544 19214 3556
rect 19245 3553 19257 3556
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 19797 3587 19855 3593
rect 19797 3553 19809 3587
rect 19843 3584 19855 3587
rect 19978 3584 19984 3596
rect 19843 3556 19984 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 3786 3516 3792 3528
rect 3651 3488 3792 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 3436 3448 3464 3479
rect 3786 3476 3792 3488
rect 3844 3516 3850 3528
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 3844 3488 5089 3516
rect 3844 3476 3850 3488
rect 5077 3485 5089 3488
rect 5123 3516 5135 3519
rect 5350 3516 5356 3528
rect 5123 3488 5356 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 6178 3516 6184 3528
rect 6091 3488 6184 3516
rect 6178 3476 6184 3488
rect 6236 3516 6242 3528
rect 6546 3516 6552 3528
rect 6236 3488 6552 3516
rect 6236 3476 6242 3488
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9950 3516 9956 3528
rect 8812 3488 9956 3516
rect 8812 3476 8818 3488
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10318 3516 10324 3528
rect 10100 3488 10324 3516
rect 10100 3476 10106 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10870 3516 10876 3528
rect 10831 3488 10876 3516
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 13722 3516 13728 3528
rect 12759 3488 13728 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 15470 3516 15476 3528
rect 13955 3488 15476 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 17034 3516 17040 3528
rect 15979 3488 17040 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 3694 3448 3700 3460
rect 3436 3420 3700 3448
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 11054 3448 11060 3460
rect 8904 3420 11060 3448
rect 8904 3408 8910 3420
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 18233 3451 18291 3457
rect 18233 3417 18245 3451
rect 18279 3448 18291 3451
rect 21174 3448 21180 3460
rect 18279 3420 21180 3448
rect 18279 3417 18291 3420
rect 18233 3411 18291 3417
rect 21174 3408 21180 3420
rect 21232 3408 21238 3460
rect 2832 3352 2912 3380
rect 2961 3383 3019 3389
rect 2832 3340 2838 3352
rect 2961 3349 2973 3383
rect 3007 3380 3019 3383
rect 4246 3380 4252 3392
rect 3007 3352 4252 3380
rect 3007 3349 3019 3352
rect 2961 3343 3019 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4706 3380 4712 3392
rect 4571 3352 4712 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 8941 3383 8999 3389
rect 8941 3349 8953 3383
rect 8987 3380 8999 3383
rect 9674 3380 9680 3392
rect 8987 3352 9680 3380
rect 8987 3349 8999 3352
rect 8941 3343 8999 3349
rect 9674 3340 9680 3352
rect 9732 3340 9738 3392
rect 10226 3380 10232 3392
rect 10187 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 15289 3383 15347 3389
rect 15289 3349 15301 3383
rect 15335 3380 15347 3383
rect 15378 3380 15384 3392
rect 15335 3352 15384 3380
rect 15335 3349 15347 3352
rect 15289 3343 15347 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18564 3352 18797 3380
rect 18564 3340 18570 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 19208 3352 19441 3380
rect 19208 3340 19214 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 19429 3343 19487 3349
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 19981 3383 20039 3389
rect 19981 3380 19993 3383
rect 19576 3352 19993 3380
rect 19576 3340 19582 3352
rect 19981 3349 19993 3352
rect 20027 3349 20039 3383
rect 19981 3343 20039 3349
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2740 3148 2973 3176
rect 2740 3136 2746 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 5350 3176 5356 3188
rect 3752 3148 5212 3176
rect 5311 3148 5356 3176
rect 3752 3136 3758 3148
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 3786 3108 3792 3120
rect 3476 3080 3792 3108
rect 3476 3068 3482 3080
rect 3786 3068 3792 3080
rect 3844 3068 3850 3120
rect 5184 3108 5212 3148
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 8628 3148 9168 3176
rect 8628 3136 8634 3148
rect 7374 3108 7380 3120
rect 5184 3080 7380 3108
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 9140 3108 9168 3148
rect 10060 3148 10640 3176
rect 10060 3108 10088 3148
rect 9140 3080 10088 3108
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 10612 3108 10640 3148
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 15194 3176 15200 3188
rect 11112 3148 15200 3176
rect 11112 3136 11118 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 10192 3080 10548 3108
rect 10612 3080 11100 3108
rect 10192 3068 10198 3080
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7340 3012 8217 3040
rect 7340 3000 7346 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 9674 3040 9680 3052
rect 8205 3003 8263 3009
rect 9223 3012 9680 3040
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1780 2944 3924 2972
rect 1486 2864 1492 2916
rect 1544 2904 1550 2916
rect 1780 2904 1808 2944
rect 1544 2876 1808 2904
rect 1848 2907 1906 2913
rect 1544 2864 1550 2876
rect 1848 2873 1860 2907
rect 1894 2904 1906 2907
rect 3510 2904 3516 2916
rect 1894 2876 3516 2904
rect 1894 2873 1906 2876
rect 1848 2867 1906 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 3896 2904 3924 2944
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4240 2975 4298 2981
rect 4028 2944 4073 2972
rect 4028 2932 4034 2944
rect 4240 2941 4252 2975
rect 4286 2972 4298 2975
rect 6546 2972 6552 2984
rect 4286 2944 6552 2972
rect 4286 2941 4298 2944
rect 4240 2935 4298 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 8472 2975 8530 2981
rect 8472 2941 8484 2975
rect 8518 2972 8530 2975
rect 9223 2972 9251 3012
rect 9674 3000 9680 3012
rect 9732 3040 9738 3052
rect 10318 3040 10324 3052
rect 9732 3012 10324 3040
rect 9732 3000 9738 3012
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10520 3049 10548 3080
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10870 3040 10876 3052
rect 10735 3012 10876 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11072 3040 11100 3080
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 15010 3108 15016 3120
rect 11480 3080 15016 3108
rect 11480 3068 11486 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 18690 3108 18696 3120
rect 18432 3080 18696 3108
rect 11072 3012 12480 3040
rect 8518 2944 9251 2972
rect 8518 2941 8530 2944
rect 8472 2935 8530 2941
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 9364 2944 11069 2972
rect 9364 2932 9370 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11422 2972 11428 2984
rect 11057 2935 11115 2941
rect 11256 2944 11428 2972
rect 5994 2904 6000 2916
rect 3896 2876 6000 2904
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 10413 2907 10471 2913
rect 10413 2904 10425 2907
rect 8588 2876 10425 2904
rect 2406 2796 2412 2848
rect 2464 2836 2470 2848
rect 2774 2836 2780 2848
rect 2464 2808 2780 2836
rect 2464 2796 2470 2808
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 2958 2796 2964 2848
rect 3016 2836 3022 2848
rect 8588 2836 8616 2876
rect 10413 2873 10425 2876
rect 10459 2904 10471 2907
rect 11256 2904 11284 2944
rect 11422 2932 11428 2944
rect 11480 2932 11486 2984
rect 12452 2981 12480 3012
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 13078 2972 13084 2984
rect 13039 2944 13084 2972
rect 12437 2935 12495 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 13906 2972 13912 2984
rect 13863 2944 13912 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14139 2944 14565 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 14553 2935 14611 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15703 2944 16129 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 17218 2972 17224 2984
rect 17179 2944 17224 2972
rect 16117 2935 16175 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18432 2972 18460 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 18598 3000 18604 3052
rect 18656 3040 18662 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 18656 3012 19717 3040
rect 18656 3000 18662 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 18782 2972 18788 2984
rect 18095 2944 18460 2972
rect 18743 2944 18788 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 19521 2975 19579 2981
rect 19521 2972 19533 2975
rect 19300 2944 19533 2972
rect 19300 2932 19306 2944
rect 19521 2941 19533 2944
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 21634 2972 21640 2984
rect 20579 2944 21640 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 10459 2876 11284 2904
rect 11333 2907 11391 2913
rect 10459 2873 10471 2876
rect 10413 2867 10471 2873
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 12526 2904 12532 2916
rect 11379 2876 12532 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 12526 2864 12532 2876
rect 12584 2864 12590 2916
rect 13357 2907 13415 2913
rect 13357 2873 13369 2907
rect 13403 2904 13415 2907
rect 14458 2904 14464 2916
rect 13403 2876 14464 2904
rect 13403 2873 13415 2876
rect 13357 2867 13415 2873
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 17402 2864 17408 2916
rect 17460 2904 17466 2916
rect 17497 2907 17555 2913
rect 17497 2904 17509 2907
rect 17460 2876 17509 2904
rect 17460 2864 17466 2876
rect 17497 2873 17509 2876
rect 17543 2873 17555 2907
rect 18322 2904 18328 2916
rect 18283 2876 18328 2904
rect 17497 2867 17555 2873
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 18874 2864 18880 2916
rect 18932 2904 18938 2916
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 18932 2876 19073 2904
rect 18932 2864 18938 2876
rect 19061 2873 19073 2876
rect 19107 2873 19119 2907
rect 19061 2867 19119 2873
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 22554 2904 22560 2916
rect 19944 2876 22560 2904
rect 19944 2864 19950 2876
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 9582 2836 9588 2848
rect 3016 2808 8616 2836
rect 9543 2808 9588 2836
rect 3016 2796 3022 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10045 2839 10103 2845
rect 10045 2805 10057 2839
rect 10091 2836 10103 2839
rect 10134 2836 10140 2848
rect 10091 2808 10140 2836
rect 10091 2805 10103 2808
rect 10045 2799 10103 2805
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 13170 2836 13176 2848
rect 12667 2808 13176 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 14737 2839 14795 2845
rect 14737 2805 14749 2839
rect 14783 2836 14795 2839
rect 15378 2836 15384 2848
rect 14783 2808 15384 2836
rect 14783 2805 14795 2808
rect 14737 2799 14795 2805
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 16298 2836 16304 2848
rect 16259 2808 16304 2836
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19702 2836 19708 2848
rect 19024 2808 19708 2836
rect 19024 2796 19030 2808
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22094 2836 22100 2848
rect 20763 2808 22100 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 2400 2567 2458 2573
rect 2400 2533 2412 2567
rect 2446 2564 2458 2567
rect 3418 2564 3424 2576
rect 2446 2536 3424 2564
rect 2446 2533 2458 2536
rect 2400 2527 2458 2533
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 4080 2564 4108 2595
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4304 2604 4445 2632
rect 4304 2592 4310 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4706 2632 4712 2644
rect 4571 2604 4712 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 6546 2632 6552 2644
rect 6507 2604 6552 2632
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10042 2632 10048 2644
rect 9815 2604 10048 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 7193 2567 7251 2573
rect 4080 2536 6960 2564
rect 1578 2456 1584 2508
rect 1636 2496 1642 2508
rect 2133 2499 2191 2505
rect 2133 2496 2145 2499
rect 1636 2468 2145 2496
rect 1636 2456 1642 2468
rect 2133 2465 2145 2468
rect 2179 2496 2191 2499
rect 3970 2496 3976 2508
rect 2179 2468 3976 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 3970 2456 3976 2468
rect 4028 2496 4034 2508
rect 6932 2505 6960 2536
rect 7193 2533 7205 2567
rect 7239 2564 7251 2567
rect 8570 2564 8576 2576
rect 7239 2536 8576 2564
rect 7239 2533 7251 2536
rect 7193 2527 7251 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 10134 2564 10140 2576
rect 10095 2536 10140 2564
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 10744 2536 20116 2564
rect 10744 2524 10750 2536
rect 5169 2499 5227 2505
rect 5169 2496 5181 2499
rect 4028 2468 5181 2496
rect 4028 2456 4034 2468
rect 5169 2465 5181 2468
rect 5215 2465 5227 2499
rect 5169 2459 5227 2465
rect 5436 2499 5494 2505
rect 5436 2465 5448 2499
rect 5482 2496 5494 2499
rect 6917 2499 6975 2505
rect 5482 2468 6868 2496
rect 5482 2465 5494 2468
rect 5436 2459 5494 2465
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 6840 2428 6868 2468
rect 6917 2465 6929 2499
rect 6963 2465 6975 2499
rect 11698 2496 11704 2508
rect 11659 2468 11704 2496
rect 6917 2459 6975 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 12986 2456 12992 2508
rect 13044 2496 13050 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 13044 2468 13185 2496
rect 13044 2456 13050 2468
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13722 2496 13728 2508
rect 13683 2468 13728 2496
rect 13173 2459 13231 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 9582 2428 9588 2440
rect 6840 2400 9588 2428
rect 4617 2391 4675 2397
rect 3510 2320 3516 2372
rect 3568 2360 3574 2372
rect 4632 2360 4660 2391
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 14292 2428 14320 2459
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14516 2468 14841 2496
rect 14516 2456 14522 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 14829 2459 14887 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16114 2496 16120 2508
rect 16075 2468 16120 2496
rect 16114 2456 16120 2468
rect 16172 2456 16178 2508
rect 16393 2499 16451 2505
rect 16393 2465 16405 2499
rect 16439 2496 16451 2499
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 16439 2468 16865 2496
rect 16439 2465 16451 2468
rect 16393 2459 16451 2465
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 17402 2496 17408 2508
rect 17363 2468 17408 2496
rect 16853 2459 16911 2465
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 18322 2496 18328 2508
rect 18283 2468 18328 2496
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19886 2496 19892 2508
rect 19847 2468 19892 2496
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 20088 2437 20116 2536
rect 12023 2400 14320 2428
rect 20073 2431 20131 2437
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 3568 2332 4660 2360
rect 3568 2320 3574 2332
rect 17954 2320 17960 2372
rect 18012 2360 18018 2372
rect 19061 2363 19119 2369
rect 19061 2360 19073 2363
rect 18012 2332 19073 2360
rect 18012 2320 18018 2332
rect 19061 2329 19073 2332
rect 19107 2329 19119 2363
rect 19061 2323 19119 2329
rect 566 2252 572 2304
rect 624 2292 630 2304
rect 4982 2292 4988 2304
rect 624 2264 4988 2292
rect 624 2252 630 2264
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 8938 2292 8944 2304
rect 5592 2264 8944 2292
rect 5592 2252 5598 2264
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12768 2264 12817 2292
rect 12768 2252 12774 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 13538 2292 13544 2304
rect 13403 2264 13544 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 13998 2292 14004 2304
rect 13955 2264 14004 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14976 2264 15025 2292
rect 14976 2252 14982 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15838 2292 15844 2304
rect 15703 2264 15844 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 16666 2252 16672 2304
rect 16724 2292 16730 2304
rect 17037 2295 17095 2301
rect 17037 2292 17049 2295
rect 16724 2264 17049 2292
rect 16724 2252 16730 2264
rect 17037 2261 17049 2264
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17184 2264 17601 2292
rect 17184 2252 17190 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 17736 2264 18521 2292
rect 17736 2252 17742 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 8754 1408 8760 1420
rect 6052 1380 8760 1408
rect 6052 1368 6058 1380
rect 8754 1368 8760 1380
rect 8812 1368 8818 1420
rect 11330 1232 11336 1284
rect 11388 1272 11394 1284
rect 12158 1272 12164 1284
rect 11388 1244 12164 1272
rect 11388 1232 11394 1244
rect 12158 1232 12164 1244
rect 12216 1232 12222 1284
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 5718 1068 5724 1080
rect 4120 1040 5724 1068
rect 4120 1028 4126 1040
rect 5718 1028 5724 1040
rect 5776 1028 5782 1080
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 7196 19864 7248 19916
rect 15200 19864 15252 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20076 19864 20128 19916
rect 5172 19796 5224 19848
rect 15292 19796 15344 19848
rect 16028 19839 16080 19848
rect 16028 19805 16037 19839
rect 16037 19805 16071 19839
rect 16071 19805 16080 19839
rect 16028 19796 16080 19805
rect 2964 19728 3016 19780
rect 17960 19660 18012 19712
rect 20628 19660 20680 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 2044 19499 2096 19508
rect 2044 19465 2053 19499
rect 2053 19465 2087 19499
rect 2087 19465 2096 19499
rect 2044 19456 2096 19465
rect 4068 19456 4120 19508
rect 16028 19456 16080 19508
rect 19708 19456 19760 19508
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 5080 19252 5132 19304
rect 3608 19184 3660 19236
rect 7012 19252 7064 19304
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 10140 19295 10192 19304
rect 2872 19116 2924 19168
rect 4160 19116 4212 19168
rect 5724 19116 5776 19168
rect 7656 19184 7708 19236
rect 7748 19184 7800 19236
rect 10140 19261 10149 19295
rect 10149 19261 10183 19295
rect 10183 19261 10192 19295
rect 10140 19252 10192 19261
rect 10784 19252 10836 19304
rect 14464 19295 14516 19304
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 14464 19252 14516 19261
rect 12716 19227 12768 19236
rect 7380 19116 7432 19168
rect 7564 19159 7616 19168
rect 7564 19125 7573 19159
rect 7573 19125 7607 19159
rect 7607 19125 7616 19159
rect 7564 19116 7616 19125
rect 9864 19159 9916 19168
rect 9864 19125 9873 19159
rect 9873 19125 9907 19159
rect 9907 19125 9916 19159
rect 11520 19159 11572 19168
rect 9864 19116 9916 19125
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 17132 19252 17184 19304
rect 19156 19252 19208 19304
rect 19340 19252 19392 19304
rect 19708 19252 19760 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 15568 19184 15620 19236
rect 19064 19159 19116 19168
rect 19064 19125 19073 19159
rect 19073 19125 19107 19159
rect 19107 19125 19116 19159
rect 19064 19116 19116 19125
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 2780 18912 2832 18964
rect 3056 18955 3108 18964
rect 3056 18921 3065 18955
rect 3065 18921 3099 18955
rect 3099 18921 3108 18955
rect 3056 18912 3108 18921
rect 7748 18912 7800 18964
rect 2504 18776 2556 18828
rect 4988 18819 5040 18828
rect 4988 18785 5022 18819
rect 5022 18785 5040 18819
rect 4988 18776 5040 18785
rect 7288 18776 7340 18828
rect 3148 18708 3200 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 5632 18572 5684 18624
rect 6092 18615 6144 18624
rect 6092 18581 6101 18615
rect 6101 18581 6135 18615
rect 6135 18581 6144 18615
rect 6092 18572 6144 18581
rect 8208 18912 8260 18964
rect 10140 18912 10192 18964
rect 19248 18912 19300 18964
rect 10324 18844 10376 18896
rect 13544 18844 13596 18896
rect 16028 18887 16080 18896
rect 16028 18853 16062 18887
rect 16062 18853 16080 18887
rect 16028 18844 16080 18853
rect 19984 18844 20036 18896
rect 9680 18776 9732 18828
rect 11520 18776 11572 18828
rect 10784 18708 10836 18760
rect 9956 18640 10008 18692
rect 8208 18572 8260 18624
rect 8392 18615 8444 18624
rect 8392 18581 8401 18615
rect 8401 18581 8435 18615
rect 8435 18581 8444 18615
rect 8392 18572 8444 18581
rect 13636 18776 13688 18828
rect 14464 18776 14516 18828
rect 16580 18776 16632 18828
rect 19524 18776 19576 18828
rect 19616 18776 19668 18828
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 15568 18708 15620 18760
rect 12716 18640 12768 18692
rect 15200 18640 15252 18692
rect 14188 18572 14240 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 7012 18411 7064 18420
rect 1952 18343 2004 18352
rect 1952 18309 1961 18343
rect 1961 18309 1995 18343
rect 1995 18309 2004 18343
rect 1952 18300 2004 18309
rect 3148 18164 3200 18216
rect 4160 18164 4212 18216
rect 1860 18096 1912 18148
rect 6000 18096 6052 18148
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 4988 18071 5040 18080
rect 3056 18028 3108 18037
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 13636 18368 13688 18420
rect 20076 18368 20128 18420
rect 8392 18300 8444 18352
rect 15108 18300 15160 18352
rect 20168 18343 20220 18352
rect 20168 18309 20177 18343
rect 20177 18309 20211 18343
rect 20211 18309 20220 18343
rect 20168 18300 20220 18309
rect 7380 18207 7432 18216
rect 7380 18173 7389 18207
rect 7389 18173 7423 18207
rect 7423 18173 7432 18207
rect 7380 18164 7432 18173
rect 7656 18232 7708 18284
rect 8208 18232 8260 18284
rect 10048 18232 10100 18284
rect 13728 18232 13780 18284
rect 9864 18164 9916 18216
rect 14188 18164 14240 18216
rect 16488 18164 16540 18216
rect 16856 18164 16908 18216
rect 17868 18164 17920 18216
rect 17960 18164 18012 18216
rect 19524 18164 19576 18216
rect 20076 18164 20128 18216
rect 8760 18096 8812 18148
rect 11060 18096 11112 18148
rect 9772 18028 9824 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 10416 18028 10468 18080
rect 13728 18071 13780 18080
rect 13728 18037 13737 18071
rect 13737 18037 13771 18071
rect 13771 18037 13780 18071
rect 13728 18028 13780 18037
rect 15752 18096 15804 18148
rect 15476 18071 15528 18080
rect 15476 18037 15485 18071
rect 15485 18037 15519 18071
rect 15519 18037 15528 18071
rect 15476 18028 15528 18037
rect 16764 18028 16816 18080
rect 18972 18028 19024 18080
rect 20628 18028 20680 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 2596 17824 2648 17876
rect 2964 17867 3016 17876
rect 2964 17833 2973 17867
rect 2973 17833 3007 17867
rect 3007 17833 3016 17867
rect 2964 17824 3016 17833
rect 4988 17824 5040 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 11060 17824 11112 17876
rect 13728 17824 13780 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15752 17867 15804 17876
rect 15752 17833 15761 17867
rect 15761 17833 15795 17867
rect 15795 17833 15804 17867
rect 15752 17824 15804 17833
rect 19064 17824 19116 17876
rect 19432 17824 19484 17876
rect 4160 17756 4212 17808
rect 3332 17731 3384 17740
rect 3332 17697 3341 17731
rect 3341 17697 3375 17731
rect 3375 17697 3384 17731
rect 3332 17688 3384 17697
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3608 17663 3660 17672
rect 3608 17629 3617 17663
rect 3617 17629 3651 17663
rect 3651 17629 3660 17663
rect 3608 17620 3660 17629
rect 2044 17484 2096 17536
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 5632 17756 5684 17808
rect 8024 17688 8076 17740
rect 9864 17688 9916 17740
rect 15108 17756 15160 17808
rect 16948 17756 17000 17808
rect 20536 17756 20588 17808
rect 9772 17620 9824 17672
rect 10324 17688 10376 17740
rect 13084 17688 13136 17740
rect 17316 17688 17368 17740
rect 12716 17663 12768 17672
rect 6736 17552 6788 17604
rect 7288 17552 7340 17604
rect 10048 17552 10100 17604
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 15568 17620 15620 17672
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 13544 17552 13596 17604
rect 10140 17484 10192 17536
rect 17776 17484 17828 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 7564 17280 7616 17332
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 15476 17280 15528 17332
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 3608 17144 3660 17196
rect 6460 17144 6512 17196
rect 7288 17144 7340 17196
rect 8760 17144 8812 17196
rect 12072 17144 12124 17196
rect 16488 17144 16540 17196
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 3516 17076 3568 17128
rect 10784 17076 10836 17128
rect 7012 17008 7064 17060
rect 8392 17051 8444 17060
rect 8392 17017 8401 17051
rect 8401 17017 8435 17051
rect 8435 17017 8444 17051
rect 8392 17008 8444 17017
rect 10968 17051 11020 17060
rect 10968 17017 11002 17051
rect 11002 17017 11020 17051
rect 11704 17076 11756 17128
rect 17776 17076 17828 17128
rect 20168 17076 20220 17128
rect 10968 17008 11020 17017
rect 12624 17008 12676 17060
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 4252 16940 4304 16992
rect 4712 16940 4764 16992
rect 4896 16940 4948 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 6644 16940 6696 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 13912 17008 13964 17060
rect 17684 17008 17736 17060
rect 19432 17008 19484 17060
rect 19708 17008 19760 17060
rect 15292 16940 15344 16992
rect 16488 16983 16540 16992
rect 16488 16949 16497 16983
rect 16497 16949 16531 16983
rect 16531 16949 16540 16983
rect 16488 16940 16540 16949
rect 16948 16940 17000 16992
rect 20628 16940 20680 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 2780 16736 2832 16788
rect 2872 16736 2924 16788
rect 3332 16736 3384 16788
rect 8760 16736 8812 16788
rect 12072 16736 12124 16788
rect 15292 16779 15344 16788
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 2320 16643 2372 16652
rect 2320 16609 2329 16643
rect 2329 16609 2363 16643
rect 2363 16609 2372 16643
rect 2320 16600 2372 16609
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 4804 16600 4856 16652
rect 5356 16643 5408 16652
rect 5356 16609 5390 16643
rect 5390 16609 5408 16643
rect 8208 16668 8260 16720
rect 12440 16668 12492 16720
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 19892 16779 19944 16788
rect 19892 16745 19901 16779
rect 19901 16745 19935 16779
rect 19935 16745 19944 16779
rect 19892 16736 19944 16745
rect 16856 16668 16908 16720
rect 19800 16668 19852 16720
rect 5356 16600 5408 16609
rect 9588 16600 9640 16652
rect 14096 16600 14148 16652
rect 16028 16600 16080 16652
rect 16488 16600 16540 16652
rect 17592 16600 17644 16652
rect 19984 16600 20036 16652
rect 11152 16532 11204 16584
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 1952 16507 2004 16516
rect 1952 16473 1961 16507
rect 1961 16473 1995 16507
rect 1995 16473 2004 16507
rect 1952 16464 2004 16473
rect 10968 16464 11020 16516
rect 12624 16532 12676 16584
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 11796 16396 11848 16448
rect 17960 16464 18012 16516
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 5264 16192 5316 16244
rect 6736 16192 6788 16244
rect 4896 16124 4948 16176
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 5356 16056 5408 16108
rect 6460 16056 6512 16108
rect 9588 16192 9640 16244
rect 11704 16192 11756 16244
rect 9956 16124 10008 16176
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 12440 16099 12492 16108
rect 12440 16065 12449 16099
rect 12449 16065 12483 16099
rect 12483 16065 12492 16099
rect 12440 16056 12492 16065
rect 6920 15988 6972 16040
rect 8208 15988 8260 16040
rect 1768 15920 1820 15972
rect 5448 15963 5500 15972
rect 5448 15929 5457 15963
rect 5457 15929 5491 15963
rect 5491 15929 5500 15963
rect 5448 15920 5500 15929
rect 15384 16192 15436 16244
rect 19432 16235 19484 16244
rect 19432 16201 19441 16235
rect 19441 16201 19475 16235
rect 19475 16201 19484 16235
rect 19432 16192 19484 16201
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 10232 15920 10284 15972
rect 10968 15920 11020 15972
rect 11980 15920 12032 15972
rect 5172 15852 5224 15904
rect 6828 15852 6880 15904
rect 7380 15852 7432 15904
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 11428 15852 11480 15904
rect 14004 15920 14056 15972
rect 14096 15920 14148 15972
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 15936 15988 15988 16040
rect 17776 15988 17828 16040
rect 20536 16031 20588 16040
rect 17224 15920 17276 15972
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 19984 15920 20036 15972
rect 20260 15920 20312 15972
rect 19064 15852 19116 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 5264 15648 5316 15700
rect 5356 15648 5408 15700
rect 8484 15648 8536 15700
rect 10140 15691 10192 15700
rect 10140 15657 10149 15691
rect 10149 15657 10183 15691
rect 10183 15657 10192 15691
rect 10140 15648 10192 15657
rect 2688 15580 2740 15632
rect 6736 15580 6788 15632
rect 6828 15580 6880 15632
rect 3240 15308 3292 15360
rect 4804 15512 4856 15564
rect 7104 15512 7156 15564
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9956 15580 10008 15632
rect 11428 15648 11480 15700
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 13912 15691 13964 15700
rect 11336 15580 11388 15632
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 14004 15648 14056 15700
rect 16672 15648 16724 15700
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 20536 15648 20588 15700
rect 18512 15580 18564 15632
rect 19708 15580 19760 15632
rect 9588 15444 9640 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 15384 15512 15436 15564
rect 15936 15512 15988 15564
rect 16396 15512 16448 15564
rect 18604 15555 18656 15564
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 18696 15555 18748 15564
rect 18696 15521 18705 15555
rect 18705 15521 18739 15555
rect 18739 15521 18748 15555
rect 18696 15512 18748 15521
rect 20260 15555 20312 15564
rect 20260 15521 20269 15555
rect 20269 15521 20303 15555
rect 20303 15521 20312 15555
rect 20260 15512 20312 15521
rect 12072 15487 12124 15496
rect 12072 15453 12081 15487
rect 12081 15453 12115 15487
rect 12115 15453 12124 15487
rect 12072 15444 12124 15453
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 18880 15444 18932 15496
rect 11980 15376 12032 15428
rect 4252 15308 4304 15360
rect 4804 15308 4856 15360
rect 7288 15308 7340 15360
rect 8208 15308 8260 15360
rect 8576 15308 8628 15360
rect 10140 15308 10192 15360
rect 12900 15308 12952 15360
rect 19432 15376 19484 15428
rect 19984 15444 20036 15496
rect 20352 15444 20404 15496
rect 17960 15308 18012 15360
rect 19984 15308 20036 15360
rect 20444 15351 20496 15360
rect 20444 15317 20453 15351
rect 20453 15317 20487 15351
rect 20487 15317 20496 15351
rect 20444 15308 20496 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 1952 15147 2004 15156
rect 1952 15113 1961 15147
rect 1961 15113 1995 15147
rect 1995 15113 2004 15147
rect 1952 15104 2004 15113
rect 4252 15104 4304 15156
rect 8208 15104 8260 15156
rect 8392 15104 8444 15156
rect 13084 15104 13136 15156
rect 9588 14968 9640 15020
rect 18512 15104 18564 15156
rect 18696 15104 18748 15156
rect 7288 14943 7340 14952
rect 3792 14875 3844 14884
rect 3792 14841 3826 14875
rect 3826 14841 3844 14875
rect 3792 14832 3844 14841
rect 7288 14909 7322 14943
rect 7322 14909 7340 14943
rect 7288 14900 7340 14909
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 15016 14900 15068 14952
rect 19248 15036 19300 15088
rect 17224 14968 17276 15020
rect 18604 14968 18656 15020
rect 17960 14900 18012 14952
rect 19064 14900 19116 14952
rect 19340 14900 19392 14952
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 7564 14832 7616 14884
rect 10140 14832 10192 14884
rect 13728 14875 13780 14884
rect 13728 14841 13762 14875
rect 13762 14841 13780 14875
rect 13728 14832 13780 14841
rect 19708 14832 19760 14884
rect 20260 14875 20312 14884
rect 20260 14841 20269 14875
rect 20269 14841 20303 14875
rect 20303 14841 20312 14875
rect 20260 14832 20312 14841
rect 2688 14764 2740 14816
rect 8300 14764 8352 14816
rect 8484 14764 8536 14816
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 15108 14764 15160 14816
rect 16396 14764 16448 14816
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 19064 14764 19116 14816
rect 19800 14764 19852 14816
rect 20904 14807 20956 14816
rect 20904 14773 20913 14807
rect 20913 14773 20947 14807
rect 20947 14773 20956 14807
rect 20904 14764 20956 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 6920 14560 6972 14612
rect 15016 14560 15068 14612
rect 15384 14560 15436 14612
rect 19892 14603 19944 14612
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 6092 14492 6144 14544
rect 7748 14492 7800 14544
rect 1676 14424 1728 14476
rect 2136 14424 2188 14476
rect 4804 14424 4856 14476
rect 5356 14467 5408 14476
rect 5356 14433 5365 14467
rect 5365 14433 5399 14467
rect 5399 14433 5408 14467
rect 5356 14424 5408 14433
rect 8392 14424 8444 14476
rect 12808 14492 12860 14544
rect 13544 14492 13596 14544
rect 11888 14424 11940 14476
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 6828 14356 6880 14408
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 2596 14263 2648 14272
rect 2596 14229 2605 14263
rect 2605 14229 2639 14263
rect 2639 14229 2648 14263
rect 2596 14220 2648 14229
rect 3884 14220 3936 14272
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 7288 14288 7340 14340
rect 10508 14356 10560 14408
rect 13452 14424 13504 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 20260 14467 20312 14476
rect 20260 14433 20269 14467
rect 20269 14433 20303 14467
rect 20303 14433 20312 14467
rect 20260 14424 20312 14433
rect 14372 14399 14424 14408
rect 10600 14220 10652 14272
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 13728 14288 13780 14340
rect 17224 14356 17276 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 18880 14288 18932 14340
rect 12624 14220 12676 14272
rect 13176 14220 13228 14272
rect 14832 14220 14884 14272
rect 16856 14220 16908 14272
rect 19432 14220 19484 14272
rect 20444 14263 20496 14272
rect 20444 14229 20453 14263
rect 20453 14229 20487 14263
rect 20487 14229 20496 14263
rect 20444 14220 20496 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2136 14059 2188 14068
rect 2136 14025 2145 14059
rect 2145 14025 2179 14059
rect 2179 14025 2188 14059
rect 2136 14016 2188 14025
rect 3056 14016 3108 14068
rect 5356 14016 5408 14068
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 6920 14016 6972 14068
rect 7196 14016 7248 14068
rect 8484 14016 8536 14068
rect 8944 14016 8996 14068
rect 9588 14016 9640 14068
rect 9956 14016 10008 14068
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10140 14016 10192 14025
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 14832 14016 14884 14068
rect 3332 13991 3384 14000
rect 3332 13957 3341 13991
rect 3341 13957 3375 13991
rect 3375 13957 3384 13991
rect 3332 13948 3384 13957
rect 8300 13948 8352 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 6736 13880 6788 13932
rect 9220 13880 9272 13932
rect 2596 13812 2648 13864
rect 6092 13812 6144 13864
rect 7104 13812 7156 13864
rect 10232 13880 10284 13932
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 14096 13880 14148 13932
rect 6276 13744 6328 13796
rect 9404 13744 9456 13796
rect 10508 13787 10560 13796
rect 10508 13753 10517 13787
rect 10517 13753 10551 13787
rect 10551 13753 10560 13787
rect 10508 13744 10560 13753
rect 10600 13787 10652 13796
rect 10600 13753 10609 13787
rect 10609 13753 10643 13787
rect 10643 13753 10652 13787
rect 10600 13744 10652 13753
rect 2228 13676 2280 13728
rect 2596 13719 2648 13728
rect 2596 13685 2605 13719
rect 2605 13685 2639 13719
rect 2639 13685 2648 13719
rect 4252 13719 4304 13728
rect 2596 13676 2648 13685
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 7196 13719 7248 13728
rect 4344 13676 4396 13685
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 8944 13676 8996 13728
rect 9312 13676 9364 13728
rect 9680 13676 9732 13728
rect 11612 13719 11664 13728
rect 11612 13685 11621 13719
rect 11621 13685 11655 13719
rect 11655 13685 11664 13719
rect 11612 13676 11664 13685
rect 11796 13676 11848 13728
rect 13452 13744 13504 13796
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 13820 13676 13872 13728
rect 15384 13812 15436 13864
rect 16948 13812 17000 13864
rect 18604 14016 18656 14068
rect 20628 13948 20680 14000
rect 19064 13880 19116 13932
rect 19248 13880 19300 13932
rect 15016 13744 15068 13796
rect 19708 13744 19760 13796
rect 16120 13676 16172 13728
rect 17040 13676 17092 13728
rect 19432 13676 19484 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2228 13515 2280 13524
rect 2228 13481 2237 13515
rect 2237 13481 2271 13515
rect 2271 13481 2280 13515
rect 2228 13472 2280 13481
rect 4344 13472 4396 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 2872 13404 2924 13456
rect 9680 13472 9732 13524
rect 13636 13472 13688 13524
rect 16764 13472 16816 13524
rect 17224 13472 17276 13524
rect 17500 13472 17552 13524
rect 18512 13472 18564 13524
rect 5540 13336 5592 13388
rect 6828 13336 6880 13388
rect 9864 13404 9916 13456
rect 11612 13404 11664 13456
rect 15016 13404 15068 13456
rect 9220 13336 9272 13388
rect 2412 13268 2464 13320
rect 2964 13268 3016 13320
rect 4988 13311 5040 13320
rect 4988 13277 4997 13311
rect 4997 13277 5031 13311
rect 5031 13277 5040 13311
rect 4988 13268 5040 13277
rect 3792 13200 3844 13252
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 9312 13268 9364 13320
rect 11888 13268 11940 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 14096 13336 14148 13388
rect 17960 13336 18012 13388
rect 18512 13336 18564 13388
rect 18880 13336 18932 13388
rect 15384 13268 15436 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16120 13311 16172 13320
rect 16120 13277 16129 13311
rect 16129 13277 16163 13311
rect 16163 13277 16172 13311
rect 16120 13268 16172 13277
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17868 13268 17920 13320
rect 5080 13132 5132 13184
rect 16396 13200 16448 13252
rect 18696 13268 18748 13320
rect 7380 13132 7432 13184
rect 8300 13132 8352 13184
rect 14372 13132 14424 13184
rect 14464 13132 14516 13184
rect 16580 13132 16632 13184
rect 16764 13132 16816 13184
rect 19064 13200 19116 13252
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 7104 12971 7156 12980
rect 7104 12937 7113 12971
rect 7113 12937 7147 12971
rect 7147 12937 7156 12971
rect 7104 12928 7156 12937
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 14464 12928 14516 12980
rect 15936 12928 15988 12980
rect 16580 12928 16632 12980
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 5264 12792 5316 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 6184 12792 6236 12844
rect 7932 12835 7984 12844
rect 3148 12724 3200 12776
rect 3424 12724 3476 12776
rect 5080 12724 5132 12776
rect 7104 12724 7156 12776
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8208 12792 8260 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 12164 12792 12216 12844
rect 12440 12724 12492 12776
rect 4068 12656 4120 12708
rect 12532 12656 12584 12708
rect 13452 12792 13504 12844
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 17408 12860 17460 12912
rect 17868 12928 17920 12980
rect 20352 12928 20404 12980
rect 15108 12792 15160 12844
rect 16396 12792 16448 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 18696 12792 18748 12844
rect 19064 12792 19116 12844
rect 20352 12792 20404 12844
rect 18880 12724 18932 12776
rect 19800 12724 19852 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 17040 12656 17092 12708
rect 17592 12656 17644 12708
rect 20628 12699 20680 12708
rect 20628 12665 20637 12699
rect 20637 12665 20671 12699
rect 20671 12665 20680 12699
rect 20628 12656 20680 12665
rect 6644 12588 6696 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 11888 12588 11940 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 13544 12588 13596 12640
rect 13912 12588 13964 12640
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 17776 12588 17828 12640
rect 18788 12631 18840 12640
rect 18788 12597 18797 12631
rect 18797 12597 18831 12631
rect 18831 12597 18840 12631
rect 20260 12631 20312 12640
rect 18788 12588 18840 12597
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2596 12384 2648 12436
rect 5908 12384 5960 12436
rect 6276 12384 6328 12436
rect 7196 12384 7248 12436
rect 2596 12291 2648 12300
rect 2596 12257 2605 12291
rect 2605 12257 2639 12291
rect 2639 12257 2648 12291
rect 2596 12248 2648 12257
rect 4712 12248 4764 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 2504 12180 2556 12232
rect 2964 12180 3016 12232
rect 3700 12180 3752 12232
rect 3056 12112 3108 12164
rect 5632 12180 5684 12232
rect 5908 12248 5960 12300
rect 6920 12248 6972 12300
rect 10968 12384 11020 12436
rect 15752 12384 15804 12436
rect 16948 12384 17000 12436
rect 17776 12384 17828 12436
rect 17960 12384 18012 12436
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 8668 12316 8720 12368
rect 11244 12316 11296 12368
rect 8576 12248 8628 12300
rect 9772 12248 9824 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 7472 12180 7524 12232
rect 7656 12180 7708 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 10968 12180 11020 12232
rect 12072 12316 12124 12368
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 12440 12248 12492 12300
rect 12716 12248 12768 12300
rect 13452 12291 13504 12300
rect 13452 12257 13486 12291
rect 13486 12257 13504 12291
rect 13452 12248 13504 12257
rect 15200 12316 15252 12368
rect 15292 12248 15344 12300
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 5816 12087 5868 12096
rect 5816 12053 5825 12087
rect 5825 12053 5859 12087
rect 5859 12053 5868 12087
rect 5816 12044 5868 12053
rect 7012 12044 7064 12096
rect 7288 12044 7340 12096
rect 8852 12112 8904 12164
rect 12992 12180 13044 12232
rect 13176 12223 13228 12232
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 18696 12316 18748 12368
rect 19064 12316 19116 12368
rect 12808 12112 12860 12164
rect 17684 12180 17736 12232
rect 20352 12248 20404 12300
rect 18880 12180 18932 12232
rect 10968 12044 11020 12096
rect 11612 12044 11664 12096
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 16028 12112 16080 12164
rect 17868 12112 17920 12164
rect 20168 12044 20220 12096
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 4160 11840 4212 11892
rect 4252 11840 4304 11892
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 8760 11840 8812 11892
rect 8852 11840 8904 11892
rect 10784 11840 10836 11892
rect 12348 11840 12400 11892
rect 3700 11815 3752 11824
rect 3700 11781 3709 11815
rect 3709 11781 3743 11815
rect 3743 11781 3752 11815
rect 3700 11772 3752 11781
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 4988 11772 5040 11824
rect 5632 11704 5684 11756
rect 6368 11704 6420 11756
rect 3056 11636 3108 11688
rect 5816 11636 5868 11688
rect 7012 11636 7064 11688
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 9588 11772 9640 11824
rect 11152 11772 11204 11824
rect 8208 11704 8260 11756
rect 9772 11704 9824 11756
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 13452 11840 13504 11892
rect 19248 11840 19300 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 11888 11679 11940 11688
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 4068 11568 4120 11620
rect 15292 11704 15344 11756
rect 4804 11500 4856 11552
rect 6736 11500 6788 11552
rect 7196 11500 7248 11552
rect 7748 11500 7800 11552
rect 8944 11543 8996 11552
rect 8944 11509 8953 11543
rect 8953 11509 8987 11543
rect 8987 11509 8996 11543
rect 10232 11543 10284 11552
rect 8944 11500 8996 11509
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 11704 11500 11756 11552
rect 12072 11500 12124 11552
rect 16948 11636 17000 11688
rect 18880 11704 18932 11756
rect 12992 11568 13044 11620
rect 16672 11568 16724 11620
rect 17592 11568 17644 11620
rect 18696 11568 18748 11620
rect 18880 11568 18932 11620
rect 19248 11611 19300 11620
rect 19248 11577 19282 11611
rect 19282 11577 19300 11611
rect 19248 11568 19300 11577
rect 13176 11500 13228 11552
rect 13268 11500 13320 11552
rect 17040 11500 17092 11552
rect 17960 11500 18012 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2504 11339 2556 11348
rect 2504 11305 2513 11339
rect 2513 11305 2547 11339
rect 2547 11305 2556 11339
rect 2504 11296 2556 11305
rect 7104 11296 7156 11348
rect 8208 11296 8260 11348
rect 8852 11296 8904 11348
rect 9312 11296 9364 11348
rect 12532 11296 12584 11348
rect 13268 11296 13320 11348
rect 13820 11296 13872 11348
rect 17316 11296 17368 11348
rect 18604 11296 18656 11348
rect 2964 11228 3016 11280
rect 3516 11228 3568 11280
rect 5448 11228 5500 11280
rect 7472 11228 7524 11280
rect 9588 11228 9640 11280
rect 1952 11160 2004 11212
rect 5724 11160 5776 11212
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 7104 11160 7156 11212
rect 7748 11160 7800 11212
rect 10692 11160 10744 11212
rect 15660 11203 15712 11212
rect 2780 11024 2832 11076
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 5448 11135 5500 11144
rect 3056 11092 3108 11101
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 5448 11092 5500 11101
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6736 11092 6788 11144
rect 3240 11024 3292 11076
rect 7288 11024 7340 11076
rect 4160 10956 4212 11008
rect 7104 10956 7156 11008
rect 7564 10956 7616 11008
rect 8392 11092 8444 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 17500 11203 17552 11212
rect 17500 11169 17534 11203
rect 17534 11169 17552 11203
rect 17500 11160 17552 11169
rect 18512 11160 18564 11212
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 16856 11092 16908 11144
rect 18696 11092 18748 11144
rect 19248 11024 19300 11076
rect 8944 10956 8996 11008
rect 15476 10956 15528 11008
rect 19616 10956 19668 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2596 10752 2648 10804
rect 4068 10752 4120 10804
rect 4988 10752 5040 10804
rect 5632 10752 5684 10804
rect 6460 10752 6512 10804
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3792 10616 3844 10668
rect 4160 10548 4212 10600
rect 13912 10752 13964 10804
rect 15660 10752 15712 10804
rect 18512 10752 18564 10804
rect 13176 10684 13228 10736
rect 14464 10684 14516 10736
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7564 10616 7616 10668
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 18696 10684 18748 10736
rect 16212 10616 16264 10668
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 19616 10616 19668 10668
rect 20536 10616 20588 10668
rect 2780 10480 2832 10532
rect 3884 10480 3936 10532
rect 3976 10480 4028 10532
rect 9864 10548 9916 10600
rect 10508 10591 10560 10600
rect 10508 10557 10542 10591
rect 10542 10557 10560 10591
rect 10508 10548 10560 10557
rect 10784 10548 10836 10600
rect 17408 10591 17460 10600
rect 5448 10480 5500 10532
rect 3608 10412 3660 10464
rect 7196 10455 7248 10464
rect 7196 10421 7205 10455
rect 7205 10421 7239 10455
rect 7239 10421 7248 10455
rect 7196 10412 7248 10421
rect 7380 10412 7432 10464
rect 11704 10412 11756 10464
rect 13912 10412 13964 10464
rect 17408 10557 17417 10591
rect 17417 10557 17451 10591
rect 17451 10557 17460 10591
rect 17408 10548 17460 10557
rect 17960 10548 18012 10600
rect 18880 10548 18932 10600
rect 19984 10480 20036 10532
rect 16672 10412 16724 10464
rect 18696 10412 18748 10464
rect 19064 10412 19116 10464
rect 19524 10412 19576 10464
rect 20076 10455 20128 10464
rect 20076 10421 20085 10455
rect 20085 10421 20119 10455
rect 20119 10421 20128 10455
rect 20076 10412 20128 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 2872 10208 2924 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 6368 10208 6420 10260
rect 7380 10208 7432 10260
rect 9680 10208 9732 10260
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 10232 10208 10284 10260
rect 15752 10208 15804 10260
rect 17500 10208 17552 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20076 10208 20128 10260
rect 4068 10140 4120 10192
rect 15200 10140 15252 10192
rect 15384 10140 15436 10192
rect 17960 10140 18012 10192
rect 1952 10072 2004 10124
rect 6552 10072 6604 10124
rect 6644 10072 6696 10124
rect 7564 10115 7616 10124
rect 3792 10004 3844 10056
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 5080 10004 5132 10056
rect 7564 10081 7587 10115
rect 7587 10081 7616 10115
rect 7564 10072 7616 10081
rect 9772 10072 9824 10124
rect 10784 10072 10836 10124
rect 11704 10115 11756 10124
rect 11704 10081 11738 10115
rect 11738 10081 11756 10115
rect 11704 10072 11756 10081
rect 13176 10072 13228 10124
rect 14096 10072 14148 10124
rect 17500 10072 17552 10124
rect 20260 10072 20312 10124
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10140 9936 10192 9988
rect 10784 9936 10836 9988
rect 6368 9868 6420 9920
rect 6552 9868 6604 9920
rect 10968 9868 11020 9920
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16856 10047 16908 10056
rect 14556 9936 14608 9988
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 20168 10047 20220 10056
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 20536 10004 20588 10056
rect 12532 9868 12584 9920
rect 12716 9868 12768 9920
rect 14004 9868 14056 9920
rect 15200 9868 15252 9920
rect 15292 9868 15344 9920
rect 16580 9868 16632 9920
rect 19616 9911 19668 9920
rect 19616 9877 19625 9911
rect 19625 9877 19659 9911
rect 19659 9877 19668 9911
rect 19616 9868 19668 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 7656 9664 7708 9716
rect 8300 9664 8352 9716
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 6276 9596 6328 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 3332 9460 3384 9512
rect 4068 9460 4120 9512
rect 7288 9596 7340 9648
rect 7748 9596 7800 9648
rect 9864 9664 9916 9716
rect 10508 9664 10560 9716
rect 10784 9664 10836 9716
rect 12440 9664 12492 9716
rect 15752 9664 15804 9716
rect 16580 9664 16632 9716
rect 16948 9664 17000 9716
rect 19248 9664 19300 9716
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 3056 9435 3108 9444
rect 3056 9401 3090 9435
rect 3090 9401 3108 9435
rect 3056 9392 3108 9401
rect 10968 9528 11020 9580
rect 13912 9596 13964 9648
rect 15844 9596 15896 9648
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 13360 9528 13412 9580
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 9680 9460 9732 9512
rect 10232 9460 10284 9512
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13820 9460 13872 9512
rect 14556 9460 14608 9512
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 12256 9392 12308 9444
rect 8208 9324 8260 9376
rect 9864 9324 9916 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 10876 9324 10928 9376
rect 11612 9324 11664 9376
rect 11888 9324 11940 9376
rect 14004 9392 14056 9444
rect 17684 9392 17736 9444
rect 19340 9460 19392 9512
rect 20168 9460 20220 9512
rect 19800 9392 19852 9444
rect 12532 9324 12584 9376
rect 13360 9324 13412 9376
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 16580 9324 16632 9376
rect 17224 9324 17276 9376
rect 18788 9324 18840 9376
rect 19064 9324 19116 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 5172 9120 5224 9172
rect 6184 9120 6236 9172
rect 7380 9120 7432 9172
rect 10600 9120 10652 9172
rect 12808 9120 12860 9172
rect 17500 9120 17552 9172
rect 18880 9120 18932 9172
rect 19156 9120 19208 9172
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 3332 9052 3384 9104
rect 3976 9052 4028 9104
rect 4068 9052 4120 9104
rect 5540 9052 5592 9104
rect 6736 9052 6788 9104
rect 11612 9052 11664 9104
rect 18512 9052 18564 9104
rect 19524 9095 19576 9104
rect 19524 9061 19533 9095
rect 19533 9061 19567 9095
rect 19567 9061 19576 9095
rect 19524 9052 19576 9061
rect 2964 8984 3016 9036
rect 3056 8823 3108 8832
rect 3056 8789 3065 8823
rect 3065 8789 3099 8823
rect 3099 8789 3108 8823
rect 3056 8780 3108 8789
rect 4252 8780 4304 8832
rect 5632 8984 5684 9036
rect 6828 8984 6880 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 12992 9027 13044 9036
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5448 8916 5500 8968
rect 7104 8916 7156 8968
rect 7564 8848 7616 8900
rect 11704 8916 11756 8968
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 17592 8984 17644 9036
rect 13176 8916 13228 8968
rect 13820 8916 13872 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 19800 8959 19852 8968
rect 19800 8925 19809 8959
rect 19809 8925 19843 8959
rect 19843 8925 19852 8959
rect 19800 8916 19852 8925
rect 20996 8916 21048 8968
rect 14096 8848 14148 8900
rect 5724 8780 5776 8832
rect 6644 8780 6696 8832
rect 7196 8780 7248 8832
rect 11704 8780 11756 8832
rect 12624 8823 12676 8832
rect 12624 8789 12633 8823
rect 12633 8789 12667 8823
rect 12667 8789 12676 8823
rect 12624 8780 12676 8789
rect 18788 8780 18840 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 6828 8619 6880 8628
rect 5632 8576 5684 8585
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 9680 8576 9732 8628
rect 10232 8508 10284 8560
rect 10784 8508 10836 8560
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 17224 8508 17276 8560
rect 7564 8440 7616 8492
rect 7748 8440 7800 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 3148 8372 3200 8424
rect 3976 8372 4028 8424
rect 5448 8372 5500 8424
rect 5632 8372 5684 8424
rect 3240 8304 3292 8356
rect 2320 8279 2372 8288
rect 2320 8245 2329 8279
rect 2329 8245 2363 8279
rect 2363 8245 2372 8279
rect 2320 8236 2372 8245
rect 2596 8236 2648 8288
rect 4160 8236 4212 8288
rect 6828 8304 6880 8356
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 7932 8372 7984 8424
rect 10968 8372 11020 8424
rect 12348 8372 12400 8424
rect 12532 8372 12584 8424
rect 12716 8415 12768 8424
rect 12716 8381 12750 8415
rect 12750 8381 12768 8415
rect 12716 8372 12768 8381
rect 13728 8372 13780 8424
rect 8484 8304 8536 8356
rect 4712 8236 4764 8288
rect 11888 8304 11940 8356
rect 16672 8372 16724 8424
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17592 8440 17644 8492
rect 18972 8440 19024 8492
rect 19340 8372 19392 8424
rect 19800 8372 19852 8424
rect 10784 8236 10836 8288
rect 16580 8304 16632 8356
rect 18972 8304 19024 8356
rect 12900 8236 12952 8288
rect 13176 8236 13228 8288
rect 16212 8236 16264 8288
rect 16856 8236 16908 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 20628 8279 20680 8288
rect 20628 8245 20637 8279
rect 20637 8245 20671 8279
rect 20671 8245 20680 8279
rect 20628 8236 20680 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1768 8032 1820 8084
rect 4252 8032 4304 8084
rect 7104 8032 7156 8084
rect 7288 8032 7340 8084
rect 7748 8032 7800 8084
rect 9680 8032 9732 8084
rect 9956 8032 10008 8084
rect 12348 8075 12400 8084
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 2688 7964 2740 8016
rect 3148 7964 3200 8016
rect 2228 7896 2280 7948
rect 3056 7896 3108 7948
rect 8208 7964 8260 8016
rect 2596 7828 2648 7880
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 6000 7896 6052 7948
rect 8576 7964 8628 8016
rect 13268 7964 13320 8016
rect 14004 8007 14056 8016
rect 14004 7973 14013 8007
rect 14013 7973 14047 8007
rect 14047 7973 14056 8007
rect 14004 7964 14056 7973
rect 17408 8032 17460 8084
rect 17684 8032 17736 8084
rect 18420 8032 18472 8084
rect 20352 8032 20404 8084
rect 15844 7964 15896 8016
rect 15936 7964 15988 8016
rect 2964 7828 3016 7837
rect 6736 7828 6788 7880
rect 7564 7828 7616 7880
rect 8392 7896 8444 7948
rect 13728 7896 13780 7948
rect 17408 7939 17460 7948
rect 8668 7760 8720 7812
rect 2688 7692 2740 7744
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 6184 7692 6236 7744
rect 9772 7760 9824 7812
rect 9128 7692 9180 7744
rect 10048 7760 10100 7812
rect 11980 7692 12032 7744
rect 13176 7828 13228 7880
rect 12716 7760 12768 7812
rect 13912 7828 13964 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 18052 7896 18104 7948
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 20628 7828 20680 7880
rect 13360 7760 13412 7812
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 14280 7692 14332 7744
rect 17132 7692 17184 7744
rect 19616 7692 19668 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 8760 7488 8812 7540
rect 10876 7488 10928 7540
rect 11060 7488 11112 7540
rect 12256 7488 12308 7540
rect 12440 7488 12492 7540
rect 17592 7531 17644 7540
rect 8208 7420 8260 7472
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 18512 7420 18564 7472
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 3056 7352 3108 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 7196 7352 7248 7404
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 2320 7284 2372 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9680 7327 9732 7336
rect 9128 7284 9180 7293
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 12992 7352 13044 7404
rect 6000 7216 6052 7268
rect 6368 7216 6420 7268
rect 5816 7148 5868 7200
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 10048 7216 10100 7268
rect 9772 7148 9824 7200
rect 10600 7148 10652 7200
rect 10876 7148 10928 7200
rect 12348 7284 12400 7336
rect 13820 7284 13872 7336
rect 13912 7284 13964 7336
rect 13452 7216 13504 7268
rect 15292 7216 15344 7268
rect 16212 7327 16264 7336
rect 16212 7293 16221 7327
rect 16221 7293 16255 7327
rect 16255 7293 16264 7327
rect 16212 7284 16264 7293
rect 16488 7327 16540 7336
rect 16488 7293 16522 7327
rect 16522 7293 16540 7327
rect 19340 7327 19392 7336
rect 16488 7284 16540 7293
rect 19340 7293 19349 7327
rect 19349 7293 19383 7327
rect 19383 7293 19392 7327
rect 19340 7284 19392 7293
rect 19432 7284 19484 7336
rect 20628 7284 20680 7336
rect 20536 7216 20588 7268
rect 11152 7148 11204 7200
rect 12716 7148 12768 7200
rect 13728 7148 13780 7200
rect 15476 7148 15528 7200
rect 17960 7148 18012 7200
rect 19432 7148 19484 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 5816 6987 5868 6996
rect 5816 6953 5825 6987
rect 5825 6953 5859 6987
rect 5859 6953 5868 6987
rect 5816 6944 5868 6953
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 6644 6944 6696 6996
rect 8576 6944 8628 6996
rect 1308 6876 1360 6928
rect 6368 6876 6420 6928
rect 6920 6876 6972 6928
rect 8392 6876 8444 6928
rect 4068 6808 4120 6860
rect 6184 6808 6236 6860
rect 1952 6740 2004 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 2228 6672 2280 6724
rect 5908 6740 5960 6792
rect 7932 6808 7984 6860
rect 11612 6944 11664 6996
rect 12624 6944 12676 6996
rect 13636 6944 13688 6996
rect 12348 6876 12400 6928
rect 16212 6876 16264 6928
rect 16764 6876 16816 6928
rect 7472 6740 7524 6792
rect 16580 6808 16632 6860
rect 19340 6876 19392 6928
rect 19432 6851 19484 6860
rect 19432 6817 19466 6851
rect 19466 6817 19484 6851
rect 19432 6808 19484 6817
rect 6920 6672 6972 6724
rect 7564 6672 7616 6724
rect 13728 6740 13780 6792
rect 16948 6740 17000 6792
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 12440 6672 12492 6724
rect 13912 6672 13964 6724
rect 1860 6604 1912 6656
rect 7748 6604 7800 6656
rect 7932 6604 7984 6656
rect 10784 6604 10836 6656
rect 10968 6604 11020 6656
rect 13084 6604 13136 6656
rect 13268 6604 13320 6656
rect 16488 6604 16540 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 6000 6400 6052 6452
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 5540 6264 5592 6316
rect 6000 6264 6052 6316
rect 6920 6264 6972 6316
rect 7288 6400 7340 6452
rect 7472 6400 7524 6452
rect 8484 6443 8536 6452
rect 8484 6409 8493 6443
rect 8493 6409 8527 6443
rect 8527 6409 8536 6443
rect 8484 6400 8536 6409
rect 9036 6400 9088 6452
rect 12440 6400 12492 6452
rect 12532 6400 12584 6452
rect 18512 6400 18564 6452
rect 11888 6332 11940 6384
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 11336 6264 11388 6316
rect 11612 6264 11664 6316
rect 17960 6332 18012 6384
rect 19432 6332 19484 6384
rect 13176 6264 13228 6316
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 3792 6196 3844 6248
rect 7196 6196 7248 6248
rect 8668 6196 8720 6248
rect 9220 6196 9272 6248
rect 2504 6128 2556 6180
rect 6736 6128 6788 6180
rect 9864 6196 9916 6248
rect 13268 6196 13320 6248
rect 15384 6264 15436 6316
rect 16580 6264 16632 6316
rect 17316 6264 17368 6316
rect 17868 6264 17920 6316
rect 19616 6307 19668 6316
rect 19616 6273 19625 6307
rect 19625 6273 19659 6307
rect 19659 6273 19668 6307
rect 19616 6264 19668 6273
rect 19800 6264 19852 6316
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 17040 6239 17092 6248
rect 17040 6205 17049 6239
rect 17049 6205 17083 6239
rect 17083 6205 17092 6239
rect 17040 6196 17092 6205
rect 18696 6196 18748 6248
rect 20536 6196 20588 6248
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 4160 6060 4212 6112
rect 5264 6060 5316 6112
rect 9128 6060 9180 6112
rect 9220 6060 9272 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 10784 6103 10836 6112
rect 9864 6060 9916 6069
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 13268 6060 13320 6112
rect 13544 6128 13596 6180
rect 13728 6128 13780 6180
rect 18880 6128 18932 6180
rect 18972 6128 19024 6180
rect 19340 6128 19392 6180
rect 15108 6103 15160 6112
rect 15108 6069 15117 6103
rect 15117 6069 15151 6103
rect 15151 6069 15160 6103
rect 15108 6060 15160 6069
rect 16212 6060 16264 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 18420 6103 18472 6112
rect 18420 6069 18429 6103
rect 18429 6069 18463 6103
rect 18463 6069 18472 6103
rect 18420 6060 18472 6069
rect 18696 6060 18748 6112
rect 19248 6060 19300 6112
rect 19892 6060 19944 6112
rect 20536 6103 20588 6112
rect 20536 6069 20545 6103
rect 20545 6069 20579 6103
rect 20579 6069 20588 6103
rect 20536 6060 20588 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 3976 5856 4028 5908
rect 4068 5788 4120 5840
rect 6000 5856 6052 5908
rect 7196 5856 7248 5908
rect 7748 5856 7800 5908
rect 8208 5856 8260 5908
rect 10876 5856 10928 5908
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 2504 5584 2556 5636
rect 3792 5652 3844 5704
rect 5448 5720 5500 5772
rect 6000 5763 6052 5772
rect 6000 5729 6034 5763
rect 6034 5729 6052 5763
rect 6000 5720 6052 5729
rect 5632 5652 5684 5704
rect 3884 5516 3936 5568
rect 5540 5516 5592 5568
rect 5908 5516 5960 5568
rect 9220 5788 9272 5840
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 8484 5720 8536 5772
rect 10140 5720 10192 5772
rect 11612 5788 11664 5840
rect 11888 5856 11940 5908
rect 14280 5856 14332 5908
rect 14372 5856 14424 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 15108 5788 15160 5840
rect 11336 5720 11388 5772
rect 17132 5856 17184 5908
rect 18052 5856 18104 5908
rect 20536 5856 20588 5908
rect 7196 5652 7248 5704
rect 10324 5652 10376 5704
rect 10968 5652 11020 5704
rect 12808 5652 12860 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 9772 5516 9824 5568
rect 17132 5720 17184 5772
rect 17868 5720 17920 5772
rect 12440 5516 12492 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 16120 5516 16172 5568
rect 16672 5516 16724 5568
rect 18972 5652 19024 5704
rect 19800 5652 19852 5704
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2688 5312 2740 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 11152 5312 11204 5364
rect 2228 5244 2280 5296
rect 8484 5244 8536 5296
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2504 5176 2556 5228
rect 2688 5176 2740 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 7564 5176 7616 5228
rect 16672 5176 16724 5228
rect 1584 5108 1636 5160
rect 3332 5108 3384 5160
rect 7288 5108 7340 5160
rect 10968 5108 11020 5160
rect 11612 5108 11664 5160
rect 12808 5151 12860 5160
rect 12808 5117 12842 5151
rect 12842 5117 12860 5151
rect 6920 5040 6972 5092
rect 12808 5108 12860 5117
rect 13544 5108 13596 5160
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 4160 4972 4212 5024
rect 7472 4972 7524 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 13728 5040 13780 5092
rect 13636 4972 13688 5024
rect 18972 5040 19024 5092
rect 15936 4972 15988 5024
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 20260 4972 20312 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2596 4768 2648 4820
rect 1952 4632 2004 4684
rect 1032 4564 1084 4616
rect 10140 4768 10192 4820
rect 10784 4768 10836 4820
rect 11520 4768 11572 4820
rect 12900 4768 12952 4820
rect 15200 4768 15252 4820
rect 17316 4768 17368 4820
rect 6184 4700 6236 4752
rect 12992 4700 13044 4752
rect 13268 4700 13320 4752
rect 17040 4700 17092 4752
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 8300 4675 8352 4684
rect 5448 4632 5500 4641
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 2688 4496 2740 4548
rect 5816 4564 5868 4616
rect 6184 4564 6236 4616
rect 7564 4564 7616 4616
rect 2964 4496 3016 4548
rect 3332 4496 3384 4548
rect 9680 4632 9732 4684
rect 10784 4632 10836 4684
rect 10968 4632 11020 4684
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 10600 4564 10652 4616
rect 16304 4632 16356 4684
rect 20168 4632 20220 4684
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 16672 4607 16724 4616
rect 15936 4564 15988 4573
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 9680 4496 9732 4548
rect 4160 4428 4212 4480
rect 8760 4428 8812 4480
rect 9036 4428 9088 4480
rect 13636 4428 13688 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 18512 4428 18564 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3056 4224 3108 4276
rect 7564 4267 7616 4276
rect 3976 4156 4028 4208
rect 4068 4156 4120 4208
rect 5908 4156 5960 4208
rect 1584 4020 1636 4072
rect 2688 4020 2740 4072
rect 3332 3952 3384 4004
rect 5356 4088 5408 4140
rect 6736 4156 6788 4208
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 8300 4224 8352 4276
rect 10876 4224 10928 4276
rect 18512 4224 18564 4276
rect 8208 4131 8260 4140
rect 4988 4020 5040 4072
rect 6644 4020 6696 4072
rect 2504 3884 2556 3936
rect 3700 3884 3752 3936
rect 5816 3952 5868 4004
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 9036 4131 9088 4140
rect 9036 4097 9045 4131
rect 9045 4097 9079 4131
rect 9079 4097 9088 4131
rect 9036 4088 9088 4097
rect 9312 4156 9364 4208
rect 9680 4156 9732 4208
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9128 3952 9180 4004
rect 10416 3952 10468 4004
rect 15476 4020 15528 4072
rect 18880 4088 18932 4140
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 15936 4063 15988 4072
rect 15936 4029 15970 4063
rect 15970 4029 15988 4063
rect 15936 4020 15988 4029
rect 18972 4063 19024 4072
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 19892 4063 19944 4072
rect 19892 4029 19901 4063
rect 19901 4029 19935 4063
rect 19935 4029 19944 4063
rect 19892 4020 19944 4029
rect 20628 4020 20680 4072
rect 20720 4020 20772 4072
rect 17408 3952 17460 4004
rect 5264 3884 5316 3936
rect 5632 3884 5684 3936
rect 6000 3884 6052 3936
rect 8760 3884 8812 3936
rect 10324 3884 10376 3936
rect 14556 3884 14608 3936
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 16672 3884 16724 3936
rect 17040 3927 17092 3936
rect 17040 3893 17049 3927
rect 17049 3893 17083 3927
rect 17083 3893 17092 3927
rect 17040 3884 17092 3893
rect 18696 3884 18748 3936
rect 18880 3884 18932 3936
rect 19708 3884 19760 3936
rect 19800 3884 19852 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 204 3680 256 3732
rect 2964 3680 3016 3732
rect 6460 3680 6512 3732
rect 9864 3680 9916 3732
rect 9956 3680 10008 3732
rect 15108 3680 15160 3732
rect 15384 3680 15436 3732
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 4160 3612 4212 3664
rect 5632 3612 5684 3664
rect 6920 3612 6972 3664
rect 2780 3340 2832 3392
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 7472 3612 7524 3664
rect 8208 3612 8260 3664
rect 8484 3612 8536 3664
rect 6000 3544 6052 3553
rect 7288 3544 7340 3596
rect 10232 3544 10284 3596
rect 10416 3544 10468 3596
rect 10784 3544 10836 3596
rect 12992 3612 13044 3664
rect 14556 3612 14608 3664
rect 12440 3587 12492 3596
rect 12440 3553 12449 3587
rect 12449 3553 12483 3587
rect 12483 3553 12492 3587
rect 12440 3544 12492 3553
rect 13636 3587 13688 3596
rect 13636 3553 13645 3587
rect 13645 3553 13679 3587
rect 13679 3553 13688 3587
rect 13636 3544 13688 3553
rect 15200 3544 15252 3596
rect 18604 3587 18656 3596
rect 18604 3553 18613 3587
rect 18613 3553 18647 3587
rect 18647 3553 18656 3587
rect 18604 3544 18656 3553
rect 19156 3544 19208 3596
rect 19984 3544 20036 3596
rect 3792 3476 3844 3528
rect 5356 3476 5408 3528
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 6552 3476 6604 3528
rect 8760 3476 8812 3528
rect 9956 3476 10008 3528
rect 10048 3476 10100 3528
rect 10324 3476 10376 3528
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 13728 3476 13780 3528
rect 15476 3476 15528 3528
rect 17040 3476 17092 3528
rect 3700 3408 3752 3460
rect 8852 3408 8904 3460
rect 11060 3408 11112 3460
rect 21180 3408 21232 3460
rect 4252 3340 4304 3392
rect 4712 3340 4764 3392
rect 9680 3340 9732 3392
rect 10232 3383 10284 3392
rect 10232 3349 10241 3383
rect 10241 3349 10275 3383
rect 10275 3349 10284 3383
rect 10232 3340 10284 3349
rect 15384 3340 15436 3392
rect 18512 3340 18564 3392
rect 19156 3340 19208 3392
rect 19524 3340 19576 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2688 3136 2740 3188
rect 3700 3136 3752 3188
rect 5356 3179 5408 3188
rect 3424 3068 3476 3120
rect 3792 3068 3844 3120
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 8576 3136 8628 3188
rect 7380 3068 7432 3120
rect 10140 3068 10192 3120
rect 11060 3136 11112 3188
rect 15200 3136 15252 3188
rect 7288 3000 7340 3052
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 1492 2864 1544 2916
rect 3516 2864 3568 2916
rect 3976 2975 4028 2984
rect 3976 2941 3985 2975
rect 3985 2941 4019 2975
rect 4019 2941 4028 2975
rect 3976 2932 4028 2941
rect 6552 2932 6604 2984
rect 9680 3000 9732 3052
rect 10324 3000 10376 3052
rect 10876 3000 10928 3052
rect 11428 3068 11480 3120
rect 15016 3068 15068 3120
rect 9312 2932 9364 2984
rect 6000 2864 6052 2916
rect 2412 2796 2464 2848
rect 2780 2796 2832 2848
rect 2964 2796 3016 2848
rect 11428 2932 11480 2984
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 13084 2932 13136 2941
rect 13912 2932 13964 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 18696 3068 18748 3120
rect 18604 3000 18656 3052
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 19248 2932 19300 2984
rect 21640 2932 21692 2984
rect 12532 2864 12584 2916
rect 14464 2864 14516 2916
rect 17408 2864 17460 2916
rect 18328 2907 18380 2916
rect 18328 2873 18337 2907
rect 18337 2873 18371 2907
rect 18371 2873 18380 2907
rect 18328 2864 18380 2873
rect 18880 2864 18932 2916
rect 19892 2864 19944 2916
rect 22560 2864 22612 2916
rect 9588 2839 9640 2848
rect 9588 2805 9597 2839
rect 9597 2805 9631 2839
rect 9631 2805 9640 2839
rect 9588 2796 9640 2805
rect 10140 2796 10192 2848
rect 13176 2796 13228 2848
rect 15384 2796 15436 2848
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 16304 2796 16356 2805
rect 18972 2796 19024 2848
rect 19708 2796 19760 2848
rect 22100 2796 22152 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 3424 2524 3476 2576
rect 4252 2592 4304 2644
rect 4712 2592 4764 2644
rect 6552 2635 6604 2644
rect 6552 2601 6561 2635
rect 6561 2601 6595 2635
rect 6595 2601 6604 2635
rect 6552 2592 6604 2601
rect 10048 2592 10100 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 1584 2456 1636 2508
rect 3976 2456 4028 2508
rect 8576 2524 8628 2576
rect 10140 2567 10192 2576
rect 10140 2533 10149 2567
rect 10149 2533 10183 2567
rect 10183 2533 10192 2567
rect 10140 2524 10192 2533
rect 10692 2524 10744 2576
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 12532 2456 12584 2508
rect 12992 2456 13044 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 3516 2320 3568 2372
rect 9588 2388 9640 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 14464 2456 14516 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16120 2499 16172 2508
rect 16120 2465 16129 2499
rect 16129 2465 16163 2499
rect 16163 2465 16172 2499
rect 16120 2456 16172 2465
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 17960 2320 18012 2372
rect 572 2252 624 2304
rect 4988 2252 5040 2304
rect 5540 2252 5592 2304
rect 8944 2252 8996 2304
rect 12716 2252 12768 2304
rect 13544 2252 13596 2304
rect 14004 2252 14056 2304
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 14924 2252 14976 2304
rect 15844 2252 15896 2304
rect 16672 2252 16724 2304
rect 17132 2252 17184 2304
rect 17684 2252 17736 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 6000 1368 6052 1420
rect 8760 1368 8812 1420
rect 11336 1232 11388 1284
rect 12164 1232 12216 1284
rect 4068 1028 4120 1080
rect 5724 1028 5776 1080
<< metal2 >>
rect 4250 22536 4306 22545
rect 4250 22471 4306 22480
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2778 21176 2834 21185
rect 2778 21111 2834 21120
rect 2792 20058 2820 21111
rect 2870 20224 2926 20233
rect 2870 20159 2926 20168
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2042 19816 2098 19825
rect 2042 19751 2098 19760
rect 2056 19514 2084 19751
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 2778 19272 2834 19281
rect 1872 18154 1900 19246
rect 2778 19207 2834 19216
rect 2792 18970 2820 19207
rect 2884 19174 2912 20159
rect 2976 19786 3004 21519
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 3068 18970 3096 22063
rect 4066 20632 4122 20641
rect 4066 20567 4122 20576
rect 4080 19514 4108 20567
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 1964 18873 1992 18906
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 1952 18352 2004 18358
rect 1950 18320 1952 18329
rect 2004 18320 2006 18329
rect 1950 18255 2006 18264
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1582 17912 1638 17921
rect 1582 17847 1584 17856
rect 1636 17847 1638 17856
rect 1584 17818 1636 17824
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2056 17134 2084 17478
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 15065 1716 16934
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 1780 15978 1808 16594
rect 1950 16552 2006 16561
rect 1950 16487 1952 16496
rect 2004 16487 2006 16496
rect 1952 16458 2004 16464
rect 2332 16114 2360 16594
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 1950 16008 2006 16017
rect 1768 15972 1820 15978
rect 1950 15943 2006 15952
rect 1768 15914 1820 15920
rect 1964 15706 1992 15943
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1950 15600 2006 15609
rect 1950 15535 2006 15544
rect 1964 15162 1992 15535
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 1688 13938 1716 14418
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1964 14113 1992 14214
rect 1950 14104 2006 14113
rect 2148 14074 2176 14418
rect 1950 14039 2006 14048
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2240 13530 2268 13670
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 12986 2452 13262
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2516 12322 2544 18770
rect 3160 18766 3188 19246
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3160 18222 3188 18702
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 2608 17882 2636 18022
rect 2976 17882 3004 18022
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2870 17368 2926 17377
rect 3068 17338 3096 18022
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 2870 17303 2926 17312
rect 3056 17332 3108 17338
rect 2778 16960 2834 16969
rect 2778 16895 2834 16904
rect 2792 16794 2820 16895
rect 2884 16794 2912 17303
rect 3056 17274 3108 17280
rect 3344 16794 3372 17682
rect 3620 17678 3648 19178
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4172 18222 4200 19110
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 17814 4200 18158
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2700 14822 2728 15574
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2608 13870 2636 14214
rect 2700 13938 2728 14758
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2778 13696 2834 13705
rect 2608 12442 2636 13670
rect 2778 13631 2834 13640
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2424 12294 2544 12322
rect 2596 12300 2648 12306
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 1964 10674 1992 11154
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 9586 1992 10066
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1780 8090 1808 9454
rect 2424 8401 2452 12294
rect 2596 12242 2648 12248
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11354 2544 12174
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2608 10810 2636 12242
rect 2792 11082 2820 13631
rect 2884 13462 2912 16594
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 14414 3280 15302
rect 3330 14648 3386 14657
rect 3330 14583 3386 14592
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3068 14074 3096 14350
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3344 14006 3372 14583
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2964 13320 3016 13326
rect 2870 13288 2926 13297
rect 2964 13262 3016 13268
rect 2870 13223 2926 13232
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 8650 2820 10474
rect 2884 10266 2912 13223
rect 2976 12238 3004 13262
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3068 12170 3096 12786
rect 3436 12782 3464 17614
rect 3620 17202 3648 17614
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11694 3096 12106
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2976 10146 3004 11222
rect 3068 11150 3096 11630
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10674 3096 11086
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2700 8622 2820 8650
rect 2884 10118 3004 10146
rect 2410 8392 2466 8401
rect 2410 8327 2466 8336
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2240 7546 2268 7890
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2332 7342 2360 8230
rect 2608 7886 2636 8230
rect 2700 8022 2728 8622
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 7410 2728 7686
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2042 7168 2098 7177
rect 2042 7103 2098 7112
rect 1308 6928 1360 6934
rect 1308 6870 1360 6876
rect 1320 6225 1348 6870
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5166 1624 6054
rect 1872 5234 1900 6598
rect 1964 6254 1992 6734
rect 2056 6322 2084 7103
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6322 2268 6666
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 2240 5302 2268 6258
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2516 5642 2544 6122
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2516 5234 2544 5578
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1032 4616 1084 4622
rect 1032 4558 1084 4564
rect 204 3732 256 3738
rect 204 3674 256 3680
rect 216 800 244 3674
rect 572 2304 624 2310
rect 572 2246 624 2252
rect 584 800 612 2246
rect 1044 800 1072 4558
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 2990 1624 4014
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1492 2916 1544 2922
rect 1492 2858 1544 2864
rect 1504 800 1532 2858
rect 1596 2514 1624 2926
rect 1964 2825 1992 4626
rect 2516 3942 2544 5170
rect 2608 4826 2636 5714
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5370 2728 5646
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2700 4554 2728 5170
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2700 4078 2728 4490
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2700 3194 2728 4014
rect 2792 3505 2820 8366
rect 2884 7886 2912 10118
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8945 3004 8978
rect 2962 8936 3018 8945
rect 2962 8871 3018 8880
rect 2976 8498 3004 8871
rect 3068 8838 3096 9386
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 7886 3004 8434
rect 3068 7954 3096 8774
rect 3160 8430 3188 12718
rect 3528 11286 3556 17070
rect 4264 16998 4292 22471
rect 5722 22000 5778 22800
rect 17130 22000 17186 22800
rect 17866 22536 17922 22545
rect 17866 22471 17922 22480
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 17082 4752 18702
rect 5000 18086 5028 18770
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17882 5028 18022
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4816 17338 4844 17614
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4724 17054 4844 17082
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15162 4292 15302
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 15156 4304 15162
rect 4172 15116 4252 15144
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3804 13258 3832 14826
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 11830 3740 12174
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 8922 3280 11018
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 9110 3372 9454
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3252 8894 3372 8922
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 2854 2820 3334
rect 2412 2848 2464 2854
rect 1950 2816 2006 2825
rect 2412 2790 2464 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1950 2751 2006 2760
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1964 800 1992 2751
rect 2424 800 2452 2790
rect 2884 1601 2912 7822
rect 3068 7410 3096 7890
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 3738 3004 4490
rect 3068 4282 3096 6734
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2964 2848 3016 2854
rect 2962 2816 2964 2825
rect 3016 2816 3018 2825
rect 2962 2751 3018 2760
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3068 1442 3096 4218
rect 3160 2553 3188 7958
rect 3252 7410 3280 8298
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3344 7290 3372 8894
rect 3252 7262 3372 7290
rect 3146 2544 3202 2553
rect 3146 2479 3202 2488
rect 2884 1414 3096 1442
rect 2884 800 2912 1414
rect 3252 1057 3280 7262
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3344 4554 3372 5102
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3238 1048 3294 1057
rect 3238 983 3294 992
rect 3344 800 3372 3946
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3436 2582 3464 3062
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3528 2650 3556 2858
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3528 2378 3556 2586
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 3620 2009 3648 10406
rect 3804 10062 3832 10610
rect 3896 10538 3924 14214
rect 4066 12744 4122 12753
rect 4066 12679 4068 12688
rect 4120 12679 4122 12688
rect 4068 12650 4120 12656
rect 4172 11898 4200 15116
rect 4252 15098 4304 15104
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4264 11898 4292 13670
rect 4356 13530 4384 13670
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4724 12306 4752 16934
rect 4816 16658 4844 17054
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 15570 4844 16594
rect 4908 16182 4936 16934
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4816 15366 4844 15506
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 14482 4844 15302
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4066 11792 4122 11801
rect 4816 11762 4844 12038
rect 4066 11727 4122 11736
rect 4804 11756 4856 11762
rect 4080 11626 4108 11727
rect 4804 11698 4856 11704
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4066 10840 4122 10849
rect 4066 10775 4068 10784
rect 4120 10775 4122 10784
rect 4068 10746 4120 10752
rect 4172 10606 4200 10950
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3792 10056 3844 10062
rect 3988 10033 4016 10474
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 10198 4108 10367
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4068 10056 4120 10062
rect 3792 9998 3844 10004
rect 3974 10024 4030 10033
rect 4068 9998 4120 10004
rect 3974 9959 4030 9968
rect 4080 9602 4108 9998
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 3988 9574 4108 9602
rect 3988 9110 4016 9574
rect 4068 9512 4120 9518
rect 4066 9480 4068 9489
rect 4120 9480 4122 9489
rect 4066 9415 4122 9424
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3976 9104 4028 9110
rect 4068 9104 4120 9110
rect 3976 9046 4028 9052
rect 4066 9072 4068 9081
rect 4120 9072 4122 9081
rect 3988 8430 4016 9046
rect 4066 9007 4122 9016
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4172 8294 4200 9318
rect 4712 8968 4764 8974
rect 4710 8936 4712 8945
rect 4764 8936 4766 8945
rect 4710 8871 4766 8880
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4264 8090 4292 8774
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 8129 4752 8230
rect 4710 8120 4766 8129
rect 4252 8084 4304 8090
rect 4710 8055 4766 8064
rect 4252 8026 4304 8032
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 6769 4108 6802
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3804 5710 3832 6190
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5817 4016 5850
rect 4080 5846 4108 6054
rect 4068 5840 4120 5846
rect 3974 5808 4030 5817
rect 4068 5782 4120 5788
rect 3974 5743 4030 5752
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3804 4026 3832 5646
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5234 3924 5510
rect 3974 5264 4030 5273
rect 3884 5228 3936 5234
rect 4080 5234 4108 5782
rect 3974 5199 4030 5208
rect 4068 5228 4120 5234
rect 3884 5170 3936 5176
rect 3988 4214 4016 5199
rect 4068 5170 4120 5176
rect 4172 5030 4200 6054
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4080 4214 4108 4247
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 3804 3998 4016 4026
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3466 3740 3878
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3606 2000 3662 2009
rect 3606 1935 3662 1944
rect 3712 800 3740 3130
rect 3804 3126 3832 3470
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3988 2990 4016 3998
rect 4172 3670 4200 4422
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4816 3482 4844 11494
rect 4172 3454 4844 3482
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 2514 4016 2926
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4068 1080 4120 1086
rect 4068 1022 4120 1028
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4080 649 4108 1022
rect 4172 800 4200 3454
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4264 2650 4292 3334
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4724 2650 4752 3334
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4908 1986 4936 16118
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5000 12986 5028 13262
rect 5092 13190 5120 19246
rect 5184 15910 5212 19790
rect 5736 19174 5764 22000
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5644 17814 5672 18566
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16250 5304 16934
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5368 16114 5396 16594
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5368 15706 5396 16050
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5092 12782 5120 13126
rect 5276 12850 5304 15642
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5368 14074 5396 14418
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 10810 5028 11766
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5000 2310 5028 4014
rect 5092 2961 5120 9998
rect 5184 9178 5212 12242
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5276 6118 5304 12786
rect 5460 11286 5488 15914
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 11898 5580 13330
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12238 5672 12786
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5920 12306 5948 12378
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5644 11762 5672 12174
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 10538 5488 11086
rect 5644 10810 5672 11698
rect 5828 11694 5856 12038
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 10266 5488 10474
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5736 9654 5764 11154
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5354 9480 5410 9489
rect 5354 9415 5410 9424
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5368 4842 5396 9415
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8430 5488 8910
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5552 6322 5580 9046
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8634 5672 8978
rect 5724 8832 5776 8838
rect 5920 8820 5948 12242
rect 5776 8792 5948 8820
rect 5724 8774 5776 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5644 7750 5672 8366
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5184 4814 5396 4842
rect 5078 2952 5134 2961
rect 5078 2887 5134 2896
rect 5184 2836 5212 4814
rect 5460 4690 5488 5714
rect 5644 5710 5672 7686
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5368 4146 5396 4626
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5264 3936 5316 3942
rect 5552 3924 5580 5510
rect 5316 3896 5580 3924
rect 5632 3936 5684 3942
rect 5264 3878 5316 3884
rect 5632 3878 5684 3884
rect 5644 3670 5672 3878
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5368 3194 5396 3470
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5092 2808 5212 2836
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4632 1958 4936 1986
rect 4632 800 4660 1958
rect 5092 800 5120 2808
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 800 5580 2246
rect 5736 1086 5764 8774
rect 6012 7954 6040 18090
rect 6104 14550 6132 18566
rect 7024 18426 7052 19246
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6472 16454 6500 17138
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 16114 6500 16390
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6090 14104 6146 14113
rect 6090 14039 6146 14048
rect 6104 13870 6132 14039
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6196 12220 6224 12786
rect 6288 12442 6316 13738
rect 6656 12646 6684 16934
rect 6748 16250 6776 17546
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15638 6868 15846
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6748 14278 6776 15574
rect 6932 14618 6960 15982
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13938 6776 14214
rect 6840 14074 6868 14350
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6932 13546 6960 14010
rect 6840 13518 6960 13546
rect 6840 13394 6868 13518
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6276 12232 6328 12238
rect 6196 12192 6276 12220
rect 6276 12174 6328 12180
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6288 9654 6316 12174
rect 6380 11762 6408 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 10266 6408 11154
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6472 10810 6500 11086
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6564 10130 6592 11086
rect 6656 10130 6684 12582
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11150 6776 11494
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6564 9926 6592 10066
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 7002 5856 7142
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 5574 5948 6734
rect 6012 6458 6040 7210
rect 6196 7002 6224 7686
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6196 6866 6224 6938
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5914 6040 6258
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6012 5778 6040 5850
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 6182 4856 6238 4865
rect 6182 4791 6238 4800
rect 6196 4758 6224 4791
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 5828 4010 5856 4558
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5920 3924 5948 4150
rect 6196 4146 6224 4558
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6000 3936 6052 3942
rect 5920 3896 6000 3924
rect 6000 3878 6052 3884
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6012 2922 6040 3538
rect 6196 3534 6224 4082
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 5724 1080 5776 1086
rect 5724 1022 5776 1028
rect 6012 800 6040 1362
rect 4066 640 4122 649
rect 4066 575 4122 584
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6288 241 6316 9590
rect 6380 9586 6408 9862
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8276 6684 8774
rect 6748 8344 6776 9046
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8634 6868 8978
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6828 8356 6880 8362
rect 6748 8316 6828 8344
rect 6828 8298 6880 8304
rect 6656 8248 6776 8276
rect 6748 7886 6776 8248
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6380 6934 6408 7210
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6656 4078 6684 6938
rect 6748 6186 6776 7822
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6748 4214 6776 6122
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6472 800 6500 3674
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 2990 6592 3470
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6564 2650 6592 2926
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6840 800 6868 8298
rect 6932 6934 6960 12242
rect 7024 12102 7052 17002
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7116 13870 7144 15506
rect 7208 14074 7236 19858
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7760 19242 7788 19314
rect 8484 19304 8536 19310
rect 8220 19264 8484 19292
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7300 17610 7328 18770
rect 7392 18222 7420 19110
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7300 17202 7328 17546
rect 7576 17338 7604 19110
rect 7668 18290 7696 19178
rect 7760 18970 7788 19178
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18970 8248 19264
rect 8484 19246 8536 19252
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8220 18630 8248 18906
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8220 18290 8248 18566
rect 8404 18358 8432 18566
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17338 8064 17682
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8220 16726 8248 18226
rect 8760 18148 8812 18154
rect 8760 18090 8812 18096
rect 8772 17202 8800 18090
rect 9692 17882 9720 18770
rect 9876 18222 9904 19110
rect 10152 18970 10180 19246
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9784 17678 9812 18022
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8208 16720 8260 16726
rect 8208 16662 8260 16668
rect 8220 16046 8248 16662
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14958 7328 15302
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14346 7328 14894
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 12986 7144 13806
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 11234 7052 11630
rect 7116 11354 7144 12718
rect 7208 12442 7236 13670
rect 7300 13530 7328 13670
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7392 13190 7420 15846
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15366 8248 15982
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 15162 8248 15302
rect 8404 15162 8432 17002
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 15706 8524 16934
rect 8772 16794 8800 17138
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 16250 9628 16594
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7024 11218 7144 11234
rect 7024 11212 7156 11218
rect 7024 11206 7104 11212
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6322 6960 6666
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6932 3670 6960 5034
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7024 2938 7052 11206
rect 7104 11154 7156 11160
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7116 10282 7144 10950
rect 7208 10470 7236 11494
rect 7300 11082 7328 12038
rect 7484 11694 7512 12174
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10674 7328 11018
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7116 10254 7236 10282
rect 7392 10266 7420 10406
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8090 7144 8910
rect 7208 8838 7236 10254
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7300 9654 7328 9998
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7288 8424 7340 8430
rect 7392 8412 7420 9114
rect 7340 8384 7420 8412
rect 7288 8366 7340 8372
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7208 6254 7236 7346
rect 7300 6458 7328 8026
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7208 5710 7236 5850
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7300 5166 7328 6394
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 3602 7328 5102
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7300 3058 7328 3538
rect 7392 3126 7420 8384
rect 7484 6798 7512 11222
rect 7576 11014 7604 14826
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7760 13308 7788 14486
rect 8312 14006 8340 14758
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7840 13320 7892 13326
rect 7760 13280 7840 13308
rect 7892 13280 7972 13308
rect 7840 13262 7892 13268
rect 7944 12850 7972 13280
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12238 8248 12786
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10130 7604 10610
rect 7668 10248 7696 12174
rect 8220 11762 8248 12174
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 11218 7788 11494
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7668 10220 7880 10248
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9586 7604 10066
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 8906 7604 9522
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7576 7886 7604 8434
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7484 5030 7512 6394
rect 7576 5234 7604 6666
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7668 4978 7696 9658
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7760 8498 7788 9590
rect 7852 9489 7880 10220
rect 8220 9518 8248 11290
rect 8312 9722 8340 13126
rect 8404 12986 8432 14418
rect 8496 14074 8524 14758
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8390 12336 8446 12345
rect 8588 12306 8616 15302
rect 8956 14074 8984 15506
rect 9600 15502 9628 16186
rect 9588 15496 9640 15502
rect 9876 15484 9904 17682
rect 9968 16182 9996 18634
rect 10336 18426 10364 18838
rect 10796 18766 10824 19246
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18834 11560 19110
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10060 18086 10088 18226
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10060 17610 10088 18022
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9968 15638 9996 16118
rect 10152 15706 10180 17478
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9876 15456 10088 15484
rect 9588 15438 9640 15444
rect 9600 15026 9628 15438
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9586 14104 9642 14113
rect 8944 14068 8996 14074
rect 9586 14039 9588 14048
rect 8944 14010 8996 14016
rect 9640 14039 9642 14048
rect 9956 14068 10008 14074
rect 9588 14010 9640 14016
rect 9956 14010 10008 14016
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8956 12850 8984 13670
rect 9232 13394 9260 13874
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9416 13682 9444 13738
rect 9680 13728 9732 13734
rect 9416 13676 9680 13682
rect 9416 13670 9732 13676
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8390 12271 8446 12280
rect 8576 12300 8628 12306
rect 8404 11150 8432 12271
rect 8576 12242 8628 12248
rect 8680 11665 8708 12310
rect 8772 11898 8800 12582
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8864 11898 8892 12106
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8666 11656 8722 11665
rect 8666 11591 8722 11600
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9512 8260 9518
rect 7838 9480 7894 9489
rect 8208 9454 8260 9460
rect 7838 9415 7894 9424
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7930 8528 7986 8537
rect 7748 8492 7800 8498
rect 7930 8463 7986 8472
rect 7748 8434 7800 8440
rect 7760 8090 7788 8434
rect 7944 8430 7972 8463
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8220 8022 8248 9318
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8484 8356 8536 8362
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8404 7954 8432 8327
rect 8484 8298 8536 8304
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7944 6662 7972 6802
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7760 5914 7788 6598
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5914 8248 7414
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5370 7880 5714
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7484 3670 7512 4966
rect 7668 4950 7788 4978
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4282 7604 4558
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7024 2910 7328 2938
rect 7300 800 7328 2910
rect 7760 800 7788 4950
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4282 8340 4626
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3670 8248 4082
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8404 3516 8432 6870
rect 8496 6458 8524 8298
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 7002 8616 7958
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8680 7546 8708 7754
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8772 7449 8800 7482
rect 8758 7440 8814 7449
rect 8758 7375 8814 7384
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8496 5778 8524 6394
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8496 3670 8524 5238
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8220 3488 8432 3516
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 800 8248 3488
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8588 2582 8616 3130
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8680 800 8708 6190
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 3942 8800 4422
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8864 3890 8892 11290
rect 8956 11014 8984 11494
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7342 9168 7686
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6458 9076 7142
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9232 6254 9260 13330
rect 9324 13326 9352 13670
rect 9416 13654 9720 13670
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 11354 9352 13262
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9600 11286 9628 11766
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9692 10266 9720 13466
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11762 9812 12242
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9876 10713 9904 13398
rect 9862 10704 9918 10713
rect 9862 10639 9918 10648
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9310 8936 9366 8945
rect 9310 8871 9366 8880
rect 9324 7410 9352 8871
rect 9692 8634 9720 9454
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9692 7342 9720 8026
rect 9784 7936 9812 10066
rect 9876 9722 9904 10542
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9864 9376 9916 9382
rect 9862 9344 9864 9353
rect 9916 9344 9918 9353
rect 9862 9279 9918 9288
rect 9968 8090 9996 14010
rect 10060 9636 10088 15456
rect 10152 15366 10180 15642
rect 10244 15502 10272 15914
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 14074 10180 14826
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10244 13938 10272 15438
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 10266 10272 11494
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10152 9994 10180 10202
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10060 9608 10180 9636
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9784 7908 9904 7936
rect 9770 7848 9826 7857
rect 9770 7783 9772 7792
rect 9824 7783 9826 7792
rect 9772 7754 9824 7760
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9770 7304 9826 7313
rect 9770 7239 9826 7248
rect 9784 7206 9812 7239
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9876 6440 9904 7908
rect 9692 6412 9904 6440
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 6112 9180 6118
rect 9126 6080 9128 6089
rect 9220 6112 9272 6118
rect 9180 6080 9182 6089
rect 9220 6054 9272 6060
rect 9126 6015 9182 6024
rect 9232 5846 9260 6054
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 4078 8984 4558
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9048 4146 9076 4422
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8864 3862 8984 3890
rect 8850 3632 8906 3641
rect 8850 3567 8906 3576
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 1426 8800 3470
rect 8864 3466 8892 3567
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8956 2310 8984 3862
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 9140 800 9168 3946
rect 9232 1306 9260 5782
rect 9692 4690 9720 6412
rect 9862 6352 9918 6361
rect 9862 6287 9918 6296
rect 9876 6254 9904 6287
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 5953 9904 6054
rect 9862 5944 9918 5953
rect 9862 5879 9918 5888
rect 9770 5672 9826 5681
rect 9770 5607 9826 5616
rect 9784 5574 9812 5607
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9692 4321 9720 4490
rect 9678 4312 9734 4321
rect 9678 4247 9734 4256
rect 9312 4208 9364 4214
rect 9680 4208 9732 4214
rect 9312 4150 9364 4156
rect 9416 4168 9680 4196
rect 9324 2990 9352 4150
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9416 2836 9444 4168
rect 9680 4150 9732 4156
rect 9678 3904 9734 3913
rect 9678 3839 9734 3848
rect 9692 3398 9720 3839
rect 9876 3738 9904 5879
rect 9968 3738 9996 8026
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10060 7274 10088 7754
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10060 6322 10088 7210
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10152 5896 10180 9608
rect 10244 9518 10272 9998
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10232 8560 10284 8566
rect 10336 8537 10364 17682
rect 10232 8502 10284 8508
rect 10322 8528 10378 8537
rect 10060 5868 10180 5896
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10060 3618 10088 5868
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10152 4826 10180 5714
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 9968 3590 10088 3618
rect 9968 3534 9996 3590
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9954 3360 10010 3369
rect 9692 3058 9720 3334
rect 9954 3295 10010 3304
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9588 2848 9640 2854
rect 9416 2808 9588 2836
rect 9588 2790 9640 2796
rect 9600 2446 9628 2790
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9232 1278 9628 1306
rect 9600 800 9628 1278
rect 9968 800 9996 3295
rect 10060 2650 10088 3470
rect 10152 3126 10180 4762
rect 10244 3602 10272 8502
rect 10322 8463 10378 8472
rect 10336 5710 10364 8463
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10428 4010 10456 18022
rect 10796 17134 10824 18702
rect 12728 18698 12756 19178
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 17882 11100 18090
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 16522 11008 17002
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 16114 11008 16458
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 13802 10548 14350
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13802 10640 14214
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10980 13716 11008 15914
rect 10888 13688 11008 13716
rect 10782 12200 10838 12209
rect 10782 12135 10838 12144
rect 10796 11898 10824 12135
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 10606 10548 11698
rect 10888 11336 10916 13688
rect 10966 12472 11022 12481
rect 10966 12407 10968 12416
rect 11020 12407 11022 12416
rect 10968 12378 11020 12384
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10980 12102 11008 12174
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10612 11308 10916 11336
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 9722 10548 10542
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10612 9466 10640 11308
rect 10980 11234 11008 12038
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10888 11206 11008 11234
rect 10520 9438 10640 9466
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10336 3534 10364 3878
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 2582 10180 2790
rect 10244 2650 10272 3334
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 10336 2446 10364 2994
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10428 800 10456 3538
rect 10520 2292 10548 9438
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 9178 10640 9318
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 4622 10640 7142
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10704 2582 10732 11154
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 10130 10824 10542
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10796 9722 10824 9930
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10888 9602 10916 11206
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10796 9574 10916 9602
rect 10980 9586 11008 9862
rect 10968 9580 11020 9586
rect 10796 8566 10824 9574
rect 10968 9522 11020 9528
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 6662 10824 8230
rect 10888 7546 10916 9318
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10876 7200 10928 7206
rect 10980 7188 11008 8366
rect 11072 7546 11100 17818
rect 12728 17678 12756 18634
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11164 12356 11192 16526
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11716 16250 11744 17070
rect 12084 16998 12112 17138
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12084 16794 12112 16934
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11980 16584 12032 16590
rect 11978 16552 11980 16561
rect 12032 16552 12034 16561
rect 11978 16487 12034 16496
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11348 15638 11376 15846
rect 11440 15706 11468 15846
rect 11808 15706 11836 16390
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11992 15434 12020 15914
rect 12084 15502 12112 16730
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12452 16114 12480 16662
rect 12636 16590 12664 17002
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11900 13938 11928 14418
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11624 13462 11652 13670
rect 11612 13456 11664 13462
rect 11664 13416 11744 13444
rect 11612 13398 11664 13404
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11244 12368 11296 12374
rect 11164 12328 11244 12356
rect 11244 12310 11296 12316
rect 11520 12300 11572 12306
rect 11572 12260 11652 12288
rect 11520 12242 11572 12248
rect 11624 12102 11652 12260
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11164 9042 11192 11766
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11624 9382 11652 12038
rect 11716 11558 11744 13416
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10130 11744 10406
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11624 7313 11652 9046
rect 11716 8974 11744 10066
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11610 7304 11666 7313
rect 11610 7239 11666 7248
rect 11152 7200 11204 7206
rect 10928 7160 11152 7188
rect 10876 7142 10928 7148
rect 11152 7142 11204 7148
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10796 4826 10824 6054
rect 10888 5914 10916 6054
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10980 5710 11008 6598
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6322 11652 6938
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11348 5778 11376 6258
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11336 5772 11388 5778
rect 11164 5732 11336 5760
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10980 5166 11008 5646
rect 11164 5370 11192 5732
rect 11336 5714 11388 5720
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11624 5166 11652 5782
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10980 4690 11008 5102
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10796 3602 10824 4626
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10888 3534 10916 4218
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3058 10916 3470
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 3194 11100 3402
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11440 2990 11468 3062
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 11716 2514 11744 8774
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10520 2264 10916 2292
rect 10888 800 10916 2264
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11336 1284 11388 1290
rect 11336 1226 11388 1232
rect 11348 800 11376 1226
rect 11808 800 11836 13670
rect 11900 13326 11928 13874
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 11694 11928 12582
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 8362 11928 9318
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11992 7993 12020 15370
rect 12636 14822 12664 16526
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14278 12664 14758
rect 12820 14550 12848 14894
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 12084 11762 12112 12310
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11978 7984 12034 7993
rect 11978 7919 12034 7928
rect 11980 7744 12032 7750
rect 11978 7712 11980 7721
rect 12032 7712 12034 7721
rect 11978 7647 12034 7656
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11900 5914 11928 6326
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 12084 5681 12112 11494
rect 12070 5672 12126 5681
rect 12070 5607 12126 5616
rect 12176 1290 12204 12786
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12306 12480 12718
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12360 11898 12388 12242
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12544 11354 12572 12650
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12728 10010 12756 12242
rect 12820 12170 12848 12582
rect 12808 12164 12860 12170
rect 12808 12106 12860 12112
rect 12728 9982 12848 10010
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12254 9480 12310 9489
rect 12254 9415 12256 9424
rect 12308 9415 12310 9424
rect 12256 9386 12308 9392
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12360 8090 12388 8366
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 1284 12216 1290
rect 12164 1226 12216 1232
rect 12268 800 12296 7482
rect 12360 7342 12388 8026
rect 12452 7546 12480 9658
rect 12544 9382 12572 9862
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 8430 12572 9318
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 6934 12388 7278
rect 12636 7002 12664 8774
rect 12728 8430 12756 9862
rect 12820 9178 12848 9982
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12728 7818 12756 8366
rect 12912 8294 12940 15302
rect 13096 15162 13124 17682
rect 13556 17610 13584 18838
rect 14476 18834 14504 19246
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 13648 18426 13676 18770
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11626 13032 12174
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13004 11150 13032 11562
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 9353 13032 9454
rect 12990 9344 13046 9353
rect 12990 9279 13046 9288
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 13004 7410 13032 8978
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12714 7304 12770 7313
rect 12714 7239 12770 7248
rect 12728 7206 12756 7239
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 13096 6746 13124 15098
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 12238 13216 14214
rect 13464 13802 13492 14418
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 13464 13326 13492 13738
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12306 13492 12786
rect 13556 12646 13584 14486
rect 13648 14226 13676 18362
rect 13740 18290 13768 18702
rect 15212 18698 15240 19858
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 14200 18222 14228 18566
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13740 17882 13768 18022
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 14200 17678 14228 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 15120 17814 15148 18294
rect 15304 17882 15332 19790
rect 16040 19514 16068 19790
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15580 18766 15608 19178
rect 16040 18902 16068 19450
rect 17144 19310 17172 22000
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 13924 15706 13952 17002
rect 14108 16658 14136 17614
rect 15488 17338 15516 18022
rect 15580 17678 15608 18702
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15764 17882 15792 18090
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 16500 17202 16528 18158
rect 16592 17678 16620 18770
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15304 16794 15332 16934
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 16500 16658 16528 16934
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 15978 14136 16390
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14016 15706 14044 15914
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14108 15502 14136 15914
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14346 13768 14826
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15028 14618 15056 14894
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 14612 15068 14618
rect 15016 14554 15068 14560
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13648 14198 13768 14226
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13530 13676 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13740 12458 13768 14198
rect 14292 14074 14320 14418
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13818 13832 13874 13841
rect 13818 13767 13874 13776
rect 13832 13734 13860 13767
rect 13820 13728 13872 13734
rect 13872 13676 14044 13682
rect 13820 13670 14044 13676
rect 13832 13654 14044 13670
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13731 12430 13768 12458
rect 13731 12424 13759 12430
rect 13648 12396 13759 12424
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13188 11558 13216 12174
rect 13464 11898 13492 12242
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11354 13308 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13188 10130 13216 10678
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13188 9586 13216 10066
rect 13648 9636 13676 12396
rect 13832 11354 13860 12718
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12481 13952 12582
rect 13910 12472 13966 12481
rect 13910 12407 13966 12416
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13464 9608 13676 9636
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13188 8974 13216 9522
rect 13372 9382 13400 9522
rect 13464 9489 13492 9608
rect 13832 9518 13860 11290
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13924 10690 13952 10746
rect 14016 10690 14044 13654
rect 14108 13394 14136 13874
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14384 13190 14412 14350
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 14074 14872 14214
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 13462 15056 13738
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12986 14504 13126
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 15120 12850 15148 14758
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15120 12356 15148 12786
rect 15200 12368 15252 12374
rect 15120 12328 15200 12356
rect 15200 12310 15252 12316
rect 15304 12306 15332 15846
rect 15396 15570 15424 16186
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15948 15570 15976 15982
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 15396 14618 15424 15506
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15396 13870 15424 14554
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 10962 14596 12038
rect 15304 11762 15332 12242
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14476 10934 14596 10962
rect 14476 10742 14504 10934
rect 13924 10662 14044 10690
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13924 9654 13952 10406
rect 14016 9926 14044 10662
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13820 9512 13872 9518
rect 13450 9480 13506 9489
rect 13820 9454 13872 9460
rect 13450 9415 13506 9424
rect 14004 9444 14056 9450
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7886 13216 8230
rect 13268 8016 13320 8022
rect 13266 7984 13268 7993
rect 13320 7984 13322 7993
rect 13266 7919 13322 7928
rect 13176 7880 13228 7886
rect 13228 7828 13400 7834
rect 13176 7822 13400 7828
rect 13188 7818 13400 7822
rect 13188 7812 13412 7818
rect 13188 7806 13360 7812
rect 13360 7754 13412 7760
rect 13464 7698 13492 9415
rect 14004 9386 14056 9392
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 8430 13768 9318
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8566 13860 8910
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13740 7954 13768 8366
rect 13832 7970 13860 8502
rect 14016 8022 14044 9386
rect 14108 8906 14136 10066
rect 14568 9994 14596 10610
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15396 10198 15424 13262
rect 15948 12986 15976 13262
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 12442 15792 12582
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 12209 15700 12242
rect 15658 12200 15714 12209
rect 16040 12170 16068 16594
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 14822 16436 15506
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16132 13326 16160 13670
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16408 13258 16436 14758
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16408 12850 16436 13194
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16592 12986 16620 13126
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 15658 12135 15714 12144
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15488 10674 15516 10950
rect 15672 10810 15700 11154
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15764 10266 15792 11086
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15200 10192 15252 10198
rect 15384 10192 15436 10198
rect 15252 10140 15332 10146
rect 15200 10134 15332 10140
rect 15384 10134 15436 10140
rect 15212 10118 15332 10134
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14568 9518 14596 9930
rect 15304 9926 15332 10118
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14556 9512 14608 9518
rect 14278 9480 14334 9489
rect 14556 9454 14608 9460
rect 14278 9415 14334 9424
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14004 8016 14056 8022
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13832 7942 13952 7970
rect 14004 7958 14056 7964
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 13004 6718 13124 6746
rect 13188 7670 13492 7698
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 12452 6458 12480 6666
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12544 6361 12572 6394
rect 12530 6352 12586 6361
rect 12530 6287 12586 6296
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 3602 12480 5510
rect 12820 5166 12848 5646
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12912 4826 12940 5510
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13004 4758 13032 6718
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12544 2514 12572 2858
rect 13004 2514 13032 3606
rect 13096 2990 13124 6598
rect 13188 6322 13216 7670
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13280 6254 13308 6598
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 4758 13308 6054
rect 13464 5148 13492 7210
rect 13648 7002 13676 7686
rect 13832 7342 13860 7942
rect 13924 7886 13952 7942
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 14292 7750 14320 9415
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 13820 7336 13872 7342
rect 13912 7336 13964 7342
rect 13820 7278 13872 7284
rect 13910 7304 13912 7313
rect 13964 7304 13966 7313
rect 13910 7239 13966 7248
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13740 6798 13768 7142
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13556 5710 13584 6122
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13544 5160 13596 5166
rect 13464 5120 13544 5148
rect 13544 5102 13596 5108
rect 13740 5098 13768 6122
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13648 4622 13676 4966
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 3602 13676 4422
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12728 800 12756 2246
rect 13188 800 13216 2790
rect 13740 2514 13768 3470
rect 13924 2990 13952 6666
rect 14292 5914 14320 7686
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14370 5944 14426 5953
rect 14280 5908 14332 5914
rect 14684 5936 14980 5956
rect 14370 5879 14372 5888
rect 14280 5850 14332 5856
rect 14424 5879 14426 5888
rect 14372 5850 14424 5856
rect 15120 5846 15148 6054
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15106 4856 15162 4865
rect 15212 4826 15240 9862
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15304 7274 15332 7822
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15396 6322 15424 10134
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9654 15884 11086
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15856 8022 15884 9590
rect 15844 8016 15896 8022
rect 15936 8016 15988 8022
rect 15844 7958 15896 7964
rect 15934 7984 15936 7993
rect 15988 7984 15990 7993
rect 15934 7919 15990 7928
rect 15474 7712 15530 7721
rect 15474 7647 15530 7656
rect 15488 7206 15516 7647
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15106 4791 15162 4800
rect 15200 4820 15252 4826
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14568 3670 14596 3878
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 15028 3126 15056 3878
rect 15120 3738 15148 4791
rect 15200 4762 15252 4768
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 3738 15424 4422
rect 15488 4078 15516 7142
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4622 15976 4966
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4078 15976 4558
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15212 3194 15240 3538
rect 15476 3528 15528 3534
rect 16040 3505 16068 12106
rect 16684 11626 16712 15642
rect 16776 13530 16804 18022
rect 16868 16726 16896 18158
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16960 16998 16988 17750
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16868 14278 16896 16662
rect 16960 16590 16988 16934
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16948 13864 17000 13870
rect 17144 13818 17172 18566
rect 17880 18222 17908 22471
rect 19246 22128 19302 22137
rect 19246 22063 19302 22072
rect 19062 21584 19118 21593
rect 19062 21519 19118 21528
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17972 18222 18000 19654
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 19076 19174 19104 21519
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 17236 15706 17264 15914
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17236 15026 17264 15642
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17236 14414 17264 14962
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17000 13812 17172 13818
rect 16948 13806 17172 13812
rect 16960 13790 17172 13806
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16776 13190 16804 13466
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16960 12442 16988 13262
rect 17052 12714 17080 13670
rect 17144 13326 17172 13790
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 12850 17172 13262
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16960 11694 16988 12378
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 17052 11558 17080 12650
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 9586 16252 10610
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9722 16620 9862
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8362 16620 9318
rect 16684 8430 16712 10406
rect 16868 10062 16896 11086
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 8974 16896 9998
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16868 8294 16896 8910
rect 16960 8786 16988 9658
rect 17052 9160 17080 11494
rect 17236 9382 17264 13466
rect 17328 11354 17356 17682
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17788 17134 17816 17478
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 12918 17448 14758
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13530 17540 14418
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17604 12714 17632 16594
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17696 12238 17724 17002
rect 17788 16046 17816 17070
rect 17972 16522 18000 17478
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 12866 17816 15982
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 14958 18000 15302
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18524 15162 18552 15574
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18616 15026 18644 15506
rect 18708 15162 18736 15506
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18800 14498 18828 15438
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18708 14470 18828 14498
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 13530 18552 14418
rect 18708 14414 18736 14470
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18616 14074 18644 14350
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17880 12986 17908 13262
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17788 12838 17908 12866
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12442 17816 12582
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17406 11792 17462 11801
rect 17406 11727 17462 11736
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 10713 17448 11727
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17406 10704 17462 10713
rect 17512 10674 17540 11154
rect 17406 10639 17462 10648
rect 17500 10668 17552 10674
rect 17420 10606 17448 10639
rect 17500 10610 17552 10616
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17512 9178 17540 10066
rect 17604 9194 17632 11562
rect 17696 9450 17724 12174
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17696 9353 17724 9386
rect 17682 9344 17738 9353
rect 17682 9279 17738 9288
rect 17500 9172 17552 9178
rect 17052 9132 17356 9160
rect 16960 8758 17080 8786
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16224 7342 16252 8230
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16224 6934 16252 7278
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16500 6662 16528 7278
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5914 16252 6054
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16500 5710 16528 6598
rect 16592 6322 16620 6802
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16776 6066 16804 6870
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 6254 16988 6734
rect 17052 6254 17080 8758
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16684 6038 16804 6066
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16684 5574 16712 6038
rect 17144 5914 17172 7686
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17144 5778 17172 5850
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 15476 3470 15528 3476
rect 16026 3496 16082 3505
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15396 2990 15424 3334
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14476 2514 14504 2858
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 13556 800 13584 2246
rect 14016 800 14044 2246
rect 14476 800 14504 2246
rect 14936 800 14964 2246
rect 15396 800 15424 2790
rect 15488 2514 15516 3470
rect 16026 3431 16082 3440
rect 16132 2514 16160 5510
rect 16684 5234 16712 5510
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16316 3738 16344 4626
rect 16684 4622 16712 5170
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16684 3942 16712 4558
rect 17052 3942 17080 4694
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 17052 3534 17080 3878
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17236 2990 17264 8502
rect 17328 8378 17356 9132
rect 17604 9166 17724 9194
rect 17500 9114 17552 9120
rect 17512 8498 17540 9114
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8498 17632 8978
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17328 8350 17540 8378
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 8090 17448 8230
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17328 4826 17356 6258
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17420 4010 17448 7890
rect 17408 4004 17460 4010
rect 17408 3946 17460 3952
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17408 2916 17460 2922
rect 17408 2858 17460 2864
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 800 15884 2246
rect 16316 800 16344 2790
rect 17420 2514 17448 2858
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16684 800 16712 2246
rect 17144 800 17172 2246
rect 6274 232 6330 241
rect 6274 167 6330 176
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17512 241 17540 8350
rect 17604 7886 17632 8434
rect 17696 8090 17724 9166
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7546 17632 7822
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 1170 17724 2246
rect 17788 2009 17816 12378
rect 17880 12170 17908 12838
rect 17972 12442 18000 13330
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12442 18552 13330
rect 18708 13326 18736 14350
rect 18892 14346 18920 15438
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18708 12374 18736 12786
rect 18892 12782 18920 13330
rect 18984 13297 19012 18022
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19076 17785 19104 17818
rect 19062 17776 19118 17785
rect 19062 17711 19118 17720
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19076 14958 19104 15846
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14113 19104 14758
rect 19062 14104 19118 14113
rect 19062 14039 19118 14048
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 18970 13288 19026 13297
rect 19076 13258 19104 13874
rect 18970 13223 19026 13232
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18970 13152 19026 13161
rect 18970 13087 19026 13096
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17972 10606 18000 11494
rect 18708 11393 18736 11562
rect 18694 11384 18750 11393
rect 18604 11348 18656 11354
rect 18694 11319 18750 11328
rect 18604 11290 18656 11296
rect 18512 11212 18564 11218
rect 18512 11154 18564 11160
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10810 18552 11154
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18510 10704 18566 10713
rect 18510 10639 18566 10648
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17958 10432 18014 10441
rect 17958 10367 18014 10376
rect 17972 10198 18000 10367
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17958 10024 18014 10033
rect 17958 9959 18014 9968
rect 17972 7206 18000 9959
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9110 18552 10639
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18050 8120 18106 8129
rect 18432 8090 18460 8230
rect 18050 8055 18106 8064
rect 18420 8084 18472 8090
rect 18064 7954 18092 8055
rect 18420 8026 18472 8032
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 18524 7478 18552 7511
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17958 6760 18014 6769
rect 17958 6695 18014 6704
rect 17972 6390 18000 6695
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5778 17908 6258
rect 18052 6112 18104 6118
rect 18420 6112 18472 6118
rect 18052 6054 18104 6060
rect 18418 6080 18420 6089
rect 18472 6080 18474 6089
rect 18064 5914 18092 6054
rect 18418 6015 18474 6024
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18524 5817 18552 6394
rect 18510 5808 18566 5817
rect 17868 5772 17920 5778
rect 18510 5743 18566 5752
rect 17868 5714 17920 5720
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18524 4282 18552 4422
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18616 3754 18644 11290
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10742 18736 11086
rect 18696 10736 18748 10742
rect 18696 10678 18748 10684
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 6905 18736 10406
rect 18800 9382 18828 12582
rect 18892 12345 18920 12718
rect 18878 12336 18934 12345
rect 18878 12271 18934 12280
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18892 11762 18920 12174
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18892 10606 18920 11562
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18694 6896 18750 6905
rect 18694 6831 18750 6840
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18708 6254 18736 6734
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 3942 18736 6054
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18616 3726 18736 3754
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18340 2514 18368 2858
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17774 2000 17830 2009
rect 17774 1935 17830 1944
rect 17604 1142 17724 1170
rect 17972 1170 18000 2314
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18092 1170
rect 17604 800 17632 1142
rect 18064 800 18092 1142
rect 18524 800 18552 3334
rect 18616 3058 18644 3538
rect 18708 3126 18736 3726
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18800 2990 18828 8774
rect 18892 6186 18920 9114
rect 18984 8498 19012 13087
rect 19076 12850 19104 13194
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19168 12594 19196 19246
rect 19260 18970 19288 22063
rect 19614 21176 19670 21185
rect 19614 21111 19670 21120
rect 19628 20058 19656 21111
rect 20166 20632 20222 20641
rect 20166 20567 20222 20576
rect 19706 20224 19762 20233
rect 19706 20159 19762 20168
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19260 13938 19288 15030
rect 19352 14958 19380 19246
rect 19444 17882 19472 19858
rect 19720 19514 19748 20159
rect 20180 20058 20208 20567
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19536 18329 19564 18770
rect 19522 18320 19578 18329
rect 19522 18255 19578 18264
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19444 16250 19472 17002
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19444 15434 19472 16186
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19352 13818 19380 14894
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19260 13790 19380 13818
rect 19260 12730 19288 13790
rect 19444 13734 19472 14214
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19536 13546 19564 18158
rect 19628 13682 19656 18770
rect 19720 18057 19748 19246
rect 19996 18902 20024 19858
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 20088 18426 20116 19858
rect 20166 19816 20222 19825
rect 20166 19751 20222 19760
rect 20180 19514 20208 19751
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20536 19304 20588 19310
rect 20640 19281 20668 19654
rect 20536 19246 20588 19252
rect 20626 19272 20682 19281
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20168 18352 20220 18358
rect 20166 18320 20168 18329
rect 20220 18320 20222 18329
rect 20166 18255 20222 18264
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19706 18048 19762 18057
rect 19706 17983 19762 17992
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 15638 19748 17002
rect 19890 16960 19946 16969
rect 19890 16895 19946 16904
rect 19904 16794 19932 16895
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19720 14634 19748 14826
rect 19812 14822 19840 16662
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19996 16114 20024 16594
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19984 15972 20036 15978
rect 19984 15914 20036 15920
rect 19890 15600 19946 15609
rect 19890 15535 19946 15544
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19720 14606 19840 14634
rect 19904 14618 19932 15535
rect 19996 15502 20024 15914
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 14958 20024 15302
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 13802 19748 14418
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19628 13654 19748 13682
rect 19444 13518 19564 13546
rect 19260 12702 19380 12730
rect 19168 12566 19288 12594
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 19154 12336 19210 12345
rect 19076 10470 19104 12310
rect 19154 12271 19210 12280
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18984 6186 19012 8298
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 4146 18920 5510
rect 18984 5098 19012 5646
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18880 3936 18932 3942
rect 18984 3913 19012 4014
rect 18880 3878 18932 3884
rect 18970 3904 19026 3913
rect 18892 3040 18920 3878
rect 18970 3839 19026 3848
rect 18892 3012 19012 3040
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18892 2514 18920 2858
rect 18984 2854 19012 3012
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 19076 1601 19104 9318
rect 19168 9178 19196 12271
rect 19260 11898 19288 12566
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11082 19288 11562
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19352 10962 19380 12702
rect 19444 12458 19472 13518
rect 19435 12430 19472 12458
rect 19435 12356 19463 12430
rect 19435 12328 19472 12356
rect 19260 10934 19380 10962
rect 19260 9722 19288 10934
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19154 9072 19210 9081
rect 19154 9007 19210 9016
rect 19168 3602 19196 9007
rect 19352 8430 19380 9454
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19352 7342 19380 8366
rect 19444 7342 19472 12328
rect 19614 11112 19670 11121
rect 19614 11047 19670 11056
rect 19628 11014 19656 11047
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10674 19656 10950
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 9110 19564 10406
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19628 9178 19656 9862
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19352 6934 19380 7278
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19444 6866 19472 7142
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6390 19472 6802
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19628 6322 19656 7686
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19062 1592 19118 1601
rect 19062 1527 19118 1536
rect 19168 1442 19196 3334
rect 19260 2990 19288 6054
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19352 2802 19380 6122
rect 19720 3942 19748 13654
rect 19812 12782 19840 14606
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 20088 12594 20116 18158
rect 20548 17814 20576 19246
rect 20626 19207 20682 19216
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18873 20760 19110
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17921 20668 18022
rect 20626 17912 20682 17921
rect 20626 17847 20682 17856
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20166 17368 20222 17377
rect 20166 17303 20168 17312
rect 20220 17303 20222 17312
rect 20168 17274 20220 17280
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19996 12566 20116 12594
rect 19996 12356 20024 12566
rect 19904 12328 20024 12356
rect 19904 9466 19932 12328
rect 20180 12102 20208 17070
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20640 16561 20668 16934
rect 20626 16552 20682 16561
rect 20626 16487 20682 16496
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16017 20484 16390
rect 20536 16040 20588 16046
rect 20442 16008 20498 16017
rect 20260 15972 20312 15978
rect 20536 15982 20588 15988
rect 20442 15943 20498 15952
rect 20260 15914 20312 15920
rect 20272 15570 20300 15914
rect 20548 15706 20576 15982
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20272 14482 20300 14826
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20364 12986 20392 15438
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20456 15065 20484 15302
rect 20442 15056 20498 15065
rect 20442 14991 20498 15000
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14657 20944 14758
rect 20902 14648 20958 14657
rect 20902 14583 20958 14592
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20456 14113 20484 14214
rect 20442 14104 20498 14113
rect 20442 14039 20498 14048
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20640 13705 20668 13942
rect 20626 13696 20682 13705
rect 20626 13631 20682 13640
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19996 10266 20024 10474
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20088 10266 20116 10406
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20272 10130 20300 12582
rect 20364 12306 20392 12786
rect 20720 12776 20772 12782
rect 20626 12744 20682 12753
rect 20720 12718 20772 12724
rect 20626 12679 20628 12688
rect 20680 12679 20682 12688
rect 20628 12650 20680 12656
rect 20732 12345 20760 12718
rect 20718 12336 20774 12345
rect 20352 12300 20404 12306
rect 20718 12271 20774 12280
rect 20352 12242 20404 12248
rect 20364 11898 20392 12242
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20350 10840 20406 10849
rect 20350 10775 20406 10784
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20180 9518 20208 9998
rect 19812 9450 19932 9466
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19800 9444 19932 9450
rect 19852 9438 19932 9444
rect 19800 9386 19852 9392
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19812 8430 19840 8910
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 20364 8090 20392 10775
rect 20548 10674 20576 12038
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20548 10062 20576 10610
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 8974 21036 9318
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20640 7886 20668 8230
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7342 20668 7822
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 19982 7168 20038 7177
rect 19982 7103 20038 7112
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19812 5710 19840 6258
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19904 4078 19932 6054
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 18984 1414 19196 1442
rect 19260 2774 19380 2802
rect 18984 800 19012 1414
rect 17498 232 17554 241
rect 17498 167 17554 176
rect 17590 0 17646 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19260 649 19288 2774
rect 19536 1714 19564 3334
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19444 1686 19564 1714
rect 19444 800 19472 1686
rect 19720 1057 19748 2790
rect 19706 1048 19762 1057
rect 19706 983 19762 992
rect 19812 800 19840 3878
rect 19996 3602 20024 7103
rect 20548 6254 20576 7210
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5914 20576 6054
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20626 5264 20682 5273
rect 20626 5199 20682 5208
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20180 4690 20208 4966
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20180 4146 20208 4626
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19904 2514 19932 2858
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 20272 800 20300 4966
rect 20548 4321 20576 5102
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20640 4078 20668 5199
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 800 20760 4014
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21192 800 21220 3402
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21652 800 21680 2926
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 800 22140 2790
rect 22572 800 22600 2858
rect 19246 640 19302 649
rect 19246 575 19302 584
rect 19430 0 19486 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
<< via2 >>
rect 4250 22480 4306 22536
rect 3054 22072 3110 22128
rect 2962 21528 3018 21584
rect 2778 21120 2834 21176
rect 2870 20168 2926 20224
rect 2042 19760 2098 19816
rect 2778 19216 2834 19272
rect 4066 20576 4122 20632
rect 1950 18808 2006 18864
rect 1950 18300 1952 18320
rect 1952 18300 2004 18320
rect 2004 18300 2006 18320
rect 1950 18264 2006 18300
rect 1582 17876 1638 17912
rect 1582 17856 1584 17876
rect 1584 17856 1636 17876
rect 1636 17856 1638 17876
rect 1950 16516 2006 16552
rect 1950 16496 1952 16516
rect 1952 16496 2004 16516
rect 2004 16496 2006 16516
rect 1950 15952 2006 16008
rect 1950 15544 2006 15600
rect 1674 15000 1730 15056
rect 1950 14048 2006 14104
rect 2870 17312 2926 17368
rect 2778 16904 2834 16960
rect 2778 13640 2834 13696
rect 3330 14592 3386 14648
rect 2870 13232 2926 13288
rect 2410 8336 2466 8392
rect 2042 7112 2098 7168
rect 1306 6160 1362 6216
rect 2962 8880 3018 8936
rect 17866 22480 17922 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 2778 3440 2834 3496
rect 1950 2760 2006 2816
rect 2962 2796 2964 2816
rect 2964 2796 3016 2816
rect 3016 2796 3018 2816
rect 2962 2760 3018 2796
rect 2870 1536 2926 1592
rect 3146 2488 3202 2544
rect 3238 992 3294 1048
rect 4066 12708 4122 12744
rect 4066 12688 4068 12708
rect 4068 12688 4120 12708
rect 4120 12688 4122 12708
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11736 4122 11792
rect 4066 10804 4122 10840
rect 4066 10784 4068 10804
rect 4068 10784 4120 10804
rect 4120 10784 4122 10804
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4066 10376 4122 10432
rect 3974 9968 4030 10024
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4066 9460 4068 9480
rect 4068 9460 4120 9480
rect 4120 9460 4122 9480
rect 4066 9424 4122 9460
rect 4066 9052 4068 9072
rect 4068 9052 4120 9072
rect 4120 9052 4122 9072
rect 4066 9016 4122 9052
rect 4710 8916 4712 8936
rect 4712 8916 4764 8936
rect 4764 8916 4766 8936
rect 4710 8880 4766 8916
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4710 8064 4766 8120
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4066 6704 4122 6760
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 3974 5752 4030 5808
rect 3974 5208 4030 5264
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4066 4256 4122 4312
rect 3606 1944 3662 2000
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 5354 9424 5410 9480
rect 5078 2896 5134 2952
rect 6090 14048 6146 14104
rect 6182 4800 6238 4856
rect 4066 584 4122 640
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8390 12280 8446 12336
rect 9586 14068 9642 14104
rect 9586 14048 9588 14068
rect 9588 14048 9640 14068
rect 9640 14048 9642 14068
rect 8666 11600 8722 11656
rect 7838 9424 7894 9480
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7930 8472 7986 8528
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8390 8336 8446 8392
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8758 7384 8814 7440
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9862 10648 9918 10704
rect 9310 8880 9366 8936
rect 9862 9324 9864 9344
rect 9864 9324 9916 9344
rect 9916 9324 9918 9344
rect 9862 9288 9918 9324
rect 9770 7812 9826 7848
rect 9770 7792 9772 7812
rect 9772 7792 9824 7812
rect 9824 7792 9826 7812
rect 9770 7248 9826 7304
rect 9126 6060 9128 6080
rect 9128 6060 9180 6080
rect 9180 6060 9182 6080
rect 9126 6024 9182 6060
rect 8850 3576 8906 3632
rect 9862 6296 9918 6352
rect 9862 5888 9918 5944
rect 9770 5616 9826 5672
rect 9678 4256 9734 4312
rect 9678 3848 9734 3904
rect 9954 3304 10010 3360
rect 10322 8472 10378 8528
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 10782 12144 10838 12200
rect 10966 12436 11022 12472
rect 10966 12416 10968 12436
rect 10968 12416 11020 12436
rect 11020 12416 11022 12436
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11978 16532 11980 16552
rect 11980 16532 12032 16552
rect 12032 16532 12034 16552
rect 11978 16496 12034 16532
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11610 7248 11666 7304
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11978 7928 12034 7984
rect 11978 7692 11980 7712
rect 11980 7692 12032 7712
rect 12032 7692 12034 7712
rect 11978 7656 12034 7692
rect 12070 5616 12126 5672
rect 12254 9444 12310 9480
rect 12254 9424 12256 9444
rect 12256 9424 12308 9444
rect 12308 9424 12310 9444
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 12990 9288 13046 9344
rect 12714 7248 12770 7304
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 13818 13776 13874 13832
rect 13910 12416 13966 12472
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 13450 9424 13506 9480
rect 13266 7964 13268 7984
rect 13268 7964 13320 7984
rect 13320 7964 13322 7984
rect 13266 7928 13322 7964
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 15658 12144 15714 12200
rect 14278 9424 14334 9480
rect 12530 6296 12586 6352
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 13910 7284 13912 7304
rect 13912 7284 13964 7304
rect 13964 7284 13966 7304
rect 13910 7248 13966 7284
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14370 5908 14426 5944
rect 14370 5888 14372 5908
rect 14372 5888 14424 5908
rect 14424 5888 14426 5908
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 15106 4800 15162 4856
rect 15934 7964 15936 7984
rect 15936 7964 15988 7984
rect 15988 7964 15990 7984
rect 15934 7928 15990 7964
rect 15474 7656 15530 7712
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 19246 22072 19302 22128
rect 19062 21528 19118 21584
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 17406 11736 17462 11792
rect 17406 10648 17462 10704
rect 17682 9288 17738 9344
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 16026 3440 16082 3496
rect 6274 176 6330 232
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 19062 17720 19118 17776
rect 19062 14048 19118 14104
rect 18970 13232 19026 13288
rect 18970 13096 19026 13152
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18694 11328 18750 11384
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18510 10648 18566 10704
rect 17958 10376 18014 10432
rect 17958 9968 18014 10024
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18050 8064 18106 8120
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18510 7520 18566 7576
rect 17958 6704 18014 6760
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18418 6060 18420 6080
rect 18420 6060 18472 6080
rect 18472 6060 18474 6080
rect 18418 6024 18474 6060
rect 18510 5752 18566 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18878 12280 18934 12336
rect 18694 6840 18750 6896
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17774 1944 17830 2000
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 19614 21120 19670 21176
rect 20166 20576 20222 20632
rect 19706 20168 19762 20224
rect 19522 18264 19578 18320
rect 20166 19760 20222 19816
rect 20166 18300 20168 18320
rect 20168 18300 20220 18320
rect 20220 18300 20222 18320
rect 20166 18264 20222 18300
rect 19706 17992 19762 18048
rect 19890 16904 19946 16960
rect 19890 15544 19946 15600
rect 19154 12280 19210 12336
rect 18970 3848 19026 3904
rect 19154 9016 19210 9072
rect 19614 11056 19670 11112
rect 19062 1536 19118 1592
rect 20626 19216 20682 19272
rect 20718 18808 20774 18864
rect 20626 17856 20682 17912
rect 20166 17332 20222 17368
rect 20166 17312 20168 17332
rect 20168 17312 20220 17332
rect 20220 17312 20222 17332
rect 20626 16496 20682 16552
rect 20442 15952 20498 16008
rect 20442 15000 20498 15056
rect 20902 14592 20958 14648
rect 20442 14048 20498 14104
rect 20626 13640 20682 13696
rect 20626 12708 20682 12744
rect 20626 12688 20628 12708
rect 20628 12688 20680 12708
rect 20680 12688 20682 12708
rect 20718 12280 20774 12336
rect 20350 10784 20406 10840
rect 19982 7112 20038 7168
rect 17498 176 17554 232
rect 19706 992 19762 1048
rect 20626 5208 20682 5264
rect 20534 4256 20590 4312
rect 19246 584 19302 640
<< metal3 >>
rect 0 22538 800 22568
rect 4245 22538 4311 22541
rect 0 22536 4311 22538
rect 0 22480 4250 22536
rect 4306 22480 4311 22536
rect 0 22478 4311 22480
rect 0 22448 800 22478
rect 4245 22475 4311 22478
rect 17861 22538 17927 22541
rect 22000 22538 22800 22568
rect 17861 22536 22800 22538
rect 17861 22480 17866 22536
rect 17922 22480 22800 22536
rect 17861 22478 22800 22480
rect 17861 22475 17927 22478
rect 22000 22448 22800 22478
rect 0 22130 800 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 800 22070
rect 3049 22067 3115 22070
rect 19241 22130 19307 22133
rect 22000 22130 22800 22160
rect 19241 22128 22800 22130
rect 19241 22072 19246 22128
rect 19302 22072 22800 22128
rect 19241 22070 22800 22072
rect 19241 22067 19307 22070
rect 22000 22040 22800 22070
rect 0 21586 800 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 800 21526
rect 2957 21523 3023 21526
rect 19057 21586 19123 21589
rect 22000 21586 22800 21616
rect 19057 21584 22800 21586
rect 19057 21528 19062 21584
rect 19118 21528 22800 21584
rect 19057 21526 22800 21528
rect 19057 21523 19123 21526
rect 22000 21496 22800 21526
rect 0 21178 800 21208
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 19609 21178 19675 21181
rect 22000 21178 22800 21208
rect 19609 21176 22800 21178
rect 19609 21120 19614 21176
rect 19670 21120 22800 21176
rect 19609 21118 22800 21120
rect 19609 21115 19675 21118
rect 22000 21088 22800 21118
rect 0 20634 800 20664
rect 4061 20634 4127 20637
rect 0 20632 4127 20634
rect 0 20576 4066 20632
rect 4122 20576 4127 20632
rect 0 20574 4127 20576
rect 0 20544 800 20574
rect 4061 20571 4127 20574
rect 20161 20634 20227 20637
rect 22000 20634 22800 20664
rect 20161 20632 22800 20634
rect 20161 20576 20166 20632
rect 20222 20576 22800 20632
rect 20161 20574 22800 20576
rect 20161 20571 20227 20574
rect 22000 20544 22800 20574
rect 0 20226 800 20256
rect 2865 20226 2931 20229
rect 0 20224 2931 20226
rect 0 20168 2870 20224
rect 2926 20168 2931 20224
rect 0 20166 2931 20168
rect 0 20136 800 20166
rect 2865 20163 2931 20166
rect 19701 20226 19767 20229
rect 22000 20226 22800 20256
rect 19701 20224 22800 20226
rect 19701 20168 19706 20224
rect 19762 20168 22800 20224
rect 19701 20166 22800 20168
rect 19701 20163 19767 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22000 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 800 19848
rect 2037 19818 2103 19821
rect 0 19816 2103 19818
rect 0 19760 2042 19816
rect 2098 19760 2103 19816
rect 0 19758 2103 19760
rect 0 19728 800 19758
rect 2037 19755 2103 19758
rect 20161 19818 20227 19821
rect 22000 19818 22800 19848
rect 20161 19816 22800 19818
rect 20161 19760 20166 19816
rect 20222 19760 22800 19816
rect 20161 19758 22800 19760
rect 20161 19755 20227 19758
rect 22000 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 800 19304
rect 2773 19274 2839 19277
rect 0 19272 2839 19274
rect 0 19216 2778 19272
rect 2834 19216 2839 19272
rect 0 19214 2839 19216
rect 0 19184 800 19214
rect 2773 19211 2839 19214
rect 20621 19274 20687 19277
rect 22000 19274 22800 19304
rect 20621 19272 22800 19274
rect 20621 19216 20626 19272
rect 20682 19216 22800 19272
rect 20621 19214 22800 19216
rect 20621 19211 20687 19214
rect 22000 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 800 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 800 18806
rect 1945 18803 2011 18806
rect 20713 18866 20779 18869
rect 22000 18866 22800 18896
rect 20713 18864 22800 18866
rect 20713 18808 20718 18864
rect 20774 18808 22800 18864
rect 20713 18806 22800 18808
rect 20713 18803 20779 18806
rect 22000 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 800 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 800 18262
rect 1945 18259 2011 18262
rect 19517 18322 19583 18325
rect 19742 18322 19748 18324
rect 19517 18320 19748 18322
rect 19517 18264 19522 18320
rect 19578 18264 19748 18320
rect 19517 18262 19748 18264
rect 19517 18259 19583 18262
rect 19742 18260 19748 18262
rect 19812 18260 19818 18324
rect 20161 18322 20227 18325
rect 22000 18322 22800 18352
rect 20161 18320 22800 18322
rect 20161 18264 20166 18320
rect 20222 18264 22800 18320
rect 20161 18262 22800 18264
rect 20161 18259 20227 18262
rect 22000 18232 22800 18262
rect 19374 17988 19380 18052
rect 19444 18050 19450 18052
rect 19701 18050 19767 18053
rect 19444 18048 19767 18050
rect 19444 17992 19706 18048
rect 19762 17992 19767 18048
rect 19444 17990 19767 17992
rect 19444 17988 19450 17990
rect 19701 17987 19767 17990
rect 7808 17984 8128 17985
rect 0 17914 800 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1577 17914 1643 17917
rect 0 17912 1643 17914
rect 0 17856 1582 17912
rect 1638 17856 1643 17912
rect 0 17854 1643 17856
rect 0 17824 800 17854
rect 1577 17851 1643 17854
rect 20621 17914 20687 17917
rect 22000 17914 22800 17944
rect 20621 17912 22800 17914
rect 20621 17856 20626 17912
rect 20682 17856 22800 17912
rect 20621 17854 22800 17856
rect 20621 17851 20687 17854
rect 22000 17824 22800 17854
rect 19057 17780 19123 17781
rect 19006 17716 19012 17780
rect 19076 17778 19123 17780
rect 19076 17776 19168 17778
rect 19118 17720 19168 17776
rect 19076 17718 19168 17720
rect 19076 17716 19123 17718
rect 19057 17715 19123 17716
rect 4376 17440 4696 17441
rect 0 17370 800 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 2865 17370 2931 17373
rect 0 17368 2931 17370
rect 0 17312 2870 17368
rect 2926 17312 2931 17368
rect 0 17310 2931 17312
rect 0 17280 800 17310
rect 2865 17307 2931 17310
rect 20161 17370 20227 17373
rect 22000 17370 22800 17400
rect 20161 17368 22800 17370
rect 20161 17312 20166 17368
rect 20222 17312 22800 17368
rect 20161 17310 22800 17312
rect 20161 17307 20227 17310
rect 22000 17280 22800 17310
rect 0 16962 800 16992
rect 2773 16962 2839 16965
rect 0 16960 2839 16962
rect 0 16904 2778 16960
rect 2834 16904 2839 16960
rect 0 16902 2839 16904
rect 0 16872 800 16902
rect 2773 16899 2839 16902
rect 19885 16962 19951 16965
rect 22000 16962 22800 16992
rect 19885 16960 22800 16962
rect 19885 16904 19890 16960
rect 19946 16904 22800 16960
rect 19885 16902 22800 16904
rect 19885 16899 19951 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22000 16872 22800 16902
rect 14672 16831 14992 16832
rect 0 16554 800 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 800 16494
rect 1945 16491 2011 16494
rect 11973 16554 12039 16557
rect 19006 16554 19012 16556
rect 11973 16552 19012 16554
rect 11973 16496 11978 16552
rect 12034 16496 19012 16552
rect 11973 16494 19012 16496
rect 11973 16491 12039 16494
rect 19006 16492 19012 16494
rect 19076 16492 19082 16556
rect 20621 16554 20687 16557
rect 22000 16554 22800 16584
rect 20621 16552 22800 16554
rect 20621 16496 20626 16552
rect 20682 16496 22800 16552
rect 20621 16494 22800 16496
rect 20621 16491 20687 16494
rect 22000 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 800 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 800 15950
rect 1945 15947 2011 15950
rect 20437 16010 20503 16013
rect 22000 16010 22800 16040
rect 20437 16008 22800 16010
rect 20437 15952 20442 16008
rect 20498 15952 22800 16008
rect 20437 15950 22800 15952
rect 20437 15947 20503 15950
rect 22000 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 800 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 0 15512 800 15542
rect 1945 15539 2011 15542
rect 19885 15602 19951 15605
rect 22000 15602 22800 15632
rect 19885 15600 22800 15602
rect 19885 15544 19890 15600
rect 19946 15544 22800 15600
rect 19885 15542 22800 15544
rect 19885 15539 19951 15542
rect 22000 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 800 15088
rect 1669 15058 1735 15061
rect 0 15056 1735 15058
rect 0 15000 1674 15056
rect 1730 15000 1735 15056
rect 0 14998 1735 15000
rect 0 14968 800 14998
rect 1669 14995 1735 14998
rect 20437 15058 20503 15061
rect 22000 15058 22800 15088
rect 20437 15056 22800 15058
rect 20437 15000 20442 15056
rect 20498 15000 22800 15056
rect 20437 14998 22800 15000
rect 20437 14995 20503 14998
rect 22000 14968 22800 14998
rect 7808 14720 8128 14721
rect 0 14650 800 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 3325 14650 3391 14653
rect 0 14648 3391 14650
rect 0 14592 3330 14648
rect 3386 14592 3391 14648
rect 0 14590 3391 14592
rect 0 14560 800 14590
rect 3325 14587 3391 14590
rect 20897 14650 20963 14653
rect 22000 14650 22800 14680
rect 20897 14648 22800 14650
rect 20897 14592 20902 14648
rect 20958 14592 22800 14648
rect 20897 14590 22800 14592
rect 20897 14587 20963 14590
rect 22000 14560 22800 14590
rect 4376 14176 4696 14177
rect 0 14106 800 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1945 14106 2011 14109
rect 0 14104 2011 14106
rect 0 14048 1950 14104
rect 2006 14048 2011 14104
rect 0 14046 2011 14048
rect 0 14016 800 14046
rect 1945 14043 2011 14046
rect 6085 14106 6151 14109
rect 9581 14106 9647 14109
rect 6085 14104 9647 14106
rect 6085 14048 6090 14104
rect 6146 14048 9586 14104
rect 9642 14048 9647 14104
rect 6085 14046 9647 14048
rect 6085 14043 6151 14046
rect 9581 14043 9647 14046
rect 18822 14044 18828 14108
rect 18892 14106 18898 14108
rect 19057 14106 19123 14109
rect 18892 14104 19123 14106
rect 18892 14048 19062 14104
rect 19118 14048 19123 14104
rect 18892 14046 19123 14048
rect 18892 14044 18898 14046
rect 19057 14043 19123 14046
rect 20437 14106 20503 14109
rect 22000 14106 22800 14136
rect 20437 14104 22800 14106
rect 20437 14048 20442 14104
rect 20498 14048 22800 14104
rect 20437 14046 22800 14048
rect 20437 14043 20503 14046
rect 22000 14016 22800 14046
rect 13813 13834 13879 13837
rect 19374 13834 19380 13836
rect 13813 13832 19380 13834
rect 13813 13776 13818 13832
rect 13874 13776 19380 13832
rect 13813 13774 19380 13776
rect 13813 13771 13879 13774
rect 19374 13772 19380 13774
rect 19444 13772 19450 13836
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 20621 13698 20687 13701
rect 22000 13698 22800 13728
rect 20621 13696 22800 13698
rect 20621 13640 20626 13696
rect 20682 13640 22800 13696
rect 20621 13638 22800 13640
rect 20621 13635 20687 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22000 13608 22800 13638
rect 14672 13567 14992 13568
rect 0 13290 800 13320
rect 2865 13290 2931 13293
rect 0 13288 2931 13290
rect 0 13232 2870 13288
rect 2926 13232 2931 13288
rect 0 13230 2931 13232
rect 0 13200 800 13230
rect 2865 13227 2931 13230
rect 18965 13290 19031 13293
rect 22000 13290 22800 13320
rect 18965 13288 22800 13290
rect 18965 13232 18970 13288
rect 19026 13232 22800 13288
rect 18965 13230 22800 13232
rect 18965 13227 19031 13230
rect 22000 13200 22800 13230
rect 18965 13156 19031 13157
rect 18965 13152 19012 13156
rect 19076 13154 19082 13156
rect 18965 13096 18970 13152
rect 18965 13092 19012 13096
rect 19076 13094 19122 13154
rect 19076 13092 19082 13094
rect 18965 13091 19031 13092
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 800 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 800 12686
rect 4061 12683 4127 12686
rect 20621 12746 20687 12749
rect 22000 12746 22800 12776
rect 20621 12744 22800 12746
rect 20621 12688 20626 12744
rect 20682 12688 22800 12744
rect 20621 12686 22800 12688
rect 20621 12683 20687 12686
rect 22000 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 10961 12474 11027 12477
rect 13905 12474 13971 12477
rect 10961 12472 13971 12474
rect 10961 12416 10966 12472
rect 11022 12416 13910 12472
rect 13966 12416 13971 12472
rect 10961 12414 13971 12416
rect 10961 12411 11027 12414
rect 13905 12411 13971 12414
rect 0 12338 800 12368
rect 8385 12338 8451 12341
rect 0 12336 8451 12338
rect 0 12280 8390 12336
rect 8446 12280 8451 12336
rect 0 12278 8451 12280
rect 0 12248 800 12278
rect 8385 12275 8451 12278
rect 18873 12338 18939 12341
rect 19149 12338 19215 12341
rect 18873 12336 19215 12338
rect 18873 12280 18878 12336
rect 18934 12280 19154 12336
rect 19210 12280 19215 12336
rect 18873 12278 19215 12280
rect 18873 12275 18939 12278
rect 19149 12275 19215 12278
rect 20713 12338 20779 12341
rect 22000 12338 22800 12368
rect 20713 12336 22800 12338
rect 20713 12280 20718 12336
rect 20774 12280 22800 12336
rect 20713 12278 22800 12280
rect 20713 12275 20779 12278
rect 22000 12248 22800 12278
rect 10777 12202 10843 12205
rect 15653 12202 15719 12205
rect 10777 12200 15719 12202
rect 10777 12144 10782 12200
rect 10838 12144 15658 12200
rect 15714 12144 15719 12200
rect 10777 12142 15719 12144
rect 10777 12139 10843 12142
rect 15653 12139 15719 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 800 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 800 11734
rect 4061 11731 4127 11734
rect 17401 11794 17467 11797
rect 22000 11794 22800 11824
rect 17401 11792 22800 11794
rect 17401 11736 17406 11792
rect 17462 11736 22800 11792
rect 17401 11734 22800 11736
rect 17401 11731 17467 11734
rect 22000 11704 22800 11734
rect 8661 11658 8727 11661
rect 1948 11656 8727 11658
rect 1948 11600 8666 11656
rect 8722 11600 8727 11656
rect 1948 11598 8727 11600
rect 0 11386 800 11416
rect 1948 11386 2008 11598
rect 8661 11595 8727 11598
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 0 11326 2008 11386
rect 18689 11386 18755 11389
rect 22000 11386 22800 11416
rect 18689 11384 22800 11386
rect 18689 11328 18694 11384
rect 18750 11328 22800 11384
rect 18689 11326 22800 11328
rect 0 11296 800 11326
rect 18689 11323 18755 11326
rect 22000 11296 22800 11326
rect 19609 11114 19675 11117
rect 19742 11114 19748 11116
rect 19609 11112 19748 11114
rect 19609 11056 19614 11112
rect 19670 11056 19748 11112
rect 19609 11054 19748 11056
rect 19609 11051 19675 11054
rect 19742 11052 19748 11054
rect 19812 11052 19818 11116
rect 4376 10912 4696 10913
rect 0 10842 800 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 800 10782
rect 4061 10779 4127 10782
rect 20345 10842 20411 10845
rect 22000 10842 22800 10872
rect 20345 10840 22800 10842
rect 20345 10784 20350 10840
rect 20406 10784 22800 10840
rect 20345 10782 22800 10784
rect 20345 10779 20411 10782
rect 22000 10752 22800 10782
rect 9857 10706 9923 10709
rect 17401 10706 17467 10709
rect 9857 10704 17467 10706
rect 9857 10648 9862 10704
rect 9918 10648 17406 10704
rect 17462 10648 17467 10704
rect 9857 10646 17467 10648
rect 9857 10643 9923 10646
rect 17401 10643 17467 10646
rect 18505 10706 18571 10709
rect 18822 10706 18828 10708
rect 18505 10704 18828 10706
rect 18505 10648 18510 10704
rect 18566 10648 18828 10704
rect 18505 10646 18828 10648
rect 18505 10643 18571 10646
rect 18822 10644 18828 10646
rect 18892 10644 18898 10708
rect 0 10434 800 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 800 10374
rect 4061 10371 4127 10374
rect 17953 10434 18019 10437
rect 22000 10434 22800 10464
rect 17953 10432 22800 10434
rect 17953 10376 17958 10432
rect 18014 10376 22800 10432
rect 17953 10374 22800 10376
rect 17953 10371 18019 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22000 10344 22800 10374
rect 14672 10303 14992 10304
rect 0 10026 800 10056
rect 3969 10026 4035 10029
rect 0 10024 4035 10026
rect 0 9968 3974 10024
rect 4030 9968 4035 10024
rect 0 9966 4035 9968
rect 0 9936 800 9966
rect 3969 9963 4035 9966
rect 17953 10026 18019 10029
rect 22000 10026 22800 10056
rect 17953 10024 22800 10026
rect 17953 9968 17958 10024
rect 18014 9968 22800 10024
rect 17953 9966 22800 9968
rect 17953 9963 18019 9966
rect 22000 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 0 9482 800 9512
rect 4061 9482 4127 9485
rect 0 9480 4127 9482
rect 0 9424 4066 9480
rect 4122 9424 4127 9480
rect 0 9422 4127 9424
rect 0 9392 800 9422
rect 4061 9419 4127 9422
rect 5349 9482 5415 9485
rect 7833 9482 7899 9485
rect 5349 9480 7899 9482
rect 5349 9424 5354 9480
rect 5410 9424 7838 9480
rect 7894 9424 7899 9480
rect 5349 9422 7899 9424
rect 5349 9419 5415 9422
rect 7833 9419 7899 9422
rect 12249 9482 12315 9485
rect 13445 9482 13511 9485
rect 12249 9480 13511 9482
rect 12249 9424 12254 9480
rect 12310 9424 13450 9480
rect 13506 9424 13511 9480
rect 12249 9422 13511 9424
rect 12249 9419 12315 9422
rect 13445 9419 13511 9422
rect 14273 9482 14339 9485
rect 22000 9482 22800 9512
rect 14273 9480 22800 9482
rect 14273 9424 14278 9480
rect 14334 9424 22800 9480
rect 14273 9422 22800 9424
rect 14273 9419 14339 9422
rect 22000 9392 22800 9422
rect 9857 9346 9923 9349
rect 9990 9346 9996 9348
rect 9857 9344 9996 9346
rect 9857 9288 9862 9344
rect 9918 9288 9996 9344
rect 9857 9286 9996 9288
rect 9857 9283 9923 9286
rect 9990 9284 9996 9286
rect 10060 9346 10066 9348
rect 12985 9346 13051 9349
rect 17677 9348 17743 9349
rect 17677 9346 17724 9348
rect 10060 9344 13051 9346
rect 10060 9288 12990 9344
rect 13046 9288 13051 9344
rect 10060 9286 13051 9288
rect 17632 9344 17724 9346
rect 17632 9288 17682 9344
rect 17632 9286 17724 9288
rect 10060 9284 10066 9286
rect 12985 9283 13051 9286
rect 17677 9284 17724 9286
rect 17788 9284 17794 9348
rect 17677 9283 17743 9284
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 19149 9074 19215 9077
rect 22000 9074 22800 9104
rect 19149 9072 22800 9074
rect 19149 9016 19154 9072
rect 19210 9016 22800 9072
rect 19149 9014 22800 9016
rect 19149 9011 19215 9014
rect 22000 8984 22800 9014
rect 2957 8938 3023 8941
rect 4705 8938 4771 8941
rect 9305 8938 9371 8941
rect 2957 8936 9371 8938
rect 2957 8880 2962 8936
rect 3018 8880 4710 8936
rect 4766 8880 9310 8936
rect 9366 8880 9371 8936
rect 2957 8878 9371 8880
rect 2957 8875 3023 8878
rect 4705 8875 4771 8878
rect 9305 8875 9371 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 800 8560
rect 7925 8530 7991 8533
rect 0 8528 7991 8530
rect 0 8472 7930 8528
rect 7986 8472 7991 8528
rect 0 8470 7991 8472
rect 0 8440 800 8470
rect 7925 8467 7991 8470
rect 10317 8530 10383 8533
rect 22000 8530 22800 8560
rect 10317 8528 22800 8530
rect 10317 8472 10322 8528
rect 10378 8472 22800 8528
rect 10317 8470 22800 8472
rect 10317 8467 10383 8470
rect 22000 8440 22800 8470
rect 2405 8394 2471 8397
rect 8385 8394 8451 8397
rect 2405 8392 8451 8394
rect 2405 8336 2410 8392
rect 2466 8336 8390 8392
rect 8446 8336 8451 8392
rect 2405 8334 8451 8336
rect 2405 8331 2471 8334
rect 8385 8331 8451 8334
rect 7808 8192 8128 8193
rect 0 8122 800 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 4705 8122 4771 8125
rect 0 8120 4771 8122
rect 0 8064 4710 8120
rect 4766 8064 4771 8120
rect 0 8062 4771 8064
rect 0 8032 800 8062
rect 4705 8059 4771 8062
rect 18045 8122 18111 8125
rect 22000 8122 22800 8152
rect 18045 8120 22800 8122
rect 18045 8064 18050 8120
rect 18106 8064 22800 8120
rect 18045 8062 22800 8064
rect 18045 8059 18111 8062
rect 22000 8032 22800 8062
rect 11973 7986 12039 7989
rect 9814 7984 12039 7986
rect 9814 7928 11978 7984
rect 12034 7928 12039 7984
rect 9814 7926 12039 7928
rect 9814 7853 9874 7926
rect 11973 7923 12039 7926
rect 13261 7986 13327 7989
rect 15929 7986 15995 7989
rect 13261 7984 15995 7986
rect 13261 7928 13266 7984
rect 13322 7928 15934 7984
rect 15990 7928 15995 7984
rect 13261 7926 15995 7928
rect 13261 7923 13327 7926
rect 15929 7923 15995 7926
rect 9765 7848 9874 7853
rect 9765 7792 9770 7848
rect 9826 7792 9874 7848
rect 9765 7790 9874 7792
rect 9765 7787 9831 7790
rect 11973 7714 12039 7717
rect 15469 7714 15535 7717
rect 11973 7712 15535 7714
rect 11973 7656 11978 7712
rect 12034 7656 15474 7712
rect 15530 7656 15535 7712
rect 11973 7654 15535 7656
rect 11973 7651 12039 7654
rect 15469 7651 15535 7654
rect 4376 7648 4696 7649
rect 0 7578 800 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 18505 7578 18571 7581
rect 22000 7578 22800 7608
rect 0 7518 4170 7578
rect 0 7488 800 7518
rect 4110 7442 4170 7518
rect 18505 7576 22800 7578
rect 18505 7520 18510 7576
rect 18566 7520 22800 7576
rect 18505 7518 22800 7520
rect 18505 7515 18571 7518
rect 22000 7488 22800 7518
rect 8753 7442 8819 7445
rect 4110 7440 8819 7442
rect 4110 7384 8758 7440
rect 8814 7384 8819 7440
rect 4110 7382 8819 7384
rect 8753 7379 8819 7382
rect 9765 7306 9831 7309
rect 11605 7306 11671 7309
rect 9765 7304 11671 7306
rect 9765 7248 9770 7304
rect 9826 7248 11610 7304
rect 11666 7248 11671 7304
rect 9765 7246 11671 7248
rect 9765 7243 9831 7246
rect 11605 7243 11671 7246
rect 12709 7306 12775 7309
rect 13905 7306 13971 7309
rect 12709 7304 13971 7306
rect 12709 7248 12714 7304
rect 12770 7248 13910 7304
rect 13966 7248 13971 7304
rect 12709 7246 13971 7248
rect 12709 7243 12775 7246
rect 13905 7243 13971 7246
rect 0 7170 800 7200
rect 2037 7170 2103 7173
rect 0 7168 2103 7170
rect 0 7112 2042 7168
rect 2098 7112 2103 7168
rect 0 7110 2103 7112
rect 0 7080 800 7110
rect 2037 7107 2103 7110
rect 19977 7170 20043 7173
rect 22000 7170 22800 7200
rect 19977 7168 22800 7170
rect 19977 7112 19982 7168
rect 20038 7112 22800 7168
rect 19977 7110 22800 7112
rect 19977 7107 20043 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22000 7080 22800 7110
rect 14672 7039 14992 7040
rect 18689 6900 18755 6901
rect 18638 6836 18644 6900
rect 18708 6898 18755 6900
rect 18708 6896 18800 6898
rect 18750 6840 18800 6896
rect 18708 6838 18800 6840
rect 18708 6836 18755 6838
rect 18689 6835 18755 6836
rect 0 6762 800 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 800 6702
rect 4061 6699 4127 6702
rect 17953 6762 18019 6765
rect 22000 6762 22800 6792
rect 17953 6760 22800 6762
rect 17953 6704 17958 6760
rect 18014 6704 22800 6760
rect 17953 6702 22800 6704
rect 17953 6699 18019 6702
rect 22000 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 9857 6354 9923 6357
rect 12525 6354 12591 6357
rect 9857 6352 12591 6354
rect 9857 6296 9862 6352
rect 9918 6296 12530 6352
rect 12586 6296 12591 6352
rect 9857 6294 12591 6296
rect 9857 6291 9923 6294
rect 12525 6291 12591 6294
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 22000 6218 22800 6248
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 14414 6158 22800 6218
rect 9121 6082 9187 6085
rect 14414 6082 14474 6158
rect 22000 6128 22800 6158
rect 9121 6080 14474 6082
rect 9121 6024 9126 6080
rect 9182 6024 14474 6080
rect 9121 6022 14474 6024
rect 18413 6082 18479 6085
rect 18638 6082 18644 6084
rect 18413 6080 18644 6082
rect 18413 6024 18418 6080
rect 18474 6024 18644 6080
rect 18413 6022 18644 6024
rect 9121 6019 9187 6022
rect 18413 6019 18479 6022
rect 18638 6020 18644 6022
rect 18708 6020 18714 6084
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 9857 5946 9923 5949
rect 14365 5946 14431 5949
rect 9857 5944 14431 5946
rect 9857 5888 9862 5944
rect 9918 5888 14370 5944
rect 14426 5888 14431 5944
rect 9857 5886 14431 5888
rect 9857 5883 9923 5886
rect 14365 5883 14431 5886
rect 0 5810 800 5840
rect 3969 5810 4035 5813
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 0 5720 800 5750
rect 3969 5747 4035 5750
rect 18505 5810 18571 5813
rect 22000 5810 22800 5840
rect 18505 5808 22800 5810
rect 18505 5752 18510 5808
rect 18566 5752 22800 5808
rect 18505 5750 22800 5752
rect 18505 5747 18571 5750
rect 22000 5720 22800 5750
rect 9765 5674 9831 5677
rect 12065 5674 12131 5677
rect 9765 5672 12131 5674
rect 9765 5616 9770 5672
rect 9826 5616 12070 5672
rect 12126 5616 12131 5672
rect 9765 5614 12131 5616
rect 9765 5611 9831 5614
rect 12065 5611 12131 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 800 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 800 5206
rect 3969 5203 4035 5206
rect 20621 5266 20687 5269
rect 22000 5266 22800 5296
rect 20621 5264 22800 5266
rect 20621 5208 20626 5264
rect 20682 5208 22800 5264
rect 20621 5206 22800 5208
rect 20621 5203 20687 5206
rect 22000 5176 22800 5206
rect 7808 4928 8128 4929
rect 0 4858 800 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 6177 4858 6243 4861
rect 0 4856 6243 4858
rect 0 4800 6182 4856
rect 6238 4800 6243 4856
rect 0 4798 6243 4800
rect 0 4768 800 4798
rect 6177 4795 6243 4798
rect 15101 4858 15167 4861
rect 22000 4858 22800 4888
rect 15101 4856 22800 4858
rect 15101 4800 15106 4856
rect 15162 4800 22800 4856
rect 15101 4798 22800 4800
rect 15101 4795 15167 4798
rect 22000 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 800 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 9673 4314 9739 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 800 4254
rect 4061 4251 4127 4254
rect 9630 4312 9739 4314
rect 9630 4256 9678 4312
rect 9734 4256 9739 4312
rect 9630 4251 9739 4256
rect 20529 4314 20595 4317
rect 22000 4314 22800 4344
rect 20529 4312 22800 4314
rect 20529 4256 20534 4312
rect 20590 4256 22800 4312
rect 20529 4254 22800 4256
rect 20529 4251 20595 4254
rect 0 3906 800 3936
rect 9630 3909 9690 4251
rect 22000 4224 22800 4254
rect 0 3846 4906 3906
rect 9630 3904 9739 3909
rect 9630 3848 9678 3904
rect 9734 3848 9739 3904
rect 9630 3846 9739 3848
rect 0 3816 800 3846
rect 4846 3634 4906 3846
rect 9673 3843 9739 3846
rect 18965 3906 19031 3909
rect 22000 3906 22800 3936
rect 18965 3904 22800 3906
rect 18965 3848 18970 3904
rect 19026 3848 22800 3904
rect 18965 3846 22800 3848
rect 18965 3843 19031 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22000 3816 22800 3846
rect 14672 3775 14992 3776
rect 8845 3634 8911 3637
rect 4846 3632 8911 3634
rect 4846 3576 8850 3632
rect 8906 3576 8911 3632
rect 4846 3574 8911 3576
rect 8845 3571 8911 3574
rect 0 3498 800 3528
rect 2773 3498 2839 3501
rect 0 3496 2839 3498
rect 0 3440 2778 3496
rect 2834 3440 2839 3496
rect 0 3438 2839 3440
rect 0 3408 800 3438
rect 2773 3435 2839 3438
rect 16021 3498 16087 3501
rect 22000 3498 22800 3528
rect 16021 3496 22800 3498
rect 16021 3440 16026 3496
rect 16082 3440 22800 3496
rect 16021 3438 22800 3440
rect 16021 3435 16087 3438
rect 22000 3408 22800 3438
rect 9949 3364 10015 3365
rect 9949 3360 9996 3364
rect 10060 3362 10066 3364
rect 9949 3304 9954 3360
rect 9949 3300 9996 3304
rect 10060 3302 10106 3362
rect 10060 3300 10066 3302
rect 9949 3299 10015 3300
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 800 2984
rect 5073 2954 5139 2957
rect 0 2952 5139 2954
rect 0 2896 5078 2952
rect 5134 2896 5139 2952
rect 0 2894 5139 2896
rect 0 2864 800 2894
rect 5073 2891 5139 2894
rect 18638 2892 18644 2956
rect 18708 2954 18714 2956
rect 22000 2954 22800 2984
rect 18708 2894 22800 2954
rect 18708 2892 18714 2894
rect 22000 2864 22800 2894
rect 1945 2818 2011 2821
rect 2957 2818 3023 2821
rect 1945 2816 3023 2818
rect 1945 2760 1950 2816
rect 2006 2760 2962 2816
rect 3018 2760 3023 2816
rect 1945 2758 3023 2760
rect 1945 2755 2011 2758
rect 2957 2755 3023 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 800 2576
rect 3141 2546 3207 2549
rect 0 2544 3207 2546
rect 0 2488 3146 2544
rect 3202 2488 3207 2544
rect 0 2486 3207 2488
rect 0 2456 800 2486
rect 3141 2483 3207 2486
rect 17718 2484 17724 2548
rect 17788 2546 17794 2548
rect 22000 2546 22800 2576
rect 17788 2486 22800 2546
rect 17788 2484 17794 2486
rect 22000 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 800 2032
rect 3601 2002 3667 2005
rect 0 2000 3667 2002
rect 0 1944 3606 2000
rect 3662 1944 3667 2000
rect 0 1942 3667 1944
rect 0 1912 800 1942
rect 3601 1939 3667 1942
rect 17769 2002 17835 2005
rect 22000 2002 22800 2032
rect 17769 2000 22800 2002
rect 17769 1944 17774 2000
rect 17830 1944 22800 2000
rect 17769 1942 22800 1944
rect 17769 1939 17835 1942
rect 22000 1912 22800 1942
rect 0 1594 800 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 800 1534
rect 2865 1531 2931 1534
rect 19057 1594 19123 1597
rect 22000 1594 22800 1624
rect 19057 1592 22800 1594
rect 19057 1536 19062 1592
rect 19118 1536 22800 1592
rect 19057 1534 22800 1536
rect 19057 1531 19123 1534
rect 22000 1504 22800 1534
rect 0 1050 800 1080
rect 3233 1050 3299 1053
rect 0 1048 3299 1050
rect 0 992 3238 1048
rect 3294 992 3299 1048
rect 0 990 3299 992
rect 0 960 800 990
rect 3233 987 3299 990
rect 19701 1050 19767 1053
rect 22000 1050 22800 1080
rect 19701 1048 22800 1050
rect 19701 992 19706 1048
rect 19762 992 22800 1048
rect 19701 990 22800 992
rect 19701 987 19767 990
rect 22000 960 22800 990
rect 0 642 800 672
rect 4061 642 4127 645
rect 0 640 4127 642
rect 0 584 4066 640
rect 4122 584 4127 640
rect 0 582 4127 584
rect 0 552 800 582
rect 4061 579 4127 582
rect 19241 642 19307 645
rect 22000 642 22800 672
rect 19241 640 22800 642
rect 19241 584 19246 640
rect 19302 584 22800 640
rect 19241 582 22800 584
rect 19241 579 19307 582
rect 22000 552 22800 582
rect 0 234 800 264
rect 6269 234 6335 237
rect 0 232 6335 234
rect 0 176 6274 232
rect 6330 176 6335 232
rect 0 174 6335 176
rect 0 144 800 174
rect 6269 171 6335 174
rect 17493 234 17559 237
rect 22000 234 22800 264
rect 17493 232 22800 234
rect 17493 176 17498 232
rect 17554 176 22800 232
rect 17493 174 22800 176
rect 17493 171 17559 174
rect 22000 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 19748 18260 19812 18324
rect 19380 17988 19444 18052
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 19012 17776 19076 17780
rect 19012 17720 19062 17776
rect 19062 17720 19076 17776
rect 19012 17716 19076 17720
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 19012 16492 19076 16556
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 18828 14044 18892 14108
rect 19380 13772 19444 13836
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 19012 13152 19076 13156
rect 19012 13096 19026 13152
rect 19026 13096 19076 13152
rect 19012 13092 19076 13096
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 19748 11052 19812 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 18828 10644 18892 10708
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 9996 9284 10060 9348
rect 17724 9344 17788 9348
rect 17724 9288 17738 9344
rect 17738 9288 17788 9344
rect 17724 9284 17788 9288
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 18644 6896 18708 6900
rect 18644 6840 18694 6896
rect 18694 6840 18708 6896
rect 18644 6836 18708 6840
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 18644 6020 18708 6084
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 9996 3360 10060 3364
rect 9996 3304 10010 3360
rect 10010 3304 10060 3360
rect 9996 3300 10060 3304
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 18644 2892 18708 2956
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 17724 2484 17788 2548
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 9998 3365 10058 9283
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 9995 3364 10061 3365
rect 9995 3300 9996 3364
rect 10060 3300 10061 3364
rect 9995 3299 10061 3300
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 19747 18324 19813 18325
rect 19747 18260 19748 18324
rect 19812 18260 19813 18324
rect 19747 18259 19813 18260
rect 19379 18052 19445 18053
rect 19379 17988 19380 18052
rect 19444 17988 19445 18052
rect 19379 17987 19445 17988
rect 19011 17780 19077 17781
rect 19011 17716 19012 17780
rect 19076 17716 19077 17780
rect 19011 17715 19077 17716
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 19014 16557 19074 17715
rect 19011 16556 19077 16557
rect 19011 16492 19012 16556
rect 19076 16492 19077 16556
rect 19011 16491 19077 16492
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18827 14108 18893 14109
rect 18827 14044 18828 14108
rect 18892 14044 18893 14108
rect 18827 14043 18893 14044
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18830 10709 18890 14043
rect 19014 13157 19074 16491
rect 19382 13837 19442 17987
rect 19379 13836 19445 13837
rect 19379 13772 19380 13836
rect 19444 13772 19445 13836
rect 19379 13771 19445 13772
rect 19011 13156 19077 13157
rect 19011 13092 19012 13156
rect 19076 13092 19077 13156
rect 19011 13091 19077 13092
rect 19750 11117 19810 18259
rect 19747 11116 19813 11117
rect 19747 11052 19748 11116
rect 19812 11052 19813 11116
rect 19747 11051 19813 11052
rect 18827 10708 18893 10709
rect 18827 10644 18828 10708
rect 18892 10644 18893 10708
rect 18827 10643 18893 10644
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 17723 9348 17789 9349
rect 17723 9284 17724 9348
rect 17788 9284 17789 9348
rect 17723 9283 17789 9284
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 17726 2549 17786 9283
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18643 6900 18709 6901
rect 18643 6836 18644 6900
rect 18708 6836 18709 6900
rect 18643 6835 18709 6836
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18646 6085 18706 6835
rect 18643 6084 18709 6085
rect 18643 6020 18644 6084
rect 18708 6020 18709 6084
rect 18643 6019 18709 6020
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 17723 2548 17789 2549
rect 17723 2484 17724 2548
rect 17788 2484 17789 2548
rect 17723 2483 17789 2484
rect 18104 2208 18424 3232
rect 18646 2957 18706 6019
rect 18643 2956 18709 2957
rect 18643 2892 18644 2956
rect 18708 2892 18709 2956
rect 18643 2891 18709 2892
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608762747
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608762747
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608762747
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1608762747
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1608762747
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608762747
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608762747
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608762747
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1608762747
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608762747
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp 1608762747
transform 1 0 17388 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1608762747
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1608762747
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1608762747
transform 1 0 15456 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608762747
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1608762747
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1608762747
transform 1 0 16284 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1608762747
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608762747
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608762747
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608762747
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1608762747
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608762747
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1608762747
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608762747
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1608762747
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1608762747
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608762747
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608762747
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1608762747
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608762747
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608762747
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608762747
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608762747
transform 1 0 1840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608762747
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608762747
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1608762747
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1608762747
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1608762747
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_18
timestamp 1608762747
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608762747
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608762747
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1608762747
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1608762747
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1608762747
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608762747
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608762747
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608762747
transform 1 0 18860 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1608762747
transform 1 0 18768 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1608762747
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1608762747
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608762747
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_173
timestamp 1608762747
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1608762747
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1608762747
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_161
timestamp 1608762747
transform 1 0 15916 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 14444 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_139
timestamp 1608762747
transform 1 0 13892 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608762747
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_114
timestamp 1608762747
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 10120 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1608762747
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 8464 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1608762747
transform 1 0 7084 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1608762747
transform 1 0 7912 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608762747
transform 1 0 5152 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 5704 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608762747
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1608762747
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1608762747
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1608762747
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1608762747
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 3128 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_38
timestamp 1608762747
transform 1 0 4600 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608762747
transform 1 0 1840 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608762747
transform 1 0 2392 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608762747
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1608762747
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1608762747
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_12
timestamp 1608762747
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1608762747
transform 1 0 2760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608762747
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608762747
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1608762747
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608762747
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608762747
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608762747
transform 1 0 19320 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 19872 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_195
timestamp 1608762747
transform 1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1608762747
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_175
timestamp 1608762747
transform 1 0 17204 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1608762747
transform 1 0 18308 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 15732 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608762747
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1608762747
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1608762747
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_158
timestamp 1608762747
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1608762747
transform 1 0 13064 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1608762747
transform 1 0 14076 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1608762747
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_139
timestamp 1608762747
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608762747
transform 1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 10948 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1608762747
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1608762747
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608762747
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1608762747
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1608762747
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608762747
transform 1 0 8372 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_76
timestamp 1608762747
transform 1 0 8096 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 6624 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1608762747
transform 1 0 6164 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1608762747
transform 1 0 6532 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 4692 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608762747
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1608762747
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_32
timestamp 1608762747
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1608762747
transform 1 0 4600 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608762747
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608762747
transform 1 0 2300 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608762747
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608762747
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1608762747
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1608762747
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1608762747
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608762747
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608762747
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1608762747
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1608762747
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1608762747
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608762747
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608762747
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1608762747
transform 1 0 18768 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_200
timestamp 1608762747
transform 1 0 19504 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1608762747
transform 1 0 19872 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 18216 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608762747
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1608762747
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1608762747
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1608762747
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608762747
transform 1 0 16100 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15088 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_149
timestamp 1608762747
transform 1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1608762747
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608762747
transform 1 0 13248 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1608762747
transform 1 0 13156 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_141
timestamp 1608762747
transform 1 0 14076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608762747
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_109
timestamp 1608762747
transform 1 0 11132 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1608762747
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1608762747
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1608762747
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1608762747
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608762747
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 8648 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1608762747
transform 1 0 6992 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_73
timestamp 1608762747
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_78
timestamp 1608762747
transform 1 0 8280 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608762747
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1608762747
transform 1 0 5060 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_55
timestamp 1608762747
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1608762747
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 3588 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1608762747
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608762747
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1608762747
transform 1 0 2576 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608762747
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608762747
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1608762747
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1608762747
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608762747
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608762747
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608762747
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608762747
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_196
timestamp 1608762747
transform 1 0 19136 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1608762747
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 16560 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_167
timestamp 1608762747
transform 1 0 16468 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1608762747
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608762747
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608762747
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1608762747
transform 1 0 16100 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608762747
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_128
timestamp 1608762747
transform 1 0 12880 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1608762747
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1608762747
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1608762747
transform 1 0 11592 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1608762747
transform 1 0 11960 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608762747
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608762747
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1608762747
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1608762747
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1608762747
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_78
timestamp 1608762747
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 6624 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1608762747
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1608762747
transform 1 0 6256 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608762747
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608762747
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1608762747
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1608762747
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608762747
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1608762747
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1608762747
transform 1 0 1932 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608762747
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1608762747
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1608762747
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608762747
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608762747
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608762747
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1608762747
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608762747
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608762747
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1608762747
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608762747
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1608762747
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1608762747
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608762747
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608762747
transform 1 0 19688 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608762747
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_198
timestamp 1608762747
transform 1 0 19320 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1608762747
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1608762747
transform 1 0 19596 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 18124 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608762747
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_174
timestamp 1608762747
transform 1 0 17112 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1608762747
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1608762747
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1608762747
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608762747
transform 1 0 16008 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608762747
transform 1 0 16284 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608762747
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1608762747
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1608762747
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1608762747
transform 1 0 15272 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 12696 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608762747
transform 1 0 13340 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_142
timestamp 1608762747
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp 1608762747
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_142
timestamp 1608762747
transform 1 0 14168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1608762747
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608762747
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_105
timestamp 1608762747
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_122
timestamp 1608762747
transform 1 0 12328 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608762747
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_123
timestamp 1608762747
transform 1 0 12420 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 10672 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608762747
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1608762747
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1608762747
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1608762747
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_84
timestamp 1608762747
transform 1 0 8832 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_96
timestamp 1608762747
transform 1 0 9936 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 7636 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1608762747
transform 1 0 8004 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1608762747
transform 1 0 7636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 5060 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1608762747
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608762747
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_59
timestamp 1608762747
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_49
timestamp 1608762747
transform 1 0 5612 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608762747
transform 1 0 4784 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608762747
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1608762747
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_40
timestamp 1608762747
transform 1 0 4784 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1608762747
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608762747
transform 1 0 3404 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1608762747
transform 1 0 3036 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1608762747
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1608762747
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_30
timestamp 1608762747
transform 1 0 3864 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608762747
transform 1 0 2852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1608762747
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_16
timestamp 1608762747
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_20
timestamp 1608762747
transform 1 0 2944 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1608762747
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1608762747
transform 1 0 2300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1608762747
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1608762747
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1608762747
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608762747
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608762747
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608762747
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1608762747
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 20516 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608762747
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1608762747
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1608762747
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 19780 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_200
timestamp 1608762747
transform 1 0 19504 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608762747
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_167
timestamp 1608762747
transform 1 0 16468 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1608762747
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_155
timestamp 1608762747
transform 1 0 15364 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 13892 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_126
timestamp 1608762747
transform 1 0 12696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_138
timestamp 1608762747
transform 1 0 13800 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608762747
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1608762747
transform 1 0 11316 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608762747
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1608762747
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608762747
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608762747
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1608762747
transform 1 0 9936 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 8464 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1608762747
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_79
timestamp 1608762747
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608762747
transform 1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608762747
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608762747
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608762747
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608762747
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_28
timestamp 1608762747
transform 1 0 3680 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1608762747
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608762747
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1608762747
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1608762747
transform 1 0 1932 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_16
timestamp 1608762747
transform 1 0 2576 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608762747
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608762747
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608762747
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608762747
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608762747
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608762747
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1608762747
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_195
timestamp 1608762747
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1608762747
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1608762747
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_176
timestamp 1608762747
transform 1 0 17296 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_184
timestamp 1608762747
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 15824 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608762747
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608762747
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_154
timestamp 1608762747
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1608762747
transform 1 0 13432 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_133
timestamp 1608762747
transform 1 0 13340 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_143
timestamp 1608762747
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1608762747
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1608762747
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1608762747
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608762747
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608762747
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608762747
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1608762747
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608762747
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 7820 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_67
timestamp 1608762747
transform 1 0 7268 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_76
timestamp 1608762747
transform 1 0 8096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1608762747
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_48
timestamp 1608762747
transform 1 0 5520 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 4048 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608762747
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1608762747
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1608762747
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 2300 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608762747
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1608762747
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1608762747
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608762747
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608762747
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1608762747
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1608762747
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608762747
transform 1 0 18400 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1608762747
transform 1 0 18860 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 19964 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1608762747
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_202
timestamp 1608762747
transform 1 0 19688 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1608762747
transform 1 0 16928 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608762747
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_168
timestamp 1608762747
transform 1 0 16560 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608762747
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1608762747
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 15088 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1608762747
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 13432 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_23_128
timestamp 1608762747
transform 1 0 12880 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608762747
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 12604 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1608762747
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1608762747
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1608762747
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_91
timestamp 1608762747
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_103
timestamp 1608762747
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 6992 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1608762747
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1608762747
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608762747
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1608762747
transform 1 0 4968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_54
timestamp 1608762747
transform 1 0 6072 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608762747
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1608762747
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 3496 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_23
timestamp 1608762747
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1608762747
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608762747
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1608762747
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_11
timestamp 1608762747
transform 1 0 2116 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608762747
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608762747
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608762747
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608762747
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608762747
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608762747
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608762747
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_194
timestamp 1608762747
transform 1 0 18952 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1608762747
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608762747
transform 1 0 18124 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608762747
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1608762747
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608762747
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_148
timestamp 1608762747
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1608762747
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_166
timestamp 1608762747
transform 1 0 16376 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1608762747
transform 1 0 13892 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1608762747
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 12236 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1608762747
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1608762747
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608762747
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1608762747
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608762747
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1608762747
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1608762747
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1608762747
transform 1 0 6992 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_73
timestamp 1608762747
transform 1 0 7820 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 5336 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp 1608762747
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_62
timestamp 1608762747
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608762747
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_25
timestamp 1608762747
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608762747
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1608762747
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1608762747
transform 1 0 2576 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608762747
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608762747
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1608762747
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1608762747
transform 1 0 2484 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608762747
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608762747
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1608762747
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1608762747
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 20056 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608762747
transform 1 0 18768 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1608762747
transform 1 0 19596 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_205
timestamp 1608762747
transform 1 0 19964 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608762747
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_170
timestamp 1608762747
transform 1 0 16744 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608762747
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_184
timestamp 1608762747
transform 1 0 18032 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_152
timestamp 1608762747
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1608762747
transform 1 0 13248 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1608762747
transform 1 0 14260 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1608762747
transform 1 0 13156 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1608762747
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1608762747
transform 1 0 11224 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608762747
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_107
timestamp 1608762747
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1608762747
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1608762747
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608762747
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1608762747
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1608762747
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1608762747
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1608762747
transform 1 0 8096 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1608762747
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1608762747
transform 1 0 8004 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608762747
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608762747
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 5980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1608762747
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_56
timestamp 1608762747
transform 1 0 6256 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608762747
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1608762747
transform 1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608762747
transform 1 0 3864 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_26
timestamp 1608762747
transform 1 0 3496 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608762747
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1608762747
transform 1 0 2116 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608762747
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1608762747
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1608762747
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608762747
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608762747
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608762747
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1608762747
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608762747
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608762747
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608762747
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608762747
transform 1 0 20240 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608762747
transform 1 0 18676 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1608762747
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1608762747
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_200
timestamp 1608762747
transform 1 0 19504 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608762747
transform 1 0 16468 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608762747
transform 1 0 16468 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608762747
transform 1 0 18308 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608762747
transform 1 0 17664 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608762747
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_176
timestamp 1608762747
transform 1 0 17296 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1608762747
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1608762747
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1608762747
transform 1 0 17296 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1608762747
transform 1 0 15272 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608762747
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1608762747
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1608762747
transform 1 0 16100 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1608762747
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_165
timestamp 1608762747
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608762747
transform 1 0 13800 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608762747
transform 1 0 12788 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1608762747
transform 1 0 14260 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 13616 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1608762747
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1608762747
transform 1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1608762747
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608762747
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608762747
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1608762747
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608762747
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_108
timestamp 1608762747
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1608762747
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608762747
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_117
timestamp 1608762747
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1608762747
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608762747
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608762747
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_88
timestamp 1608762747
transform 1 0 9200 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_100
timestamp 1608762747
transform 1 0 10304 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1608762747
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1608762747
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608762747
transform 1 0 7268 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1608762747
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1608762747
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 7084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1608762747
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1608762747
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_76
timestamp 1608762747
transform 1 0 8096 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608762747
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608762747
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608762747
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608762747
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1608762747
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_46
timestamp 1608762747
transform 1 0 5336 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1608762747
transform 1 0 6440 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_23
timestamp 1608762747
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608762747
transform 1 0 4508 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1608762747
transform 1 0 4324 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_41
timestamp 1608762747
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608762747
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1608762747
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608762747
transform 1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608762747
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1608762747
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1608762747
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608762747
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1608762747
transform 1 0 2392 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1608762747
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608762747
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608762747
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1608762747
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1608762747
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1608762747
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1608762747
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608762747
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608762747
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608762747
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608762747
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608762747
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 19136 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1608762747
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608762747
transform 1 0 18124 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_175
timestamp 1608762747
transform 1 0 17204 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1608762747
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1608762747
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608762747
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1608762747
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_163
timestamp 1608762747
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 13156 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1608762747
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1608762747
transform 1 0 11132 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1608762747
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608762747
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1608762747
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1608762747
transform 1 0 7084 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608762747
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1608762747
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1608762747
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_79
timestamp 1608762747
transform 1 0 8372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608762747
transform 1 0 5796 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1608762747
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_60
timestamp 1608762747
transform 1 0 6624 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608762747
transform 1 0 4784 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608762747
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1608762747
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1608762747
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1608762747
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1608762747
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608762747
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1608762747
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1608762747
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608762747
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_210
timestamp 1608762747
transform 1 0 20424 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1608762747
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 18952 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1608762747
transform 1 0 18860 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608762747
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608762747
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_176
timestamp 1608762747
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1608762747
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_187
timestamp 1608762747
transform 1 0 18308 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608762747
transform 1 0 15364 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1608762747
transform 1 0 14996 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_164
timestamp 1608762747
transform 1 0 16192 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1608762747
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1608762747
transform 1 0 11500 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608762747
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608762747
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_110
timestamp 1608762747
transform 1 0 11224 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608762747
transform 1 0 9844 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_89
timestamp 1608762747
transform 1 0 9292 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_104
timestamp 1608762747
transform 1 0 10672 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1608762747
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608762747
transform 1 0 8464 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_74
timestamp 1608762747
transform 1 0 7912 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608762747
transform 1 0 5520 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608762747
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_44
timestamp 1608762747
transform 1 0 5152 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1608762747
transform 1 0 6348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1608762747
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1608762747
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_29
timestamp 1608762747
transform 1 0 3772 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 2300 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608762747
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1608762747
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1608762747
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608762747
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608762747
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608762747
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608762747
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1608762747
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1608762747
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1608762747
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 17204 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608762747
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608762747
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608762747
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_163
timestamp 1608762747
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 13432 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1608762747
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_137
timestamp 1608762747
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608762747
transform 1 0 12420 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608762747
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 10580 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608762747
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1608762747
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_101
timestamp 1608762747
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_74
timestamp 1608762747
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_78
timestamp 1608762747
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1608762747
transform 1 0 5980 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_49
timestamp 1608762747
transform 1 0 5612 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1608762747
transform 1 0 6808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1608762747
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608762747
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_24
timestamp 1608762747
transform 1 0 3312 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608762747
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_32
timestamp 1608762747
transform 1 0 4048 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1608762747
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1608762747
transform 1 0 2484 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608762747
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1608762747
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1608762747
transform 1 0 2116 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608762747
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_211
timestamp 1608762747
transform 1 0 20516 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1608762747
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608762747
transform 1 0 19688 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_193
timestamp 1608762747
transform 1 0 18860 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_201
timestamp 1608762747
transform 1 0 19596 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1608762747
transform 1 0 16928 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1608762747
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608762747
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_171
timestamp 1608762747
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608762747
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608762747
transform 1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1608762747
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1608762747
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1608762747
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_165
timestamp 1608762747
transform 1 0 16284 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608762747
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1608762747
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_139
timestamp 1608762747
transform 1 0 13892 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608762747
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_115
timestamp 1608762747
transform 1 0 11684 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608762747
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1608762747
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 10212 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_88
timestamp 1608762747
transform 1 0 9200 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_96
timestamp 1608762747
transform 1 0 9936 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608762747
transform 1 0 7820 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1608762747
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_76
timestamp 1608762747
transform 1 0 8096 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1608762747
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608762747
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608762747
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608762747
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 4324 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_24
timestamp 1608762747
transform 1 0 3312 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_32
timestamp 1608762747
transform 1 0 4048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 1748 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1608762747
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608762747
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1608762747
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1608762747
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608762747
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608762747
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608762747
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608762747
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1608762747
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1608762747
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_218
timestamp 1608762747
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 19596 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608762747
transform 1 0 19596 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_196
timestamp 1608762747
transform 1 0 19136 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_200
timestamp 1608762747
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1608762747
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 16836 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608762747
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_167
timestamp 1608762747
transform 1 0 16468 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1608762747
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1608762747
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_187
timestamp 1608762747
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608762747
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608762747
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1608762747
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1608762747
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1608762747
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1608762747
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 13064 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 13984 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 13708 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_133
timestamp 1608762747
transform 1 0 13340 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp 1608762747
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1608762747
transform 1 0 12512 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608762747
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1608762747
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608762747
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1608762747
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1608762747
transform 1 0 10948 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1608762747
transform 1 0 11316 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1608762747
transform 1 0 10672 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 8924 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608762747
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608762747
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608762747
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_84
timestamp 1608762747
transform 1 0 8832 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1608762747
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608762747
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1608762747
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 7268 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608762747
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1608762747
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_78
timestamp 1608762747
transform 1 0 8280 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_65
timestamp 1608762747
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1608762747
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1608762747
transform 1 0 6256 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608762747
transform 1 0 5704 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608762747
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_46
timestamp 1608762747
transform 1 0 5336 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608762747
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1608762747
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_48
timestamp 1608762747
transform 1 0 5520 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608762747
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_34
timestamp 1608762747
transform 1 0 4232 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1608762747
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608762747
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_11
timestamp 1608762747
transform 1 0 2116 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1608762747
transform 1 0 2300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_17
timestamp 1608762747
transform 1 0 2668 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1608762747
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 1748 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608762747
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608762747
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608762747
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1608762747
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608762747
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608762747
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1608762747
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608762747
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608762747
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608762747
transform 1 0 19136 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1608762747
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_205
timestamp 1608762747
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 16836 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1608762747
transform 1 0 16744 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1608762747
transform 1 0 18308 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608762747
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1608762747
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608762747
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1608762747
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1608762747
transform 1 0 16376 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_134
timestamp 1608762747
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1608762747
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608762747
transform 1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_114
timestamp 1608762747
transform 1 0 11592 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_122
timestamp 1608762747
transform 1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608762747
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_86
timestamp 1608762747
transform 1 0 9016 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1608762747
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608762747
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608762747
transform 1 0 8188 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1608762747
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1608762747
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 5520 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1608762747
transform 1 0 5428 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608762747
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608762747
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1608762747
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1608762747
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1608762747
transform 1 0 4876 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 1656 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608762747
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1608762747
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608762747
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_213
timestamp 1608762747
transform 1 0 20700 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1608762747
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 19228 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_193
timestamp 1608762747
transform 1 0 18860 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1608762747
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1608762747
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608762747
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1608762747
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1608762747
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 15640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_151
timestamp 1608762747
transform 1 0 14996 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1608762747
transform 1 0 15548 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_161
timestamp 1608762747
transform 1 0 15916 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1608762747
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608762747
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_116
timestamp 1608762747
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_92
timestamp 1608762747
transform 1 0 9568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1608762747
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 8096 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1608762747
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp 1608762747
transform 1 0 8004 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608762747
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608762747
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_50
timestamp 1608762747
transform 1 0 5704 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1608762747
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 4232 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_22
timestamp 1608762747
transform 1 0 3128 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1608762747
transform 1 0 2300 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608762747
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1608762747
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1608762747
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608762747
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608762747
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1608762747
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608762747
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608762747
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1608762747
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_199
timestamp 1608762747
transform 1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608762747
transform 1 0 18032 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1608762747
transform 1 0 17020 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_170
timestamp 1608762747
transform 1 0 16744 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1608762747
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1608762747
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608762747
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1608762747
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1608762747
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1608762747
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1608762747
transform 1 0 12604 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 12328 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_116
timestamp 1608762747
transform 1 0 11776 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608762747
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608762747
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1608762747
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608762747
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_104
timestamp 1608762747
transform 1 0 10672 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 8096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_69
timestamp 1608762747
transform 1 0 7452 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_75
timestamp 1608762747
transform 1 0 8004 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_79
timestamp 1608762747
transform 1 0 8372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608762747
transform 1 0 6624 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762747
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1608762747
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_52
timestamp 1608762747
transform 1 0 5888 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608762747
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608762747
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1608762747
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1608762747
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1608762747
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1608762747
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608762747
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1608762747
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608762747
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 1608762747
transform 1 0 20792 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 19320 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1608762747
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608762747
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1608762747
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1608762747
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 16192 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_148
timestamp 1608762747
transform 1 0 14720 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1608762747
transform 1 0 15824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608762747
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 13248 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_130
timestamp 1608762747
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608762747
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_109
timestamp 1608762747
transform 1 0 11132 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608762747
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1608762747
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 9660 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1608762747
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608762747
transform 1 0 8648 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_74
timestamp 1608762747
transform 1 0 7912 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1608762747
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608762747
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608762747
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608762747
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1608762747
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1608762747
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 1608762747
transform 1 0 3496 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 1608762747
transform 1 0 4600 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1608762747
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608762747
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1608762747
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1608762747
transform 1 0 2116 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608762747
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608762747
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608762747
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608762747
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608762747
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608762747
transform 1 0 18676 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_188
timestamp 1608762747
transform 1 0 18400 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1608762747
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608762747
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp 1608762747
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_176
timestamp 1608762747
transform 1 0 17296 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608762747
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_133
timestamp 1608762747
transform 1 0 13340 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1608762747
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1608762747
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_119
timestamp 1608762747
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_123
timestamp 1608762747
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 10580 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608762747
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608762747
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1608762747
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1608762747
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1608762747
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_72
timestamp 1608762747
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_82
timestamp 1608762747
transform 1 0 8648 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1608762747
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_44
timestamp 1608762747
transform 1 0 5152 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_50
timestamp 1608762747
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_60
timestamp 1608762747
transform 1 0 6624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608762747
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1608762747
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608762747
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608762747
transform 1 0 1840 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608762747
transform 1 0 2576 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608762747
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1608762747
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1608762747
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1608762747
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_11
timestamp 1608762747
transform 1 0 2116 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608762747
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608762747
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608762747
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1608762747
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1608762747
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608762747
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608762747
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_216
timestamp 1608762747
transform 1 0 20976 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608762747
transform 1 0 20056 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1608762747
transform 1 0 19136 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608762747
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1608762747
transform 1 0 20148 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1608762747
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_202
timestamp 1608762747
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp 1608762747
transform 1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1608762747
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 17204 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1608762747
transform 1 0 16560 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608762747
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608762747
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_169
timestamp 1608762747
transform 1 0 16652 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1608762747
transform 1 0 16468 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_177
timestamp 1608762747
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1608762747
transform 1 0 15088 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608762747
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608762747
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_154
timestamp 1608762747
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_151
timestamp 1608762747
transform 1 0 14996 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1608762747
transform 1 0 15916 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608762747
transform 1 0 13984 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1608762747
transform 1 0 12880 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1608762747
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1608762747
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1608762747
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_137
timestamp 1608762747
transform 1 0 13708 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1608762747
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1608762747
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_143
timestamp 1608762747
transform 1 0 14260 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 11224 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608762747
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_107
timestamp 1608762747
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1608762747
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp 1608762747
transform 1 0 12420 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1608762747
transform 1 0 10120 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1608762747
transform 1 0 10396 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608762747
transform 1 0 9384 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608762747
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1608762747
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1608762747
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1608762747
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_89
timestamp 1608762747
transform 1 0 9292 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1608762747
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 7084 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1608762747
transform 1 0 7452 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1608762747
transform 1 0 8464 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_66
timestamp 1608762747
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_78
timestamp 1608762747
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_81
timestamp 1608762747
transform 1 0 8556 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1608762747
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 5704 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1608762747
transform 1 0 5244 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608762747
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1608762747
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1608762747
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608762747
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1608762747
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608762747
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_21
timestamp 1608762747
transform 1 0 3036 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1608762747
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_33
timestamp 1608762747
transform 1 0 4140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 2668 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1608762747
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608762747
transform 1 0 2208 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608762747
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608762747
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1608762747
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1608762747
transform 1 0 2116 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1608762747
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_14
timestamp 1608762747
transform 1 0 2392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608762747
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608762747
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1608762747
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1608762747
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 18768 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp 1608762747
transform 1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608762747
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_170
timestamp 1608762747
transform 1 0 16744 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1608762747
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1608762747
transform 1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_158
timestamp 1608762747
transform 1 0 15640 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 14168 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1608762747
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608762747
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 12512 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608762747
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_111
timestamp 1608762747
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1608762747
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1608762747
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 9844 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_94
timestamp 1608762747
transform 1 0 9752 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1608762747
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_70
timestamp 1608762747
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1608762747
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608762747
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_46
timestamp 1608762747
transform 1 0 5336 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_58
timestamp 1608762747
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1608762747
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608762747
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1608762747
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_34
timestamp 1608762747
transform 1 0 4232 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608762747
transform 1 0 2392 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608762747
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608762747
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1608762747
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608762747
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608762747
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608762747
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608762747
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608762747
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1608762747
transform 1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 16652 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1608762747
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1608762747
transform 1 0 18124 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608762747
transform 1 0 15364 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608762747
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1608762747
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_154
timestamp 1608762747
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1608762747
transform 1 0 16192 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1608762747
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_128
timestamp 1608762747
transform 1 0 12880 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_138
timestamp 1608762747
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_112
timestamp 1608762747
transform 1 0 11408 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1608762747
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608762747
transform 1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1608762747
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608762747
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1608762747
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1608762747
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1608762747
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608762747
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_63
timestamp 1608762747
transform 1 0 6900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_71
timestamp 1608762747
transform 1 0 7636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1608762747
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1608762747
transform 1 0 4968 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_51
timestamp 1608762747
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608762747
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_22
timestamp 1608762747
transform 1 0 3128 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1608762747
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1608762747
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1608762747
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608762747
transform 1 0 2300 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608762747
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1608762747
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1608762747
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608762747
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608762747
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1608762747
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1608762747
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1608762747
transform 1 0 21252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608762747
transform 1 0 18952 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1608762747
transform 1 0 19504 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1608762747
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_198
timestamp 1608762747
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608762747
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_174
timestamp 1608762747
transform 1 0 17112 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_182
timestamp 1608762747
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1608762747
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 15640 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608762747
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_156
timestamp 1608762747
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608762747
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608762747
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1608762747
transform 1 0 11500 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1608762747
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608762747
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608762747
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1608762747
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_101
timestamp 1608762747
transform 1 0 10396 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608762747
transform 1 0 7544 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1608762747
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1608762747
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608762747
transform 1 0 5060 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608762747
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608762747
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_46
timestamp 1608762747
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1608762747
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1608762747
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1608762747
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_28
timestamp 1608762747
transform 1 0 3680 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_40
timestamp 1608762747
transform 1 0 4784 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 1472 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608762747
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608762747
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_20
timestamp 1608762747
transform 1 0 2944 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608762747
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608762747
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1608762747
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1608762747
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1608762747
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608762747
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608762747
transform 1 0 19228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608762747
transform 1 0 19780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1608762747
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_194
timestamp 1608762747
transform 1 0 18952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1608762747
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_207
timestamp 1608762747
transform 1 0 20148 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608762747
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1608762747
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1608762747
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608762747
transform 1 0 16284 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608762747
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608762747
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1608762747
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1608762747
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 13616 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_129
timestamp 1608762747
transform 1 0 12972 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1608762747
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_142
timestamp 1608762747
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 11684 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 12420 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_108
timestamp 1608762747
transform 1 0 11040 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_114
timestamp 1608762747
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1608762747
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608762747
transform 1 0 10212 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608762747
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_86
timestamp 1608762747
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93
timestamp 1608762747
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 7544 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1608762747
transform 1 0 7452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608762747
transform 1 0 5520 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_46
timestamp 1608762747
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_57
timestamp 1608762747
transform 1 0 6348 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608762747
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608762747
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1608762747
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1608762747
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1608762747
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608762747
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608762747
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608762747
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1608762747
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_19
timestamp 1608762747
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1608762747
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608762747
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608762747
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608762747
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1608762747
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608762747
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_210
timestamp 1608762747
transform 1 0 20424 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1608762747
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1608762747
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608762747
transform 1 0 19688 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 19504 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1608762747
transform 1 0 19596 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1608762747
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1608762747
transform 1 0 20056 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608762747
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 18768 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1608762747
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1608762747
transform 1 0 19228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1608762747
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608762747
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608762747
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1608762747
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608762747
transform 1 0 17388 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608762747
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1608762747
transform 1 0 17756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608762747
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608762747
transform 1 0 16836 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1608762747
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1608762747
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_167
timestamp 1608762747
transform 1 0 16468 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608762747
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 16100 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_160
timestamp 1608762747
transform 1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1608762747
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608762747
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 15364 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608762747
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1608762747
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_154
timestamp 1608762747
transform 1 0 15272 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608762747
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608762747
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1608762747
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1608762747
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608762747
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1608762747
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1608762747
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608762747
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 13800 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1608762747
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_136
timestamp 1608762747
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608762747
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 13064 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1608762747
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_127
timestamp 1608762747
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608762747
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608762747
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 11040 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 11684 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608762747
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608762747
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1608762747
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1608762747
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1608762747
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608762747
transform 1 0 10028 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608762747
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608762747
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_103
timestamp 1608762747
transform 1 0 10580 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1608762747
transform 1 0 9660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762747
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1608762747
transform 1 0 7452 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1608762747
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_74
timestamp 1608762747
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 5152 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608762747
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608762747
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1608762747
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_47
timestamp 1608762747
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608762747
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608762747
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762747
transform 1 0 3956 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608762747
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608762747
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608762747
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp 1608762747
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_21
timestamp 1608762747
transform 1 0 3036 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1608762747
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762747
transform 1 0 2116 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762747
transform 1 0 1564 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608762747
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608762747
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3
timestamp 1608762747
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1608762747
transform 1 0 1380 0 1 2720
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 800 4 SC_IN_BOT
port 1 nsew
rlabel metal2 s 22098 0 22154 800 4 SC_OUT_BOT
port 2 nsew
rlabel metal2 s 202 0 258 800 4 bottom_left_grid_pin_42_
port 3 nsew
rlabel metal2 s 570 0 626 800 4 bottom_left_grid_pin_43_
port 4 nsew
rlabel metal2 s 1030 0 1086 800 4 bottom_left_grid_pin_44_
port 5 nsew
rlabel metal2 s 1490 0 1546 800 4 bottom_left_grid_pin_45_
port 6 nsew
rlabel metal2 s 1950 0 2006 800 4 bottom_left_grid_pin_46_
port 7 nsew
rlabel metal2 s 2410 0 2466 800 4 bottom_left_grid_pin_47_
port 8 nsew
rlabel metal2 s 2870 0 2926 800 4 bottom_left_grid_pin_48_
port 9 nsew
rlabel metal2 s 3330 0 3386 800 4 bottom_left_grid_pin_49_
port 10 nsew
rlabel metal2 s 5722 22000 5778 22800 4 ccff_head
port 11 nsew
rlabel metal2 s 17130 22000 17186 22800 4 ccff_tail
port 12 nsew
rlabel metal3 s 0 3816 800 3936 4 chanx_left_in[0]
port 13 nsew
rlabel metal3 s 0 8440 800 8560 4 chanx_left_in[10]
port 14 nsew
rlabel metal3 s 0 8984 800 9104 4 chanx_left_in[11]
port 15 nsew
rlabel metal3 s 0 9392 800 9512 4 chanx_left_in[12]
port 16 nsew
rlabel metal3 s 0 9936 800 10056 4 chanx_left_in[13]
port 17 nsew
rlabel metal3 s 0 10344 800 10464 4 chanx_left_in[14]
port 18 nsew
rlabel metal3 s 0 10752 800 10872 4 chanx_left_in[15]
port 19 nsew
rlabel metal3 s 0 11296 800 11416 4 chanx_left_in[16]
port 20 nsew
rlabel metal3 s 0 11704 800 11824 4 chanx_left_in[17]
port 21 nsew
rlabel metal3 s 0 12248 800 12368 4 chanx_left_in[18]
port 22 nsew
rlabel metal3 s 0 12656 800 12776 4 chanx_left_in[19]
port 23 nsew
rlabel metal3 s 0 4224 800 4344 4 chanx_left_in[1]
port 24 nsew
rlabel metal3 s 0 4768 800 4888 4 chanx_left_in[2]
port 25 nsew
rlabel metal3 s 0 5176 800 5296 4 chanx_left_in[3]
port 26 nsew
rlabel metal3 s 0 5720 800 5840 4 chanx_left_in[4]
port 27 nsew
rlabel metal3 s 0 6128 800 6248 4 chanx_left_in[5]
port 28 nsew
rlabel metal3 s 0 6672 800 6792 4 chanx_left_in[6]
port 29 nsew
rlabel metal3 s 0 7080 800 7200 4 chanx_left_in[7]
port 30 nsew
rlabel metal3 s 0 7488 800 7608 4 chanx_left_in[8]
port 31 nsew
rlabel metal3 s 0 8032 800 8152 4 chanx_left_in[9]
port 32 nsew
rlabel metal3 s 0 13200 800 13320 4 chanx_left_out[0]
port 33 nsew
rlabel metal3 s 0 17824 800 17944 4 chanx_left_out[10]
port 34 nsew
rlabel metal3 s 0 18232 800 18352 4 chanx_left_out[11]
port 35 nsew
rlabel metal3 s 0 18776 800 18896 4 chanx_left_out[12]
port 36 nsew
rlabel metal3 s 0 19184 800 19304 4 chanx_left_out[13]
port 37 nsew
rlabel metal3 s 0 19728 800 19848 4 chanx_left_out[14]
port 38 nsew
rlabel metal3 s 0 20136 800 20256 4 chanx_left_out[15]
port 39 nsew
rlabel metal3 s 0 20544 800 20664 4 chanx_left_out[16]
port 40 nsew
rlabel metal3 s 0 21088 800 21208 4 chanx_left_out[17]
port 41 nsew
rlabel metal3 s 0 21496 800 21616 4 chanx_left_out[18]
port 42 nsew
rlabel metal3 s 0 22040 800 22160 4 chanx_left_out[19]
port 43 nsew
rlabel metal3 s 0 13608 800 13728 4 chanx_left_out[1]
port 44 nsew
rlabel metal3 s 0 14016 800 14136 4 chanx_left_out[2]
port 45 nsew
rlabel metal3 s 0 14560 800 14680 4 chanx_left_out[3]
port 46 nsew
rlabel metal3 s 0 14968 800 15088 4 chanx_left_out[4]
port 47 nsew
rlabel metal3 s 0 15512 800 15632 4 chanx_left_out[5]
port 48 nsew
rlabel metal3 s 0 15920 800 16040 4 chanx_left_out[6]
port 49 nsew
rlabel metal3 s 0 16464 800 16584 4 chanx_left_out[7]
port 50 nsew
rlabel metal3 s 0 16872 800 16992 4 chanx_left_out[8]
port 51 nsew
rlabel metal3 s 0 17280 800 17400 4 chanx_left_out[9]
port 52 nsew
rlabel metal3 s 22000 3816 22800 3936 4 chanx_right_in[0]
port 53 nsew
rlabel metal3 s 22000 8440 22800 8560 4 chanx_right_in[10]
port 54 nsew
rlabel metal3 s 22000 8984 22800 9104 4 chanx_right_in[11]
port 55 nsew
rlabel metal3 s 22000 9392 22800 9512 4 chanx_right_in[12]
port 56 nsew
rlabel metal3 s 22000 9936 22800 10056 4 chanx_right_in[13]
port 57 nsew
rlabel metal3 s 22000 10344 22800 10464 4 chanx_right_in[14]
port 58 nsew
rlabel metal3 s 22000 10752 22800 10872 4 chanx_right_in[15]
port 59 nsew
rlabel metal3 s 22000 11296 22800 11416 4 chanx_right_in[16]
port 60 nsew
rlabel metal3 s 22000 11704 22800 11824 4 chanx_right_in[17]
port 61 nsew
rlabel metal3 s 22000 12248 22800 12368 4 chanx_right_in[18]
port 62 nsew
rlabel metal3 s 22000 12656 22800 12776 4 chanx_right_in[19]
port 63 nsew
rlabel metal3 s 22000 4224 22800 4344 4 chanx_right_in[1]
port 64 nsew
rlabel metal3 s 22000 4768 22800 4888 4 chanx_right_in[2]
port 65 nsew
rlabel metal3 s 22000 5176 22800 5296 4 chanx_right_in[3]
port 66 nsew
rlabel metal3 s 22000 5720 22800 5840 4 chanx_right_in[4]
port 67 nsew
rlabel metal3 s 22000 6128 22800 6248 4 chanx_right_in[5]
port 68 nsew
rlabel metal3 s 22000 6672 22800 6792 4 chanx_right_in[6]
port 69 nsew
rlabel metal3 s 22000 7080 22800 7200 4 chanx_right_in[7]
port 70 nsew
rlabel metal3 s 22000 7488 22800 7608 4 chanx_right_in[8]
port 71 nsew
rlabel metal3 s 22000 8032 22800 8152 4 chanx_right_in[9]
port 72 nsew
rlabel metal3 s 22000 13200 22800 13320 4 chanx_right_out[0]
port 73 nsew
rlabel metal3 s 22000 17824 22800 17944 4 chanx_right_out[10]
port 74 nsew
rlabel metal3 s 22000 18232 22800 18352 4 chanx_right_out[11]
port 75 nsew
rlabel metal3 s 22000 18776 22800 18896 4 chanx_right_out[12]
port 76 nsew
rlabel metal3 s 22000 19184 22800 19304 4 chanx_right_out[13]
port 77 nsew
rlabel metal3 s 22000 19728 22800 19848 4 chanx_right_out[14]
port 78 nsew
rlabel metal3 s 22000 20136 22800 20256 4 chanx_right_out[15]
port 79 nsew
rlabel metal3 s 22000 20544 22800 20664 4 chanx_right_out[16]
port 80 nsew
rlabel metal3 s 22000 21088 22800 21208 4 chanx_right_out[17]
port 81 nsew
rlabel metal3 s 22000 21496 22800 21616 4 chanx_right_out[18]
port 82 nsew
rlabel metal3 s 22000 22040 22800 22160 4 chanx_right_out[19]
port 83 nsew
rlabel metal3 s 22000 13608 22800 13728 4 chanx_right_out[1]
port 84 nsew
rlabel metal3 s 22000 14016 22800 14136 4 chanx_right_out[2]
port 85 nsew
rlabel metal3 s 22000 14560 22800 14680 4 chanx_right_out[3]
port 86 nsew
rlabel metal3 s 22000 14968 22800 15088 4 chanx_right_out[4]
port 87 nsew
rlabel metal3 s 22000 15512 22800 15632 4 chanx_right_out[5]
port 88 nsew
rlabel metal3 s 22000 15920 22800 16040 4 chanx_right_out[6]
port 89 nsew
rlabel metal3 s 22000 16464 22800 16584 4 chanx_right_out[7]
port 90 nsew
rlabel metal3 s 22000 16872 22800 16992 4 chanx_right_out[8]
port 91 nsew
rlabel metal3 s 22000 17280 22800 17400 4 chanx_right_out[9]
port 92 nsew
rlabel metal2 s 3698 0 3754 800 4 chany_bottom_in[0]
port 93 nsew
rlabel metal2 s 8206 0 8262 800 4 chany_bottom_in[10]
port 94 nsew
rlabel metal2 s 8666 0 8722 800 4 chany_bottom_in[11]
port 95 nsew
rlabel metal2 s 9126 0 9182 800 4 chany_bottom_in[12]
port 96 nsew
rlabel metal2 s 9586 0 9642 800 4 chany_bottom_in[13]
port 97 nsew
rlabel metal2 s 9954 0 10010 800 4 chany_bottom_in[14]
port 98 nsew
rlabel metal2 s 10414 0 10470 800 4 chany_bottom_in[15]
port 99 nsew
rlabel metal2 s 10874 0 10930 800 4 chany_bottom_in[16]
port 100 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_in[17]
port 101 nsew
rlabel metal2 s 11794 0 11850 800 4 chany_bottom_in[18]
port 102 nsew
rlabel metal2 s 12254 0 12310 800 4 chany_bottom_in[19]
port 103 nsew
rlabel metal2 s 4158 0 4214 800 4 chany_bottom_in[1]
port 104 nsew
rlabel metal2 s 4618 0 4674 800 4 chany_bottom_in[2]
port 105 nsew
rlabel metal2 s 5078 0 5134 800 4 chany_bottom_in[3]
port 106 nsew
rlabel metal2 s 5538 0 5594 800 4 chany_bottom_in[4]
port 107 nsew
rlabel metal2 s 5998 0 6054 800 4 chany_bottom_in[5]
port 108 nsew
rlabel metal2 s 6458 0 6514 800 4 chany_bottom_in[6]
port 109 nsew
rlabel metal2 s 6826 0 6882 800 4 chany_bottom_in[7]
port 110 nsew
rlabel metal2 s 7286 0 7342 800 4 chany_bottom_in[8]
port 111 nsew
rlabel metal2 s 7746 0 7802 800 4 chany_bottom_in[9]
port 112 nsew
rlabel metal2 s 12714 0 12770 800 4 chany_bottom_out[0]
port 113 nsew
rlabel metal2 s 17130 0 17186 800 4 chany_bottom_out[10]
port 114 nsew
rlabel metal2 s 17590 0 17646 800 4 chany_bottom_out[11]
port 115 nsew
rlabel metal2 s 18050 0 18106 800 4 chany_bottom_out[12]
port 116 nsew
rlabel metal2 s 18510 0 18566 800 4 chany_bottom_out[13]
port 117 nsew
rlabel metal2 s 18970 0 19026 800 4 chany_bottom_out[14]
port 118 nsew
rlabel metal2 s 19430 0 19486 800 4 chany_bottom_out[15]
port 119 nsew
rlabel metal2 s 19798 0 19854 800 4 chany_bottom_out[16]
port 120 nsew
rlabel metal2 s 20258 0 20314 800 4 chany_bottom_out[17]
port 121 nsew
rlabel metal2 s 20718 0 20774 800 4 chany_bottom_out[18]
port 122 nsew
rlabel metal2 s 21178 0 21234 800 4 chany_bottom_out[19]
port 123 nsew
rlabel metal2 s 13174 0 13230 800 4 chany_bottom_out[1]
port 124 nsew
rlabel metal2 s 13542 0 13598 800 4 chany_bottom_out[2]
port 125 nsew
rlabel metal2 s 14002 0 14058 800 4 chany_bottom_out[3]
port 126 nsew
rlabel metal2 s 14462 0 14518 800 4 chany_bottom_out[4]
port 127 nsew
rlabel metal2 s 14922 0 14978 800 4 chany_bottom_out[5]
port 128 nsew
rlabel metal2 s 15382 0 15438 800 4 chany_bottom_out[6]
port 129 nsew
rlabel metal2 s 15842 0 15898 800 4 chany_bottom_out[7]
port 130 nsew
rlabel metal2 s 16302 0 16358 800 4 chany_bottom_out[8]
port 131 nsew
rlabel metal2 s 16670 0 16726 800 4 chany_bottom_out[9]
port 132 nsew
rlabel metal3 s 0 144 800 264 4 left_bottom_grid_pin_34_
port 133 nsew
rlabel metal3 s 0 552 800 672 4 left_bottom_grid_pin_35_
port 134 nsew
rlabel metal3 s 0 960 800 1080 4 left_bottom_grid_pin_36_
port 135 nsew
rlabel metal3 s 0 1504 800 1624 4 left_bottom_grid_pin_37_
port 136 nsew
rlabel metal3 s 0 1912 800 2032 4 left_bottom_grid_pin_38_
port 137 nsew
rlabel metal3 s 0 2456 800 2576 4 left_bottom_grid_pin_39_
port 138 nsew
rlabel metal3 s 0 2864 800 2984 4 left_bottom_grid_pin_40_
port 139 nsew
rlabel metal3 s 0 3408 800 3528 4 left_bottom_grid_pin_41_
port 140 nsew
rlabel metal3 s 0 22448 800 22568 4 left_top_grid_pin_1_
port 141 nsew
rlabel metal2 s 22558 0 22614 800 4 prog_clk_0_S_in
port 142 nsew
rlabel metal3 s 22000 144 22800 264 4 right_bottom_grid_pin_34_
port 143 nsew
rlabel metal3 s 22000 552 22800 672 4 right_bottom_grid_pin_35_
port 144 nsew
rlabel metal3 s 22000 960 22800 1080 4 right_bottom_grid_pin_36_
port 145 nsew
rlabel metal3 s 22000 1504 22800 1624 4 right_bottom_grid_pin_37_
port 146 nsew
rlabel metal3 s 22000 1912 22800 2032 4 right_bottom_grid_pin_38_
port 147 nsew
rlabel metal3 s 22000 2456 22800 2576 4 right_bottom_grid_pin_39_
port 148 nsew
rlabel metal3 s 22000 2864 22800 2984 4 right_bottom_grid_pin_40_
port 149 nsew
rlabel metal3 s 22000 3408 22800 3528 4 right_bottom_grid_pin_41_
port 150 nsew
rlabel metal3 s 22000 22448 22800 22568 4 right_top_grid_pin_1_
port 151 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 152 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 153 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_1__2_/results/magic/sb_1__2_.gds
string GDS_END 1165972
string GDS_START 81916
<< end >>
